//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(G2106), .B1(G567), .B2(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G113), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(G2105), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n467), .A2(new_n469), .B1(G101), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n468), .A2(G137), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(KEYINPUT3), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(new_n466), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(KEYINPUT68), .ZN(new_n479));
  OAI211_X1 g054(.A(KEYINPUT69), .B(G2104), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n472), .A2(new_n475), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n471), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n475), .A2(new_n481), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n486), .A2(new_n480), .A3(new_n469), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G2105), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n486), .A2(new_n490), .A3(new_n480), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n491), .A2(new_n494), .A3(G136), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G162));
  NAND4_X1  g071(.A1(new_n475), .A2(G126), .A3(new_n480), .A4(new_n481), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n468), .A2(new_n463), .A3(G138), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n500), .A2(new_n501), .B1(G102), .B2(new_n470), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n490), .A2(KEYINPUT67), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  AND4_X1   g080(.A1(KEYINPUT4), .A2(new_n503), .A3(new_n505), .A4(G138), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n475), .A2(new_n506), .A3(new_n480), .A4(new_n481), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n499), .A2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n511), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(G651), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT73), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  NAND3_X1  g102(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G51), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI221_X1 g105(.A(new_n528), .B1(new_n514), .B2(new_n529), .C1(new_n530), .C2(new_n512), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n512), .A2(new_n533), .B1(new_n514), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT74), .Z(new_n536));
  AOI22_X1  g111(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT75), .B(G43), .Z(new_n543));
  OAI22_X1  g118(.A1(new_n512), .A2(new_n542), .B1(new_n514), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n538), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AND2_X1   g128(.A1(new_n510), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(new_n512), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G91), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n556), .B(new_n558), .C1(new_n538), .C2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G168), .ZN(G286));
  INV_X1    g136(.A(G166), .ZN(G303));
  INV_X1    g137(.A(G87), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n512), .A2(KEYINPUT76), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n512), .B2(new_n563), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G49), .B2(new_n554), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT77), .Z(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G288));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n512), .A2(new_n570), .B1(new_n514), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n538), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT78), .Z(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  INV_X1    g152(.A(G85), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n512), .A2(new_n578), .B1(new_n514), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT80), .Z(new_n581));
  NAND2_X1  g156(.A1(G72), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G60), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n518), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n538), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(new_n585), .B2(new_n584), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n518), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n538), .B1(new_n592), .B2(KEYINPUT83), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(KEYINPUT83), .B2(new_n592), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n595), .B1(new_n514), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(new_n514), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n511), .A2(new_n510), .A3(G92), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(KEYINPUT10), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n589), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n589), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(KEYINPUT84), .B1(new_n607), .B2(new_n547), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT84), .B2(new_n614), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT85), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n463), .A2(new_n470), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2100), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n491), .A2(G135), .ZN(new_n623));
  OAI221_X1 g198(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n624));
  INV_X1    g199(.A(G123), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n623), .B(new_n624), .C1(new_n487), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT14), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n635), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(G401));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT86), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n444), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(KEYINPUT17), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n647), .A3(new_n649), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT87), .Z(new_n657));
  INV_X1    g232(.A(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n649), .B1(new_n658), .B2(new_n648), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n648), .B2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT20), .Z(new_n674));
  AOI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT89), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n576), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT91), .Z(new_n686));
  XOR2_X1   g261(.A(KEYINPUT32), .B(G1981), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G22), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G166), .B2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(KEYINPUT92), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n692), .B2(KEYINPUT92), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n688), .A2(KEYINPUT34), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT34), .B1(new_n688), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n491), .A2(G131), .ZN(new_n704));
  OAI221_X1 g279(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n705));
  INV_X1    g280(.A(G119), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n704), .B(new_n705), .C1(new_n487), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G25), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n694), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G290), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n694), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT90), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n702), .A2(new_n703), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT36), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n702), .A2(new_n720), .A3(new_n703), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n694), .A2(G20), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT23), .Z(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G299), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1956), .ZN(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n728), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n726), .B1(new_n733), .B2(KEYINPUT94), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(KEYINPUT94), .B2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n626), .A2(new_n728), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n694), .A2(G5), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G171), .B2(new_n694), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1961), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n743), .A2(new_n744), .B1(G105), .B2(new_n470), .ZN(new_n745));
  INV_X1    g320(.A(G129), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n487), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G141), .B2(new_n491), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n728), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n728), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n737), .B(new_n740), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n694), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n752), .B(new_n757), .C1(new_n750), .C2(new_n751), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n728), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n491), .A2(G140), .ZN(new_n761));
  OAI221_X1 g336(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n762));
  INV_X1    g337(.A(G128), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n761), .B(new_n762), .C1(new_n487), .C2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(new_n728), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n728), .B1(new_n768), .B2(G28), .ZN(new_n770));
  AND2_X1   g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NOR2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n694), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n694), .B2(G19), .ZN(new_n775));
  INV_X1    g350(.A(G1341), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n776), .B2(new_n775), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n694), .A2(G21), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G168), .B2(new_n694), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1966), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n728), .B1(KEYINPUT24), .B2(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(KEYINPUT24), .B2(G34), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n483), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n778), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n728), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n728), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(new_n443), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n728), .A2(G33), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n468), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n491), .B2(G139), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n791), .B1(new_n796), .B2(new_n728), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(new_n442), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n787), .A2(new_n790), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n758), .A2(new_n767), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n735), .A2(KEYINPUT95), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n731), .A2(new_n727), .A3(new_n732), .ZN(new_n802));
  AND4_X1   g377(.A1(new_n736), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n722), .A2(new_n803), .ZN(G311));
  AND3_X1   g379(.A1(new_n722), .A2(KEYINPUT96), .A3(new_n803), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT96), .B1(new_n722), .B2(new_n803), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(G150));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G67), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n518), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n538), .B1(new_n810), .B2(KEYINPUT97), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT97), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n554), .A2(G55), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n557), .A2(G93), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT99), .B(G860), .Z(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n547), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n604), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT98), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n823), .B2(new_n824), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n764), .B(G164), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n748), .ZN(new_n830));
  INV_X1    g405(.A(new_n796), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n707), .B(KEYINPUT101), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(new_n620), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n620), .ZN(new_n837));
  OAI221_X1 g412(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n838));
  INV_X1    g413(.A(G130), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n487), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G142), .B2(new_n491), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OR3_X1    g417(.A1(new_n836), .A2(new_n837), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n836), .B2(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT103), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n832), .A2(new_n843), .A3(new_n844), .A4(new_n833), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT102), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n626), .B(G160), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(G162), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT104), .B(G37), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n854), .B1(new_n845), .B2(new_n834), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n849), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n855), .A2(new_n859), .A3(KEYINPUT40), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT40), .B1(new_n855), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(G395));
  XNOR2_X1  g437(.A(new_n576), .B(new_n696), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n713), .B(G166), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n604), .B(G299), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n755), .B(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n613), .B(new_n820), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n875), .B2(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n867), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n867), .ZN(new_n882));
  OAI21_X1  g457(.A(G868), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n815), .A2(new_n607), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(G295));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(G331));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  XNOR2_X1  g462(.A(G301), .B(G286), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n820), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n889), .A2(new_n872), .ZN(new_n890));
  INV_X1    g465(.A(new_n873), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n871), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(KEYINPUT108), .A3(new_n820), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n889), .B2(KEYINPUT108), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n865), .B(new_n890), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n856), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n870), .A2(new_n873), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(new_n889), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g475(.A1(new_n898), .A2(new_n899), .B1(new_n868), .B2(new_n894), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n865), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT110), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  INV_X1    g479(.A(new_n865), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT110), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n906), .A2(new_n907), .A3(new_n856), .A4(new_n895), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n887), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n905), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n911), .A2(new_n912), .A3(new_n895), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n906), .A2(new_n887), .A3(new_n856), .A4(new_n895), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n913), .B2(new_n887), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(G397));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n499), .B2(new_n508), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n471), .A2(G40), .A3(new_n482), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n924), .A2(KEYINPUT111), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT111), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n713), .A2(new_n681), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT112), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n713), .A2(new_n681), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n748), .B(G1996), .ZN(new_n934));
  INV_X1    g509(.A(G2067), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n764), .B(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n707), .B(new_n709), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n929), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT45), .B(new_n921), .C1(new_n499), .C2(new_n508), .ZN(new_n941));
  INV_X1    g516(.A(new_n925), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n924), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n922), .A2(KEYINPUT113), .A3(new_n923), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT53), .B1(new_n947), .B2(new_n443), .ZN(new_n948));
  NOR2_X1   g523(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(new_n499), .B2(new_n508), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n925), .B1(new_n950), .B2(KEYINPUT114), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n497), .A2(new_n498), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G2105), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n502), .A2(new_n507), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n949), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1961), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n941), .A2(new_n942), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n924), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(G171), .B1(new_n948), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n522), .A2(new_n523), .A3(G8), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n955), .B2(new_n921), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n942), .A2(new_n950), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n971), .A2(new_n972), .A3(G2090), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n922), .A2(KEYINPUT113), .A3(new_n923), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT113), .B1(new_n922), .B2(new_n923), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n962), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n976), .B2(new_n691), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT115), .B(G8), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n969), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n945), .A2(new_n946), .ZN(new_n980));
  AOI21_X1  g555(.A(G1971), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n959), .A2(G2090), .ZN(new_n982));
  OAI211_X1 g557(.A(G8), .B(new_n968), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n922), .A2(new_n925), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n696), .A2(G1976), .ZN(new_n986));
  INV_X1    g561(.A(new_n978), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT52), .ZN(new_n989));
  INV_X1    g564(.A(G1976), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n986), .A3(new_n991), .A4(new_n987), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n575), .A2(G1981), .ZN(new_n993));
  OR3_X1    g568(.A1(new_n572), .A2(new_n574), .A3(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n985), .A2(new_n997), .A3(new_n987), .A4(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n989), .A2(new_n992), .A3(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n979), .A2(new_n983), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1966), .ZN(new_n1002));
  INV_X1    g577(.A(new_n924), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n943), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n951), .A2(new_n957), .A3(new_n785), .A4(new_n958), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G168), .A2(new_n978), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT118), .Z(new_n1009));
  AOI21_X1  g584(.A(new_n978), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1010), .A2(KEYINPUT120), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1007), .A2(KEYINPUT51), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT120), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1007), .B(KEYINPUT119), .Z(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1006), .B2(G8), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1011), .A2(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n965), .B(new_n1001), .C1(new_n1018), .C2(KEYINPUT62), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(KEYINPUT62), .B2(new_n1018), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1000), .B(KEYINPUT116), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1010), .A2(G168), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n981), .B2(new_n982), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n969), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n983), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(new_n1001), .B2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n999), .A2(new_n990), .A3(new_n696), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n978), .B(new_n984), .C1(new_n1030), .C2(new_n994), .ZN(new_n1031));
  INV_X1    g606(.A(new_n983), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT56), .B(G2072), .Z(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n980), .A2(new_n962), .A3(new_n1036), .ZN(new_n1037));
  XOR2_X1   g612(.A(G299), .B(KEYINPUT57), .Z(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT117), .B(G1956), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n971), .B2(new_n972), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1348), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n959), .A2(new_n1043), .B1(new_n935), .B2(new_n984), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(new_n755), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n976), .B2(new_n1035), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1038), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1042), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n755), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(new_n1050), .A3(new_n604), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(new_n962), .C1(new_n974), .C2(new_n975), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT58), .B(G1341), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n985), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n547), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1053), .B1(KEYINPUT59), .B2(new_n1058), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1058), .A2(KEYINPUT59), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1052), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1048), .A2(KEYINPUT61), .A3(new_n1041), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT61), .B1(new_n1048), .B2(new_n1041), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1049), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n1066));
  OR2_X1    g641(.A1(KEYINPUT122), .A2(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(KEYINPUT122), .A2(G2078), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n924), .A2(new_n942), .A3(new_n941), .A4(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n443), .B(new_n962), .C1(new_n974), .C2(new_n975), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1066), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n959), .B2(new_n960), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n959), .A2(new_n1073), .A3(new_n960), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n948), .A2(new_n964), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(G301), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1001), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1072), .B(G301), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n965), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT123), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1085), .B(KEYINPUT54), .C1(new_n1082), .C2(new_n965), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1081), .B(new_n1018), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1065), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n965), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT123), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1091), .A2(KEYINPUT124), .A3(new_n1018), .A4(new_n1081), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1034), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1020), .B1(new_n1093), .B2(KEYINPUT125), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1095), .B(new_n1034), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n940), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n707), .A2(new_n710), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n937), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n765), .A2(new_n935), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n928), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT48), .B1(new_n931), .B2(new_n929), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n939), .B2(new_n929), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n931), .A2(KEYINPUT48), .A3(new_n929), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n928), .B1(new_n936), .B2(new_n748), .ZN(new_n1106));
  XOR2_X1   g681(.A(new_n1106), .B(KEYINPUT126), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n929), .A2(new_n1054), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT46), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT47), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1105), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1111), .B2(new_n1110), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1097), .A2(new_n1113), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g689(.A1(new_n664), .A2(G319), .A3(new_n644), .ZN(new_n1116));
  XOR2_X1   g690(.A(new_n1116), .B(KEYINPUT127), .Z(new_n1117));
  NOR2_X1   g691(.A1(new_n1117), .A2(G229), .ZN(new_n1118));
  AOI21_X1  g692(.A(new_n853), .B1(new_n847), .B2(new_n849), .ZN(new_n1119));
  INV_X1    g693(.A(new_n859), .ZN(new_n1120));
  OAI211_X1 g694(.A(new_n917), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G225));
  INV_X1    g695(.A(G225), .ZN(G308));
endmodule


