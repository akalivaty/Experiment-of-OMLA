//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(new_n195), .A3(new_n199), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n204), .A2(new_n205), .B1(G104), .B2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(G104), .A3(new_n206), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT80), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(G104), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(new_n203), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n210), .A4(new_n208), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(G101), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G101), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n219), .A3(new_n210), .A4(new_n208), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT64), .A3(G143), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(G146), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n223), .A2(G143), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n229), .A2(new_n232), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n212), .A2(new_n236), .A3(G101), .A4(new_n217), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n222), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n213), .A2(new_n210), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n223), .A2(G143), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n242), .B(KEYINPUT1), .C1(new_n226), .C2(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n229), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n226), .A2(G146), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n248), .A3(new_n249), .A4(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n241), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n250), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT1), .B1(new_n226), .B2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(G128), .A3(new_n245), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n254), .B1(new_n257), .B2(new_n229), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n220), .A2(KEYINPUT10), .A3(new_n240), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT81), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n249), .B1(G143), .B2(new_n223), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n250), .B1(new_n264), .B2(new_n234), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n220), .A3(new_n240), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT10), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND4_X1   g082(.A1(new_n202), .A2(new_n238), .A3(new_n261), .A4(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n253), .A2(new_n260), .B1(new_n267), .B2(new_n266), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n202), .B1(new_n270), .B2(new_n238), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n190), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n238), .A2(new_n261), .A3(new_n202), .A4(new_n268), .ZN(new_n273));
  INV_X1    g087(.A(new_n190), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n220), .A2(new_n240), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n250), .A3(new_n247), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n266), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n277), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n201), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n202), .B1(new_n276), .B2(new_n266), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(KEYINPUT12), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT82), .B1(new_n279), .B2(KEYINPUT12), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n273), .B(new_n274), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G469), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n272), .B2(new_n282), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT83), .A3(new_n284), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n201), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT12), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n278), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n274), .B1(new_n296), .B2(new_n273), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n269), .A2(new_n271), .A3(new_n190), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n285), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n288), .A2(new_n290), .B1(G469), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n301), .B(KEYINPUT84), .Z(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n229), .A2(new_n232), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n234), .A2(new_n230), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G125), .ZN(new_n307));
  INV_X1    g121(.A(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n258), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G224), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G953), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT66), .B1(new_n314), .B2(G119), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G113), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G113), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT67), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n317), .B2(G116), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n314), .A2(KEYINPUT67), .A3(G119), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n319), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT68), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n326), .A2(new_n327), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n324), .A4(new_n319), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n324), .B1(new_n330), .B2(new_n319), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n222), .A3(new_n237), .ZN(new_n337));
  INV_X1    g151(.A(new_n275), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(KEYINPUT5), .A3(new_n319), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n314), .A2(G119), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n320), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT86), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT85), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n344), .A4(new_n348), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n345), .B2(new_n349), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n313), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G210), .B1(G237), .B2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n348), .B(KEYINPUT8), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n333), .A2(new_n338), .A3(new_n343), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n338), .B1(new_n333), .B2(new_n343), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT87), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT87), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n361), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n312), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT7), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n310), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT7), .A4(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n237), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n334), .B1(new_n329), .B2(new_n332), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n357), .B1(new_n371), .B2(new_n222), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n368), .B1(new_n372), .B2(new_n348), .ZN(new_n373));
  AOI21_X1  g187(.A(G902), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n354), .A2(new_n355), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n355), .B1(new_n354), .B2(new_n374), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n303), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  OAI21_X1  g192(.A(G221), .B1(new_n378), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n300), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n192), .A2(G137), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n194), .A2(G134), .ZN(new_n384));
  OAI21_X1  g198(.A(G131), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n200), .A2(new_n385), .ZN(new_n386));
  OAI22_X1  g200(.A1(new_n202), .A2(new_n306), .B1(new_n258), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n336), .ZN(new_n388));
  INV_X1    g202(.A(new_n386), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n263), .B1(new_n262), .B2(new_n242), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n243), .B1(new_n233), .B2(new_n225), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n390), .A2(new_n256), .B1(new_n391), .B2(new_n224), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n389), .B1(new_n392), .B2(new_n254), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n235), .A2(new_n201), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n370), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n382), .B1(new_n388), .B2(new_n395), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n395), .A2(new_n382), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT72), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n387), .A2(new_n336), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n393), .A2(new_n394), .B1(new_n333), .B2(new_n335), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n404));
  NOR2_X1   g218(.A1(G237), .A2(G953), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G210), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n404), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT26), .B(G101), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n403), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n285), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT73), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(new_n285), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n396), .A2(new_n397), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n409), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n370), .B1(new_n387), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n235), .B2(new_n201), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n421), .A2(new_n393), .A3(KEYINPUT69), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT69), .B1(new_n421), .B2(new_n393), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT70), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n420), .B(new_n426), .C1(new_n423), .C2(new_n422), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n399), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n418), .B1(new_n428), .B2(new_n409), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n414), .B(new_n416), .C1(KEYINPUT29), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G472), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n399), .A2(new_n409), .ZN(new_n432));
  INV_X1    g246(.A(new_n427), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n394), .A2(KEYINPUT30), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n258), .A2(new_n386), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n421), .A2(new_n393), .A3(KEYINPUT69), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n426), .B1(new_n439), .B2(new_n420), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT31), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n409), .B1(new_n396), .B2(new_n397), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n425), .A2(new_n427), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT31), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n432), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(G472), .A2(G902), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n447), .A2(KEYINPUT32), .A3(new_n448), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n431), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G217), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(G234), .B2(new_n285), .ZN(new_n455));
  INV_X1    g269(.A(G140), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n308), .A2(G140), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT16), .ZN(new_n459));
  OR3_X1    g273(.A1(new_n308), .A2(KEYINPUT16), .A3(G140), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n223), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n458), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n223), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT23), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n317), .B2(G128), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n317), .A2(G128), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n263), .A2(KEYINPUT23), .A3(G119), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G110), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT74), .B1(new_n263), .B2(G119), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT74), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n317), .A3(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n263), .A2(G119), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT24), .B(G110), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n472), .A2(new_n479), .A3(KEYINPUT76), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT76), .B1(new_n472), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n465), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n477), .A2(KEYINPUT75), .A3(new_n478), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT75), .B1(new_n477), .B2(new_n478), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n470), .A2(new_n471), .ZN(new_n486));
  AOI21_X1  g300(.A(G146), .B1(new_n459), .B2(new_n460), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n462), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT22), .B(G137), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n482), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n482), .B2(new_n488), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT25), .B1(new_n494), .B2(new_n285), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n482), .A2(new_n488), .ZN(new_n496));
  INV_X1    g310(.A(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n488), .A3(new_n491), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n498), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n455), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n494), .B(KEYINPUT77), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n455), .A2(G902), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT78), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n502), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n188), .A3(G214), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n226), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n405), .B2(G214), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n226), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n405), .A2(G143), .A3(G214), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n199), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n462), .A2(new_n487), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n513), .A2(KEYINPUT91), .A3(new_n514), .A4(new_n517), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n513), .A2(new_n514), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n463), .A2(KEYINPUT88), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n463), .A2(KEYINPUT88), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(G146), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n464), .A2(new_n223), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n515), .B(new_n516), .C1(new_n530), .C2(new_n199), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT18), .B(G131), .C1(new_n511), .C2(new_n512), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G113), .B(G122), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT90), .B(G104), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n534), .B(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n524), .A2(new_n533), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n524), .B2(new_n533), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n285), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(KEYINPUT92), .B(new_n285), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(G475), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n525), .A2(KEYINPUT19), .A3(new_n526), .ZN(new_n544));
  OR3_X1    g358(.A1(new_n463), .A2(KEYINPUT89), .A3(KEYINPUT19), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT89), .B1(new_n463), .B2(KEYINPUT19), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n544), .A2(new_n223), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n462), .B1(new_n513), .B2(new_n517), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n536), .B1(new_n549), .B2(new_n533), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n537), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G475), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n285), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT20), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n524), .A2(new_n533), .A3(new_n536), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n532), .A2(new_n531), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n528), .B2(new_n527), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n547), .B2(new_n548), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n555), .B1(new_n558), .B2(new_n536), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n552), .A4(new_n285), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n543), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n226), .A2(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n263), .A2(G143), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n192), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(G134), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n572), .A3(G134), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(new_n568), .A3(new_n572), .A4(G134), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n314), .A2(G122), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT93), .ZN(new_n577));
  INV_X1    g391(.A(G122), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G116), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n577), .A2(new_n206), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n206), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n574), .B(new_n575), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n577), .A2(KEYINPUT14), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n577), .A2(KEYINPUT14), .B1(G116), .B2(new_n578), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n206), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n577), .A2(new_n206), .A3(new_n579), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n570), .A3(new_n571), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n582), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n378), .A2(new_n454), .A3(G953), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n582), .B(new_n589), .C1(new_n585), .C2(new_n587), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n566), .B1(new_n593), .B2(new_n285), .ZN(new_n594));
  AOI211_X1 g408(.A(G902), .B(new_n565), .C1(new_n591), .C2(new_n592), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G234), .A2(G237), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(G952), .A3(new_n188), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT94), .Z(new_n600));
  AND3_X1   g414(.A1(new_n598), .A2(G902), .A3(G953), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT21), .B(G898), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n563), .A2(new_n597), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n381), .A2(new_n453), .A3(new_n508), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  INV_X1    g421(.A(new_n449), .ZN(new_n608));
  INV_X1    g422(.A(G472), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n447), .B2(new_n285), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n604), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n303), .B(new_n612), .C1(new_n375), .C2(new_n376), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n593), .A2(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n591), .A2(new_n615), .A3(new_n592), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(G478), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n564), .A2(new_n285), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n591), .B2(new_n592), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n564), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n563), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n288), .A2(new_n290), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n299), .A2(G469), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n380), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n611), .A2(new_n624), .A3(new_n627), .A4(new_n508), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  AND2_X1   g444(.A1(new_n543), .A2(new_n562), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n597), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n611), .A2(new_n633), .A3(new_n627), .A4(new_n508), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT95), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n496), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n505), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n502), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n455), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n498), .A2(new_n285), .A3(new_n499), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT25), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n643), .B1(new_n646), .B2(new_n500), .ZN(new_n647));
  INV_X1    g461(.A(new_n641), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT96), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n608), .A2(new_n610), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n381), .A2(new_n651), .A3(new_n605), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  AND3_X1   g468(.A1(new_n447), .A2(KEYINPUT32), .A3(new_n448), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT32), .B1(new_n447), .B2(new_n448), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n650), .B1(new_n657), .B2(new_n431), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n289), .A2(KEYINPUT83), .A3(new_n284), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT83), .B1(new_n289), .B2(new_n284), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n626), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n354), .A2(new_n374), .ZN(new_n662));
  INV_X1    g476(.A(new_n355), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n354), .A2(new_n374), .A3(new_n355), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n302), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n601), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n600), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n563), .A2(new_n596), .A3(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n379), .A2(new_n661), .A3(new_n666), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n658), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT97), .B(G128), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G30));
  INV_X1    g488(.A(new_n428), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n410), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n409), .A2(new_n388), .A3(new_n395), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n428), .B2(new_n409), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(KEYINPUT98), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n609), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n655), .A3(new_n656), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n375), .A2(new_n376), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n375), .B2(new_n376), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n596), .B1(new_n543), .B2(new_n562), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n647), .A2(new_n648), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n303), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n683), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n669), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n627), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  NOR3_X1   g512(.A1(new_n650), .A2(new_n623), .A3(new_n669), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n381), .A2(new_n453), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n381), .A2(new_n453), .A3(KEYINPUT99), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  NAND3_X1  g519(.A1(new_n238), .A2(new_n261), .A3(new_n268), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n201), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n273), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n273), .A2(new_n274), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n190), .A2(new_n708), .B1(new_n709), .B2(new_n296), .ZN(new_n710));
  OAI211_X1 g524(.A(KEYINPUT100), .B(G469), .C1(new_n710), .C2(G902), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n289), .B2(new_n284), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n625), .A2(new_n714), .A3(new_n379), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n453), .A2(new_n624), .A3(new_n715), .A4(new_n508), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n453), .A2(new_n508), .A3(new_n715), .A4(new_n633), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT101), .B(G116), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G18));
  INV_X1    g535(.A(new_n650), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n453), .A2(new_n605), .A3(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n666), .A2(new_n379), .A3(new_n625), .A4(new_n714), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n288), .A2(new_n290), .B1(new_n711), .B2(new_n713), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(KEYINPUT102), .A3(new_n379), .A4(new_n666), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n723), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n317), .ZN(G21));
  OAI211_X1 g544(.A(new_n689), .B(new_n303), .C1(new_n375), .C2(new_n376), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n604), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n447), .A2(new_n285), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n398), .A2(new_n403), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n442), .B(new_n446), .C1(new_n410), .C2(new_n734), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n733), .A2(G472), .B1(new_n448), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n715), .A2(new_n732), .A3(new_n508), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NAND2_X1  g552(.A1(new_n726), .A2(new_n728), .ZN(new_n739));
  INV_X1    g553(.A(new_n690), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n623), .A2(new_n669), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  AOI21_X1  g558(.A(new_n507), .B1(new_n657), .B2(new_n431), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n375), .A2(new_n376), .A3(new_n302), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n661), .A2(new_n746), .A3(new_n379), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n627), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n745), .A2(new_n741), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n452), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n447), .A2(KEYINPUT104), .A3(KEYINPUT32), .A4(new_n448), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n431), .A3(new_n451), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n623), .A2(new_n752), .A3(new_n669), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n508), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n749), .B1(new_n627), .B2(new_n746), .ZN(new_n760));
  AND4_X1   g574(.A1(new_n749), .A2(new_n661), .A3(new_n379), .A4(new_n746), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n762), .A3(KEYINPUT105), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n748), .A2(new_n750), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n757), .A2(new_n508), .A3(new_n758), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G131), .ZN(G33));
  NAND4_X1  g583(.A1(new_n745), .A2(new_n670), .A3(new_n748), .A4(new_n750), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n709), .A2(new_n707), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n296), .A2(new_n273), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT45), .B(new_n772), .C1(new_n773), .C2(new_n274), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n297), .B2(new_n298), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(G469), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT106), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n774), .A2(new_n776), .A3(KEYINPUT106), .A4(G469), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(G469), .A2(G902), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT107), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n625), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n781), .A2(new_n782), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n783), .B1(new_n779), .B2(new_n780), .ZN(new_n791));
  INV_X1    g605(.A(new_n625), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT107), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n787), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n379), .A3(new_n693), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n563), .B2(new_n621), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT43), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n608), .A2(new_n610), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n740), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT44), .A4(new_n740), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n746), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n795), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n194), .ZN(G39));
  XNOR2_X1  g620(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n794), .A2(new_n379), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n794), .B2(new_n379), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n741), .A2(new_n746), .A3(new_n507), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n453), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  XOR2_X1   g629(.A(new_n727), .B(KEYINPUT49), .Z(new_n816));
  INV_X1    g630(.A(new_n683), .ZN(new_n817));
  INV_X1    g631(.A(new_n688), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n507), .A2(new_n380), .A3(new_n302), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n631), .A3(new_n622), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT110), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  INV_X1    g638(.A(new_n669), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n690), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n731), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n627), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n683), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n702), .B2(new_n703), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n739), .A2(new_n742), .B1(new_n658), .B2(new_n671), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n824), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n833));
  INV_X1    g647(.A(new_n829), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n631), .A2(new_n621), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n649), .A3(new_n642), .A4(new_n825), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n657), .B2(new_n431), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT99), .B1(new_n837), .B2(new_n381), .ZN(new_n838));
  INV_X1    g652(.A(new_n703), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n743), .A2(new_n672), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n831), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n832), .B1(new_n844), .B2(new_n824), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n652), .A2(new_n737), .A3(new_n634), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n716), .A2(new_n719), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n729), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n606), .A2(new_n628), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n606), .A2(KEYINPUT111), .A3(new_n628), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n631), .A2(new_n596), .A3(new_n825), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT112), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n658), .A2(new_n627), .A3(new_n746), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n742), .A2(new_n748), .A3(new_n750), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n770), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n768), .A2(new_n848), .A3(new_n853), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT113), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n768), .A2(new_n848), .A3(new_n853), .A4(new_n858), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n845), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(KEYINPUT114), .A2(new_n704), .A3(new_n831), .A4(new_n834), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT114), .B1(new_n830), .B2(new_n831), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n824), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n843), .ZN(new_n870));
  AND4_X1   g684(.A1(KEYINPUT53), .A2(new_n869), .A3(new_n859), .A4(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n823), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n600), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n798), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n715), .A2(new_n746), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n508), .A3(new_n757), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n188), .A2(G952), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n508), .A2(new_n874), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n817), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n880), .B1(new_n882), .B2(new_n835), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n736), .A2(new_n508), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(new_n739), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n879), .B(new_n883), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n877), .A2(new_n740), .A3(new_n736), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n563), .A2(new_n622), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n882), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n882), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT50), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n303), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n688), .A2(new_n715), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n896), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n746), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n875), .A2(new_n884), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n727), .A2(new_n380), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n811), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n890), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n896), .A2(new_n903), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT115), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n808), .B2(new_n810), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n915), .A3(new_n908), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n912), .B1(new_n916), .B2(new_n907), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n911), .B1(new_n917), .B2(KEYINPUT51), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n869), .A2(new_n859), .A3(new_n870), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n865), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n861), .A2(new_n865), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n845), .A2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n920), .A2(new_n823), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n873), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n822), .B1(new_n924), .B2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n920), .A2(new_n922), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(G210), .A3(G902), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n352), .A2(new_n353), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT119), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n313), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n928), .B2(new_n929), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n188), .A2(G952), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(G51));
  XOR2_X1   g751(.A(new_n782), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n823), .B1(new_n920), .B2(new_n922), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n923), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n283), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n927), .A2(G902), .A3(new_n779), .A4(new_n780), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n927), .A2(G902), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n551), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n945), .B2(new_n551), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n927), .A2(G902), .A3(new_n559), .A4(new_n944), .ZN(new_n949));
  INV_X1    g763(.A(new_n936), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(G60));
  NAND2_X1  g766(.A1(new_n614), .A2(new_n616), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n919), .A2(new_n865), .B1(new_n845), .B2(new_n921), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n823), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n871), .B1(new_n865), .B2(new_n864), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n823), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n618), .B(KEYINPUT59), .Z(new_n958));
  AOI21_X1  g772(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n953), .A2(new_n958), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n923), .B2(new_n939), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n950), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n959), .A2(new_n962), .ZN(G63));
  XNOR2_X1  g777(.A(new_n503), .B(KEYINPUT122), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n454), .A2(new_n285), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n954), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n927), .A2(new_n640), .A3(new_n967), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n969), .A2(new_n970), .A3(new_n950), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT61), .A4(new_n950), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G66));
  AND2_X1   g789(.A1(new_n848), .A2(new_n853), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(G953), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT123), .ZN(new_n978));
  OAI21_X1  g792(.A(G953), .B1(new_n602), .B2(new_n311), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n931), .B1(G898), .B2(new_n188), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  NAND3_X1  g796(.A1(new_n697), .A2(new_n704), .A3(new_n831), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n697), .A2(new_n704), .A3(new_n831), .A4(KEYINPUT62), .ZN(new_n986));
  AOI22_X1  g800(.A1(new_n985), .A2(new_n986), .B1(new_n811), .B2(new_n813), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n906), .B1(new_n623), .B2(new_n632), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n745), .A2(new_n627), .A3(new_n988), .A4(new_n693), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n795), .B2(new_n804), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(KEYINPUT124), .B(new_n989), .C1(new_n795), .C2(new_n804), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT125), .B1(new_n987), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n188), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n387), .A2(new_n419), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n439), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n704), .A2(new_n831), .ZN(new_n1004));
  OR3_X1    g818(.A1(new_n805), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n805), .B2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n757), .A2(new_n508), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n795), .A2(new_n731), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n1009), .A2(new_n768), .A3(new_n770), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1007), .A2(new_n188), .A3(new_n814), .A4(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1002), .B1(G900), .B2(G953), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n997), .A2(new_n1002), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1013), .B(new_n1017), .ZN(G72));
  NOR2_X1   g832(.A1(new_n995), .A2(new_n996), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n976), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  AOI21_X1  g836(.A(new_n676), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1022), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n814), .A2(new_n768), .A3(new_n770), .A4(new_n1009), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1024), .B1(new_n1026), .B2(new_n976), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n675), .A2(new_n410), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n950), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n676), .A3(new_n1022), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n956), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n1023), .A2(new_n1030), .A3(new_n1032), .ZN(G57));
endmodule


