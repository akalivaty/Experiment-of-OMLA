//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n442, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1161,
    new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G108), .ZN(new_n442));
  INV_X1    g017(.A(new_n442), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n442), .A2(G57), .A3(G69), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT65), .Z(new_n453));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT66), .Z(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n462), .ZN(new_n468));
  OAI22_X1  g043(.A1(new_n464), .A2(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(new_n468), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  XOR2_X1   g050(.A(KEYINPUT3), .B(G2104), .Z(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND3_X1  g057(.A1(new_n467), .A2(G138), .A3(new_n462), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n467), .A2(KEYINPUT67), .A3(G138), .A4(new_n462), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n462), .A2(G102), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n476), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n488), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n483), .A2(new_n484), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n487), .A2(new_n492), .A3(new_n497), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n502), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n502), .A2(G543), .A3(new_n510), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n508), .A2(G62), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n511), .A2(G89), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n505), .B2(new_n507), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n522), .A2(new_n523), .A3(new_n527), .A4(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n524), .A2(new_n525), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(KEYINPUT73), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(G543), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n505), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(G64), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n542), .A2(new_n543), .A3(new_n534), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n536), .A2(G651), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n502), .A2(G52), .A3(G543), .A4(new_n510), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n502), .A2(G90), .A3(new_n508), .A4(new_n510), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n546), .B1(new_n545), .B2(new_n550), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n509), .ZN(new_n556));
  AOI22_X1  g131(.A1(G43), .A2(new_n521), .B1(new_n511), .B2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND3_X1  g140(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n511), .A2(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n514), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n509), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n566), .A2(new_n567), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G299));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND2_X1  g155(.A1(new_n521), .A2(G49), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n511), .A2(G87), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT76), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n583), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AND2_X1   g162(.A1(new_n508), .A2(G61), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(G651), .A2(new_n590), .B1(new_n521), .B2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n511), .A2(G86), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n511), .A2(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n514), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n526), .A2(G60), .ZN(new_n597));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n509), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n511), .A2(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n521), .A2(G54), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n508), .A2(G66), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n602), .B1(G868), .B2(new_n611), .ZN(G284));
  OAI21_X1  g187(.A(new_n602), .B1(G868), .B2(new_n611), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n578), .B(KEYINPUT78), .Z(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g198(.A(new_n463), .B(KEYINPUT66), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n467), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n474), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(G123), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT80), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT80), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G111), .C2(new_n462), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT82), .B(KEYINPUT14), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT81), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n653), .A2(KEYINPUT83), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n650), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(KEYINPUT83), .ZN(new_n656));
  NAND4_X1  g231(.A1(new_n654), .A2(G14), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT84), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n663), .B(KEYINPUT17), .Z(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n661), .A3(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n663), .A3(new_n659), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n676), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT85), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n681), .B1(new_n684), .B2(KEYINPUT20), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n680), .A3(new_n682), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n686), .C1(KEYINPUT20), .C2(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G32), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n474), .A2(G141), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n477), .A2(G129), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n624), .A2(G105), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT26), .Z(new_n700));
  NAND4_X1  g275(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n695), .B1(new_n702), .B2(new_n694), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT87), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT27), .B(G1996), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(G168), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G21), .ZN(new_n710));
  INV_X1    g285(.A(G1966), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n694), .A2(G26), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n474), .A2(G140), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n477), .A2(G128), .ZN(new_n715));
  OR2_X1    g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n694), .ZN(new_n720));
  MUX2_X1   g295(.A(new_n713), .B(new_n720), .S(KEYINPUT28), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G2067), .ZN(new_n722));
  AND4_X1   g297(.A1(new_n707), .A2(new_n708), .A3(new_n712), .A4(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(KEYINPUT24), .A2(G34), .ZN(new_n724));
  NAND2_X1  g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n694), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G160), .B2(new_n694), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n721), .A2(G2067), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n694), .A2(G33), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n474), .A2(G139), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT25), .Z(new_n734));
  AOI22_X1  g309(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n734), .C1(new_n462), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(G2072), .ZN(new_n739));
  INV_X1    g314(.A(new_n636), .ZN(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n740), .A2(G29), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G11), .ZN(new_n747));
  INV_X1    g322(.A(G2072), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n748), .C2(new_n737), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n559), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G19), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n739), .B(new_n749), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n723), .A2(new_n729), .A3(new_n730), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n694), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n694), .ZN(new_n756));
  MUX2_X1   g331(.A(new_n755), .B(new_n756), .S(KEYINPUT91), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT29), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2090), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n751), .A2(new_n752), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n710), .A2(new_n711), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT88), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n754), .A2(new_n759), .A3(new_n760), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G4), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n611), .B2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(G1348), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G5), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G171), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n764), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT92), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT23), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  INV_X1    g351(.A(G1956), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G27), .A2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2078), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n763), .A2(new_n768), .A3(new_n772), .A4(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n474), .A2(G131), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n477), .A2(G119), .ZN(new_n786));
  NOR2_X1   g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  MUX2_X1   g364(.A(G25), .B(new_n789), .S(G29), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT35), .B(G1991), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  NOR2_X1   g367(.A1(new_n600), .A2(new_n764), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n764), .B2(G24), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G22), .ZN(new_n797));
  OAI21_X1  g372(.A(KEYINPUT86), .B1(new_n797), .B2(G16), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n797), .A2(KEYINPUT86), .A3(G16), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(G166), .C2(new_n764), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n764), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(G288), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n764), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n801), .B1(new_n806), .B2(G1976), .ZN(new_n807));
  MUX2_X1   g382(.A(G6), .B(G305), .S(G16), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT32), .B(G1981), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n810), .C1(G1976), .C2(new_n806), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n796), .B1(new_n811), .B2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n794), .A2(new_n795), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n812), .B(new_n813), .C1(KEYINPUT34), .C2(new_n811), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n784), .B1(new_n815), .B2(new_n816), .ZN(G311));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n815), .ZN(new_n818));
  INV_X1    g393(.A(new_n784), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(G150));
  NAND2_X1  g395(.A1(new_n511), .A2(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n822), .B2(new_n514), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n526), .A2(G67), .ZN(new_n824));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n509), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT95), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n559), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n827), .A2(new_n558), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT38), .Z(new_n835));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n618), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  AOI21_X1  g413(.A(G860), .B1(new_n838), .B2(KEYINPUT94), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(KEYINPUT94), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(G145));
  XNOR2_X1  g417(.A(new_n495), .B(new_n718), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n702), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n474), .A2(KEYINPUT96), .A3(G142), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n477), .A2(G130), .ZN(new_n846));
  OR2_X1    g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  INV_X1    g424(.A(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n468), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n846), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n844), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n740), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n626), .B(KEYINPUT97), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n789), .B(KEYINPUT98), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n481), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n736), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g443(.A(G166), .B(new_n600), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(G305), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n803), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT42), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n611), .B1(new_n576), .B2(new_n577), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n578), .A2(new_n610), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n578), .B2(new_n610), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n875), .B2(new_n876), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT101), .A4(KEYINPUT41), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n620), .B(new_n834), .ZN(new_n885));
  MUX2_X1   g460(.A(new_n875), .B(new_n884), .S(new_n885), .Z(new_n886));
  AND2_X1   g461(.A1(new_n872), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n872), .A2(new_n886), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g465(.A(new_n889), .B1(G868), .B2(new_n827), .ZN(G331));
  OAI21_X1  g466(.A(KEYINPUT102), .B1(new_n551), .B2(new_n552), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n542), .A2(new_n543), .A3(new_n534), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n543), .B1(new_n542), .B2(new_n534), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(new_n509), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT74), .B1(new_n895), .B2(new_n549), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n892), .A2(G286), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g475(.A(G168), .B(KEYINPUT102), .C1(new_n551), .C2(new_n552), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n900), .A2(new_n834), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n834), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n901), .ZN(new_n906));
  INV_X1    g481(.A(new_n834), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(KEYINPUT103), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n875), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n871), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n884), .B1(new_n903), .B2(new_n902), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT104), .B(new_n875), .C1(new_n905), .C2(new_n909), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n916), .A2(new_n862), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(new_n914), .A3(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n871), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT43), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n905), .A2(new_n909), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n877), .A2(new_n879), .A3(new_n876), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n875), .A2(new_n876), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n875), .A2(new_n925), .A3(new_n876), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n922), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n902), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(new_n875), .A3(new_n908), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n871), .ZN(new_n932));
  AND4_X1   g507(.A1(KEYINPUT43), .A2(new_n932), .A3(new_n916), .A4(new_n862), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n917), .B2(new_n919), .ZN(new_n937));
  AND4_X1   g512(.A1(new_n936), .A2(new_n932), .A3(new_n916), .A4(new_n862), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(G397));
  AND2_X1   g515(.A1(G160), .A2(G40), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n495), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(G1996), .A3(new_n701), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n718), .B(G2067), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n945), .A2(G1996), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n702), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n789), .A2(new_n791), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n953), .A2(new_n954), .B1(G2067), .B2(new_n718), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(new_n946), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n946), .A2(new_n701), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT125), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n958), .B2(KEYINPUT46), .ZN(new_n959));
  XOR2_X1   g534(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n945), .B2(G1996), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n957), .A2(new_n949), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  INV_X1    g538(.A(new_n953), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n789), .B(new_n791), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n946), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT126), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n945), .A2(G290), .A3(G1986), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n969), .B(KEYINPUT127), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT48), .Z(new_n971));
  AOI211_X1 g546(.A(new_n956), .B(new_n963), .C1(new_n968), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  INV_X1    g548(.A(new_n511), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT112), .B(G86), .Z(new_n975));
  OAI21_X1  g550(.A(new_n591), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G1981), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(KEYINPUT49), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT113), .ZN(new_n979));
  NAND2_X1  g554(.A1(G160), .A2(G40), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n943), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n495), .A2(KEYINPUT107), .A3(new_n942), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n973), .A2(new_n977), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n979), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n583), .A2(new_n585), .A3(G1976), .A4(new_n586), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT110), .B(G1976), .Z(new_n994));
  NAND2_X1  g569(.A1(G288), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n982), .A2(new_n983), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n941), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n999), .A2(new_n992), .A3(G8), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n991), .A4(new_n995), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT109), .B1(new_n1000), .B2(new_n991), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n986), .A2(new_n992), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(KEYINPUT52), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n990), .A2(new_n1003), .A3(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n941), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n496), .A2(new_n942), .A3(new_n498), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n944), .B2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1013), .A2(G1971), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n496), .A2(new_n1015), .A3(new_n942), .A4(new_n498), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI221_X1 g594(.A(new_n941), .B1(new_n1015), .B2(new_n998), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1014), .B1(new_n1020), .B2(G2090), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G166), .A2(new_n985), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT55), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT108), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n998), .B2(new_n1015), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n495), .A2(KEYINPUT107), .A3(new_n942), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT107), .B1(new_n495), .B2(new_n942), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1027), .B(new_n1015), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n941), .B(new_n1026), .C1(new_n1028), .C2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1014), .B1(new_n1033), .B2(G2090), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1024), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(G8), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1015), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT108), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1031), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1039), .A2(new_n728), .A3(new_n941), .A4(new_n1026), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n982), .A2(new_n944), .A3(new_n983), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1041), .B(new_n941), .C1(new_n944), .C2(new_n1012), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n711), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(G286), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1009), .A2(new_n1025), .A3(new_n1036), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AND4_X1   g624(.A1(new_n1036), .A2(new_n1008), .A3(new_n990), .A4(new_n1003), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1034), .A2(G8), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1051), .B2(new_n1024), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1009), .A2(G8), .A3(new_n1035), .A4(new_n1034), .ZN(new_n1055));
  INV_X1    g630(.A(new_n990), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G288), .A2(G1976), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT114), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n973), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n986), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G286), .A2(G8), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1063), .B(KEYINPUT121), .Z(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n985), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1064), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1062), .A2(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1045), .A2(KEYINPUT51), .A3(new_n1064), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1068), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n1013), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1033), .B2(new_n771), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1042), .A2(new_n1079), .A3(G2078), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G301), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1070), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1073), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(G301), .A3(new_n1080), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n943), .A2(new_n944), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1079), .A2(G2078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1087), .A2(new_n941), .A3(new_n1010), .A4(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT122), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1077), .B(new_n1090), .C1(new_n771), .C2(new_n1033), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1086), .B(KEYINPUT54), .C1(new_n1091), .C2(G301), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT123), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1090), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1078), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1096), .B2(G171), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n1086), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1078), .A2(G301), .A3(new_n1095), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1081), .B2(G301), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(new_n1094), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n573), .B1(KEYINPUT116), .B2(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(KEYINPUT116), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1106), .B(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1013), .A2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1108), .B(new_n1110), .C1(new_n1020), .C2(new_n777), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1108), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1020), .A2(new_n777), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1110), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1104), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1033), .A2(new_n767), .ZN(new_n1117));
  INV_X1    g692(.A(G2067), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n984), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n610), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1119), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n611), .B(new_n1121), .C1(new_n1033), .C2(new_n767), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT60), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1113), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1033), .B2(new_n767), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1124), .A2(KEYINPUT61), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(KEYINPUT119), .B(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1013), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT58), .B(G1341), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n999), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n558), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT59), .Z(new_n1133));
  AND4_X1   g708(.A1(new_n1116), .A2(new_n1123), .A3(new_n1127), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1120), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT117), .B1(new_n1125), .B2(new_n610), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT118), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1113), .A2(new_n1141), .A3(new_n1114), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1108), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1111), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1100), .B(new_n1103), .C1(new_n1134), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1085), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1050), .A2(new_n1025), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1061), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n600), .B(G1986), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n964), .B(new_n966), .C1(new_n945), .C2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n972), .B1(new_n1148), .B2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g726(.A1(G229), .A2(new_n460), .ZN(new_n1153));
  NOR2_X1   g727(.A1(G401), .A2(G227), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n863), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g729(.A(new_n919), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n862), .ZN(new_n1157));
  OAI21_X1  g731(.A(KEYINPUT43), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n936), .A3(new_n932), .ZN(new_n1159));
  AOI211_X1 g733(.A(new_n1153), .B(new_n1155), .C1(new_n1158), .C2(new_n1159), .ZN(G308));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1161));
  INV_X1    g735(.A(new_n1155), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1162), .ZN(G225));
endmodule


