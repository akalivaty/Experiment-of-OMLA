

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n974), .A2(n724), .ZN(n721) );
  INV_X1 U557 ( .A(n707), .ZN(n736) );
  NOR2_X1 U558 ( .A1(n751), .A2(n750), .ZN(n757) );
  NAND2_X1 U559 ( .A1(G8), .A2(n759), .ZN(n780) );
  NOR2_X2 U560 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NOR2_X1 U561 ( .A1(n727), .A2(n973), .ZN(n712) );
  INV_X1 U562 ( .A(KEYINPUT28), .ZN(n711) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NOR2_X1 U564 ( .A1(n797), .A2(n796), .ZN(n808) );
  NOR2_X1 U565 ( .A1(n539), .A2(n538), .ZN(G160) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n524), .Z(n897) );
  NAND2_X1 U567 ( .A1(G138), .A2(n897), .ZN(n526) );
  INV_X1 U568 ( .A(G2105), .ZN(n528) );
  XNOR2_X1 U569 ( .A(KEYINPUT66), .B(G2104), .ZN(n527) );
  NOR2_X1 U570 ( .A1(n528), .A2(n527), .ZN(n892) );
  NAND2_X1 U571 ( .A1(G126), .A2(n892), .ZN(n525) );
  NAND2_X1 U572 ( .A1(n526), .A2(n525), .ZN(n532) );
  AND2_X2 U573 ( .A1(n528), .A2(n527), .ZN(n895) );
  NAND2_X1 U574 ( .A1(G102), .A2(n895), .ZN(n530) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U576 ( .A1(G114), .A2(n891), .ZN(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n532), .A2(n531), .ZN(G164) );
  NAND2_X1 U579 ( .A1(n891), .A2(G113), .ZN(n535) );
  NAND2_X1 U580 ( .A1(G101), .A2(n895), .ZN(n533) );
  XOR2_X1 U581 ( .A(KEYINPUT23), .B(n533), .Z(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U583 ( .A1(G137), .A2(n897), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G125), .A2(n892), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n647) );
  NAND2_X1 U587 ( .A1(n647), .A2(G89), .ZN(n540) );
  XNOR2_X1 U588 ( .A(n540), .B(KEYINPUT4), .ZN(n543) );
  INV_X1 U589 ( .A(G651), .ZN(n545) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  OR2_X1 U591 ( .A1(n545), .A2(n628), .ZN(n541) );
  XNOR2_X2 U592 ( .A(KEYINPUT67), .B(n541), .ZN(n645) );
  NAND2_X1 U593 ( .A1(G76), .A2(n645), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n544), .ZN(n553) );
  NOR2_X1 U596 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n546), .Z(n651) );
  NAND2_X1 U598 ( .A1(n651), .A2(G63), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT81), .B(n547), .Z(n550) );
  NOR2_X1 U600 ( .A1(G651), .A2(n628), .ZN(n548) );
  XOR2_X1 U601 ( .A(KEYINPUT65), .B(n548), .Z(n654) );
  NAND2_X1 U602 ( .A1(n654), .A2(G51), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U606 ( .A(KEYINPUT7), .B(n554), .ZN(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  NAND2_X1 U611 ( .A1(G94), .A2(G452), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U613 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U615 ( .A(G223), .ZN(n823) );
  NAND2_X1 U616 ( .A1(n823), .A2(G567), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U618 ( .A1(n651), .A2(G56), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT14), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G43), .A2(n654), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n570) );
  XNOR2_X1 U622 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT13), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n645), .A2(G68), .ZN(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT76), .B(n562), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n564) );
  NAND2_X1 U627 ( .A1(G81), .A2(n647), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U630 ( .A(n568), .B(n567), .ZN(n569) );
  NOR2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X2 U632 ( .A(KEYINPUT79), .B(n571), .Z(n986) );
  NAND2_X1 U633 ( .A1(n986), .A2(G860), .ZN(G153) );
  NAND2_X1 U634 ( .A1(G64), .A2(n651), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT72), .B(n572), .Z(n577) );
  NAND2_X1 U636 ( .A1(G77), .A2(n645), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G90), .A2(n647), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  NOR2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n654), .A2(G52), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n579), .A2(n578), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G79), .A2(n645), .ZN(n581) );
  NAND2_X1 U644 ( .A1(G92), .A2(n647), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U646 ( .A1(G66), .A2(n651), .ZN(n583) );
  NAND2_X1 U647 ( .A1(G54), .A2(n654), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT15), .ZN(n974) );
  INV_X1 U651 ( .A(G868), .ZN(n602) );
  NAND2_X1 U652 ( .A1(n974), .A2(n602), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT80), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G65), .A2(n651), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G53), .A2(n654), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U659 ( .A(KEYINPUT74), .B(n592), .Z(n596) );
  NAND2_X1 U660 ( .A1(G78), .A2(n645), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G91), .A2(n647), .ZN(n593) );
  AND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U664 ( .A1(G286), .A2(n602), .ZN(n598) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(G297) );
  INV_X1 U667 ( .A(G860), .ZN(n617) );
  NAND2_X1 U668 ( .A1(n617), .A2(G559), .ZN(n599) );
  INV_X1 U669 ( .A(n974), .ZN(n615) );
  NAND2_X1 U670 ( .A1(n599), .A2(n615), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G559), .A2(n974), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n604) );
  NOR2_X1 U674 ( .A1(n986), .A2(G868), .ZN(n603) );
  OR2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G111), .A2(n891), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G135), .A2(n897), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n611) );
  NAND2_X1 U679 ( .A1(G123), .A2(n892), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n895), .A2(G99), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n925) );
  XNOR2_X1 U684 ( .A(n925), .B(G2096), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT82), .ZN(n614) );
  INV_X1 U686 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U688 ( .A1(G559), .A2(n615), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(n986), .ZN(n665) );
  NAND2_X1 U690 ( .A1(n617), .A2(n665), .ZN(n624) );
  NAND2_X1 U691 ( .A1(G67), .A2(n651), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G55), .A2(n654), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G80), .A2(n645), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G93), .A2(n647), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n667) );
  XOR2_X1 U698 ( .A(n624), .B(n667), .Z(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n654), .ZN(n626) );
  NAND2_X1 U700 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n651), .A2(n627), .ZN(n630) );
  NAND2_X1 U703 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G62), .A2(n651), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G50), .A2(n654), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G75), .A2(n645), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G88), .A2(n647), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U712 ( .A(KEYINPUT83), .B(n637), .Z(G166) );
  NAND2_X1 U713 ( .A1(G48), .A2(n654), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G86), .A2(n647), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U716 ( .A1(G73), .A2(n645), .ZN(n640) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n651), .A2(G61), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U721 ( .A1(n645), .A2(G72), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(KEYINPUT68), .ZN(n649) );
  NAND2_X1 U723 ( .A1(G85), .A2(n647), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT69), .ZN(n653) );
  NAND2_X1 U726 ( .A1(G60), .A2(n651), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n654), .A2(G47), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT70), .B(n655), .Z(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT71), .B(n658), .ZN(G290) );
  XNOR2_X1 U732 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U733 ( .A(G288), .B(G166), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n667), .B(n661), .ZN(n663) );
  INV_X1 U736 ( .A(G299), .ZN(n973) );
  XNOR2_X1 U737 ( .A(G305), .B(n973), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n663), .B(n662), .ZN(n664) );
  XOR2_X1 U739 ( .A(n664), .B(G290), .Z(n908) );
  XNOR2_X1 U740 ( .A(n908), .B(n665), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n666), .A2(G868), .ZN(n669) );
  OR2_X1 U742 ( .A1(G868), .A2(n667), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n671), .ZN(n673) );
  XOR2_X1 U747 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n672) );
  XNOR2_X1 U748 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G2072), .A2(n674), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n675) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n675), .Z(n676) );
  NOR2_X1 U753 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G96), .A2(n677), .ZN(n827) );
  AND2_X1 U755 ( .A1(G2106), .A2(n827), .ZN(n682) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U757 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G108), .A2(n679), .ZN(n828) );
  NAND2_X1 U759 ( .A1(G567), .A2(n828), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT86), .B(n680), .Z(n681) );
  NOR2_X1 U761 ( .A1(n682), .A2(n681), .ZN(G319) );
  INV_X1 U762 ( .A(G319), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n683) );
  XOR2_X1 U764 ( .A(KEYINPUT87), .B(n683), .Z(n684) );
  NOR2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n826) );
  NAND2_X1 U766 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G166), .ZN(G303) );
  INV_X1 U768 ( .A(G301), .ZN(G171) );
  NAND2_X1 U769 ( .A1(G107), .A2(n891), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G131), .A2(n897), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U772 ( .A1(G95), .A2(n895), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G119), .A2(n892), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n690) );
  OR2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n876) );
  AND2_X1 U776 ( .A1(n876), .A2(G1991), .ZN(n700) );
  NAND2_X1 U777 ( .A1(G117), .A2(n891), .ZN(n693) );
  NAND2_X1 U778 ( .A1(G141), .A2(n897), .ZN(n692) );
  NAND2_X1 U779 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n895), .A2(G105), .ZN(n694) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n694), .Z(n695) );
  NOR2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U783 ( .A1(n892), .A2(G129), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n874) );
  AND2_X1 U785 ( .A1(n874), .A2(G1996), .ZN(n699) );
  NOR2_X1 U786 ( .A1(n700), .A2(n699), .ZN(n922) );
  NAND2_X1 U787 ( .A1(G160), .A2(G40), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n819) );
  INV_X1 U789 ( .A(n819), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n922), .A2(n701), .ZN(n811) );
  INV_X1 U791 ( .A(n811), .ZN(n794) );
  INV_X1 U792 ( .A(n702), .ZN(n704) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n707) );
  BUF_X2 U794 ( .A(n707), .Z(n759) );
  NOR2_X1 U795 ( .A1(G2090), .A2(G303), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n705), .B(KEYINPUT100), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n706), .A2(G8), .ZN(n769) );
  NOR2_X1 U798 ( .A1(G1966), .A2(n780), .ZN(n752) );
  XOR2_X1 U799 ( .A(n736), .B(KEYINPUT90), .Z(n735) );
  INV_X1 U800 ( .A(n735), .ZN(n718) );
  NAND2_X1 U801 ( .A1(G2072), .A2(n718), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U803 ( .A(G1956), .B(KEYINPUT93), .ZN(n1002) );
  NOR2_X1 U804 ( .A1(n718), .A2(n1002), .ZN(n709) );
  NOR2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n727) );
  XNOR2_X1 U806 ( .A(n712), .B(n711), .ZN(n731) );
  AND2_X1 U807 ( .A1(n736), .A2(G1996), .ZN(n714) );
  XOR2_X1 U808 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n713) );
  XNOR2_X1 U809 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n759), .A2(G1341), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n723) );
  NAND2_X1 U812 ( .A1(G1348), .A2(n759), .ZN(n717) );
  XNOR2_X1 U813 ( .A(n717), .B(KEYINPUT94), .ZN(n720) );
  NAND2_X1 U814 ( .A1(G2067), .A2(n718), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n986), .A2(n721), .ZN(n722) );
  NOR2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U818 ( .A1(n724), .A2(n974), .ZN(n725) );
  NOR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n727), .A2(n973), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n733) );
  XOR2_X1 U823 ( .A(KEYINPUT95), .B(KEYINPUT29), .Z(n732) );
  XNOR2_X1 U824 ( .A(n733), .B(n732), .ZN(n741) );
  XNOR2_X1 U825 ( .A(G2078), .B(KEYINPUT25), .ZN(n734) );
  XNOR2_X1 U826 ( .A(n734), .B(KEYINPUT91), .ZN(n949) );
  NOR2_X1 U827 ( .A1(n949), .A2(n735), .ZN(n738) );
  NOR2_X1 U828 ( .A1(n736), .A2(G1961), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U830 ( .A(KEYINPUT92), .B(n739), .Z(n742) );
  AND2_X1 U831 ( .A1(n742), .A2(G171), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n751) );
  NOR2_X1 U833 ( .A1(G171), .A2(n742), .ZN(n747) );
  NOR2_X1 U834 ( .A1(G2084), .A2(n759), .ZN(n753) );
  NOR2_X1 U835 ( .A1(n752), .A2(n753), .ZN(n743) );
  NAND2_X1 U836 ( .A1(G8), .A2(n743), .ZN(n744) );
  XNOR2_X1 U837 ( .A(KEYINPUT30), .B(n744), .ZN(n745) );
  NOR2_X1 U838 ( .A1(G168), .A2(n745), .ZN(n746) );
  NOR2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U840 ( .A(KEYINPUT96), .B(n748), .ZN(n749) );
  XNOR2_X1 U841 ( .A(KEYINPUT31), .B(n749), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n752), .A2(n757), .ZN(n755) );
  NAND2_X1 U843 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U845 ( .A(KEYINPUT97), .B(n756), .Z(n768) );
  INV_X1 U846 ( .A(n757), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n758), .A2(G286), .ZN(n764) );
  NOR2_X1 U848 ( .A1(G1971), .A2(n780), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G303), .A2(n762), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(G8), .ZN(n766) );
  XNOR2_X1 U854 ( .A(n766), .B(KEYINPUT32), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n775) );
  NAND2_X1 U856 ( .A1(n769), .A2(n775), .ZN(n770) );
  NAND2_X1 U857 ( .A1(n780), .A2(n770), .ZN(n771) );
  XOR2_X1 U858 ( .A(KEYINPUT101), .B(n771), .Z(n792) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U860 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U861 ( .A1(n780), .A2(n773), .ZN(n790) );
  XNOR2_X1 U862 ( .A(G1981), .B(G305), .ZN(n969) );
  NOR2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G1971), .A2(G303), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n781), .A2(n774), .ZN(n977) );
  NAND2_X1 U866 ( .A1(n775), .A2(n977), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G288), .A2(G1976), .ZN(n776) );
  XOR2_X1 U868 ( .A(KEYINPUT98), .B(n776), .Z(n972) );
  NOR2_X1 U869 ( .A1(n972), .A2(n780), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  INV_X1 U871 ( .A(KEYINPUT33), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n779), .A2(n784), .ZN(n787) );
  INV_X1 U873 ( .A(n780), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U876 ( .A(n785), .B(KEYINPUT99), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U878 ( .A1(n969), .A2(n788), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n797) );
  XNOR2_X1 U882 ( .A(G1986), .B(G290), .ZN(n984) );
  NAND2_X1 U883 ( .A1(n984), .A2(n819), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(n795), .Z(n796) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NAND2_X1 U886 ( .A1(G104), .A2(n895), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G140), .A2(n897), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n800), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G116), .A2(n891), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G128), .A2(n892), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U893 ( .A(n803), .B(KEYINPUT35), .Z(n804) );
  NOR2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U895 ( .A(KEYINPUT36), .B(n806), .Z(n807) );
  XNOR2_X1 U896 ( .A(KEYINPUT89), .B(n807), .ZN(n871) );
  NOR2_X1 U897 ( .A1(n816), .A2(n871), .ZN(n932) );
  NAND2_X1 U898 ( .A1(n819), .A2(n932), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n808), .A2(n814), .ZN(n821) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n874), .ZN(n920) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n876), .ZN(n924) );
  NOR2_X1 U903 ( .A1(n809), .A2(n924), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n920), .A2(n812), .ZN(n813) );
  XNOR2_X1 U906 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n816), .A2(n871), .ZN(n934) );
  NAND2_X1 U909 ( .A1(n817), .A2(n934), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U912 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U916 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G69), .ZN(G235) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U924 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U925 ( .A(G2454), .B(G2451), .ZN(n838) );
  XNOR2_X1 U926 ( .A(G2430), .B(G2446), .ZN(n836) );
  XOR2_X1 U927 ( .A(G2435), .B(G2427), .Z(n831) );
  XNOR2_X1 U928 ( .A(KEYINPUT102), .B(G2438), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U930 ( .A(n832), .B(G2443), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1348), .B(G1341), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U933 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n839), .A2(G14), .ZN(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT103), .B(n840), .ZN(n915) );
  XNOR2_X1 U937 ( .A(n915), .B(KEYINPUT104), .ZN(G401) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2090), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2067), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1986), .B(G1956), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1971), .B(G1961), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n860) );
  XOR2_X1 U950 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1996), .B(KEYINPUT41), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(G1991), .B(G1966), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1981), .B(G1976), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2474), .B(KEYINPUT106), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U960 ( .A1(n892), .A2(G124), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G136), .A2(n897), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT109), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G100), .A2(n895), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n891), .A2(G112), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT110), .B(n867), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U970 ( .A(G160), .B(n925), .Z(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n880) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n878) );
  XOR2_X1 U976 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(n880), .B(n879), .Z(n890) );
  NAND2_X1 U979 ( .A1(G103), .A2(n895), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G139), .A2(n897), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G115), .A2(n891), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G127), .A2(n892), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT113), .B(n888), .Z(n936) );
  XNOR2_X1 U988 ( .A(n936), .B(G162), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U990 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U993 ( .A1(n895), .A2(G106), .ZN(n896) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n896), .Z(n899) );
  NAND2_X1 U995 ( .A1(n897), .A2(G142), .ZN(n898) );
  NAND2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT45), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n974), .B(G286), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(G171), .B(n986), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n910), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(n913), .A2(G319), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT116), .B(n916), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1013 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n921), .Z(n930) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n928) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT117), .B(n926), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1025 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1026 ( .A(n933), .B(KEYINPUT118), .ZN(n935) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n941) );
  XOR2_X1 U1028 ( .A(G2072), .B(n936), .Z(n938) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n937) );
  NOR2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n939), .Z(n940) );
  NOR2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n942), .ZN(n944) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n945), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1037 ( .A(G29), .B(KEYINPUT121), .ZN(n966) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n956) );
  XOR2_X1 U1041 ( .A(G2072), .B(G33), .Z(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(n949), .B(G27), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(G32), .B(G1996), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n952), .B(KEYINPUT119), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n957), .ZN(n961) );
  XOR2_X1 U1050 ( .A(G34), .B(KEYINPUT120), .Z(n959) );
  XNOR2_X1 U1051 ( .A(G2084), .B(KEYINPUT54), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(n959), .B(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1054 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n964), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(G11), .A2(n967), .ZN(n1023) );
  XNOR2_X1 U1059 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XOR2_X1 U1060 ( .A(G1966), .B(G168), .Z(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT57), .B(n970), .Z(n990) );
  AND2_X1 U1063 ( .A1(G303), .A2(G1971), .ZN(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n982) );
  XNOR2_X1 U1065 ( .A(n973), .B(G1956), .ZN(n976) );
  XOR2_X1 U1066 ( .A(G1348), .B(n974), .Z(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1073 ( .A(KEYINPUT122), .B(n985), .Z(n988) );
  XOR2_X1 U1074 ( .A(n986), .B(G1341), .Z(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n1021) );
  INV_X1 U1078 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1079 ( .A(G1981), .B(G6), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n993), .B(KEYINPUT124), .ZN(n996) );
  XOR2_X1 U1081 ( .A(G1341), .B(G19), .Z(n994) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n994), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1084 ( .A(KEYINPUT125), .B(n997), .Z(n1001) );
  XNOR2_X1 U1085 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(n998), .B(G4), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1348), .B(n999), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(G20), .B(n1002), .Z(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G24), .B(G1986), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G1976), .B(G23), .Z(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1026), .B(KEYINPUT127), .ZN(n1027) );
  XNOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

