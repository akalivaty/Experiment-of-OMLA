//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G146), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G110), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT23), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n192), .A2(new_n195), .A3(KEYINPUT23), .A4(G119), .ZN(new_n200));
  AND4_X1   g014(.A1(new_n191), .A2(new_n197), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n196), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT76), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n196), .A3(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT24), .A2(G110), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT24), .A2(G110), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(KEYINPUT77), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n210));
  INV_X1    g024(.A(new_n208), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n211), .B2(new_n206), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n203), .A2(new_n205), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n190), .B1(new_n201), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT79), .A2(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT79), .A2(G125), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G140), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(G125), .A2(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n223));
  INV_X1    g037(.A(G140), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n220), .A2(G146), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n187), .B1(new_n214), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G146), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n223), .B1(new_n217), .B2(new_n218), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n221), .A2(KEYINPUT16), .A3(G140), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n203), .A2(new_n205), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n209), .A2(new_n212), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G110), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n234), .A2(new_n235), .B1(G110), .B2(new_n237), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(KEYINPUT80), .A3(new_n190), .A4(new_n226), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n228), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(G221), .A2(G234), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT22), .B1(new_n243), .B2(G953), .ZN(new_n244));
  OR3_X1    g058(.A1(new_n243), .A2(KEYINPUT22), .A3(G953), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n244), .A2(G137), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(G137), .B1(new_n245), .B2(new_n244), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT75), .B(G902), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n228), .A2(new_n239), .A3(new_n241), .A4(new_n248), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT25), .ZN(new_n255));
  INV_X1    g069(.A(G217), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(new_n252), .B2(G234), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(new_n258), .A3(new_n252), .A4(new_n253), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT81), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n255), .A2(new_n262), .A3(new_n257), .A4(new_n259), .ZN(new_n263));
  INV_X1    g077(.A(new_n250), .ZN(new_n264));
  INV_X1    g078(.A(new_n253), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT82), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n257), .A2(G902), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n250), .A2(new_n268), .A3(new_n253), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n261), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT0), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n195), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n229), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT64), .A2(G146), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n229), .A2(G143), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n273), .A2(new_n195), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n229), .A2(G143), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n188), .B2(G143), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n281), .A2(new_n282), .B1(new_n284), .B2(new_n274), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT65), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT11), .ZN(new_n288));
  INV_X1    g102(.A(G137), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .A4(G134), .ZN(new_n290));
  INV_X1    g104(.A(G134), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n291), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n291), .A2(G137), .B1(KEYINPUT65), .B2(KEYINPUT11), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n286), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n286), .A3(new_n294), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n285), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n291), .A2(G137), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT66), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n289), .B2(G134), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n300), .B(G131), .C1(new_n299), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT67), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT67), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n296), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(KEYINPUT64), .A2(G146), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT64), .A2(G146), .ZN(new_n310));
  OAI21_X1  g124(.A(G143), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n283), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n313), .A2(KEYINPUT1), .A3(new_n195), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n277), .B1(new_n276), .B2(new_n278), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT68), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n318), .A3(KEYINPUT1), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(G128), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n279), .A2(new_n280), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n314), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n298), .B1(new_n308), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT69), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n324), .B1(new_n325), .B2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n198), .A2(KEYINPUT69), .A3(G116), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT2), .B(G113), .Z(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n331), .B(new_n298), .C1(new_n322), .C2(new_n304), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n272), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n298), .B1(new_n322), .B2(new_n304), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n338), .B(new_n298), .C1(new_n322), .C2(new_n304), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n272), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT26), .B(G101), .Z(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G210), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n342), .B(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT72), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n272), .ZN(new_n350));
  INV_X1    g164(.A(new_n307), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n306), .B1(new_n296), .B2(new_n303), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n319), .A2(G128), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n318), .B1(new_n311), .B2(KEYINPUT1), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n321), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n284), .A2(new_n316), .A3(G128), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n331), .B1(new_n359), .B2(new_n298), .ZN(new_n360));
  INV_X1    g174(.A(new_n334), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT28), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(new_n347), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT30), .B(new_n298), .C1(new_n322), .C2(new_n304), .ZN(new_n366));
  INV_X1    g180(.A(new_n323), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n332), .B(new_n366), .C1(new_n367), .C2(KEYINPUT30), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n334), .A3(new_n348), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT31), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n368), .A2(KEYINPUT31), .A3(new_n334), .A4(new_n348), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n349), .A2(new_n365), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(G472), .A2(G902), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT32), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n364), .B1(new_n363), .B2(new_n347), .ZN(new_n378));
  AOI211_X1 g192(.A(KEYINPUT72), .B(new_n348), .C1(new_n350), .C2(new_n362), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT32), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n374), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n336), .A2(new_n332), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n336), .A2(new_n386), .A3(new_n332), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n334), .B(KEYINPUT73), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n272), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(KEYINPUT29), .A3(new_n348), .A4(new_n350), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n368), .A2(new_n334), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n347), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n394), .B(new_n395), .C1(new_n347), .C2(new_n363), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n252), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G472), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n271), .B1(new_n383), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n322), .A2(new_n221), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n281), .A2(new_n282), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n284), .A2(new_n274), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n222), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT7), .ZN(new_n409));
  INV_X1    g223(.A(G224), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G953), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G110), .B(G122), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT8), .Z(new_n414));
  INV_X1    g228(.A(G113), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n325), .A2(G119), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n329), .B2(new_n416), .ZN(new_n419));
  INV_X1    g233(.A(new_n329), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n330), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G104), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G107), .ZN(new_n424));
  INV_X1    g238(.A(G107), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G104), .ZN(new_n426));
  OAI21_X1  g240(.A(G101), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT3), .B1(new_n423), .B2(G107), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n425), .B2(G104), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n425), .A3(G104), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n423), .A2(KEYINPUT84), .A3(G107), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n427), .B1(new_n434), .B2(G101), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n414), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n439), .A2(new_n418), .B1(new_n330), .B2(new_n420), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n436), .B1(new_n440), .B2(new_n435), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT88), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n406), .B2(new_n222), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n285), .A2(KEYINPUT88), .A3(new_n221), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n411), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(KEYINPUT7), .A3(new_n446), .A4(new_n403), .ZN(new_n447));
  INV_X1    g261(.A(new_n435), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n422), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n428), .A2(new_n432), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n430), .A2(new_n433), .ZN(new_n451));
  INV_X1    g265(.A(G101), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n434), .A2(G101), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(KEYINPUT4), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n434), .A2(new_n456), .A3(G101), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n332), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n458), .A3(new_n413), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n412), .A2(new_n441), .A3(new_n447), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n449), .A2(new_n458), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n413), .B(KEYINPUT87), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT6), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n463), .B1(new_n465), .B2(KEYINPUT6), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n407), .A2(KEYINPUT88), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n406), .A2(new_n442), .A3(new_n222), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n403), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n411), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n446), .B1(new_n445), .B2(new_n403), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n402), .B(new_n460), .C1(new_n466), .C2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(KEYINPUT90), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n464), .B2(new_n459), .ZN(new_n478));
  OAI22_X1  g292(.A1(new_n478), .A2(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n402), .A3(new_n480), .A4(new_n460), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n401), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT94), .Z(new_n484));
  XNOR2_X1  g298(.A(G113), .B(G122), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n423), .ZN(new_n486));
  INV_X1    g300(.A(G237), .ZN(new_n487));
  INV_X1    g301(.A(G953), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(G214), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n277), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n286), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(G131), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n286), .A4(new_n491), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT93), .B1(new_n189), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n219), .B2(new_n500), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n217), .A2(KEYINPUT93), .A3(KEYINPUT19), .A4(new_n218), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n188), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT92), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n494), .A2(new_n496), .A3(new_n506), .A4(new_n497), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n499), .A2(new_n505), .A3(new_n226), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n495), .B(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n190), .B1(new_n219), .B2(new_n229), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n486), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n494), .A2(new_n496), .A3(new_n514), .A4(new_n497), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n495), .A2(KEYINPUT17), .A3(G131), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(new_n232), .A3(new_n226), .A4(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n517), .A2(new_n512), .A3(new_n486), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n484), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT20), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT20), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(new_n484), .C1(new_n513), .C2(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n486), .B1(new_n517), .B2(new_n512), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n402), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n520), .A2(new_n522), .B1(new_n524), .B2(G475), .ZN(new_n525));
  INV_X1    g339(.A(G952), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n526), .A2(G953), .ZN(new_n527));
  NAND2_X1  g341(.A1(G234), .A2(G237), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n251), .A2(G953), .A3(new_n528), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT21), .B(G898), .Z(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT9), .B(G234), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n533), .A2(new_n256), .A3(G953), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n277), .A2(G128), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n277), .A2(G128), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n195), .B2(G143), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n277), .A2(KEYINPUT95), .A3(KEYINPUT13), .A4(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G134), .ZN(new_n543));
  XNOR2_X1  g357(.A(G128), .B(G143), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n291), .ZN(new_n545));
  XNOR2_X1  g359(.A(G116), .B(G122), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(new_n425), .ZN(new_n547));
  INV_X1    g361(.A(new_n546), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G107), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n543), .B(new_n545), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n544), .B(new_n291), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n325), .A2(KEYINPUT14), .A3(G122), .ZN(new_n552));
  OAI211_X1 g366(.A(G107), .B(new_n552), .C1(new_n548), .C2(KEYINPUT14), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n553), .C1(G107), .C2(new_n548), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n534), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n554), .A3(new_n534), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n252), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n559), .A2(new_n561), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n525), .A2(new_n532), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G221), .B1(new_n533), .B2(G902), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT83), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G469), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n356), .A2(new_n357), .A3(new_n435), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT1), .B1(new_n277), .B2(G146), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT85), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT85), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n280), .A2(new_n573), .A3(KEYINPUT1), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(G128), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n313), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n357), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n448), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n570), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n297), .A2(new_n295), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT12), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n583), .B(new_n580), .C1(new_n570), .C2(new_n578), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n358), .A2(KEYINPUT10), .A3(new_n448), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n455), .A2(new_n285), .A3(new_n457), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n586), .A2(new_n580), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n488), .A2(G227), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n322), .A2(new_n587), .A3(new_n435), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n435), .B1(new_n576), .B2(new_n357), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n589), .B1(KEYINPUT10), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n581), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n599), .B2(new_n590), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n569), .B(new_n252), .C1(new_n595), .C2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n593), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n596), .A2(new_n598), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n580), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n599), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n597), .B1(new_n322), .B2(new_n435), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n583), .B1(new_n606), .B2(new_n580), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n579), .A2(KEYINPUT12), .A3(new_n581), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n609), .A2(new_n590), .ZN(new_n610));
  OAI211_X1 g424(.A(G469), .B(new_n605), .C1(new_n610), .C2(new_n593), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n569), .A2(new_n402), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n601), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n482), .A2(new_n565), .A3(new_n568), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n399), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  AND2_X1   g432(.A1(new_n482), .A2(new_n532), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n558), .A2(new_n560), .A3(new_n252), .ZN(new_n621));
  INV_X1    g435(.A(new_n557), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT33), .B1(new_n622), .B2(new_n555), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n556), .A2(new_n624), .A3(new_n557), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n251), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n621), .B1(new_n626), .B2(new_n560), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n525), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n380), .B2(new_n252), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n349), .A2(new_n365), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n375), .B1(new_n633), .B2(new_n377), .ZN(new_n634));
  INV_X1    g448(.A(new_n614), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n271), .A2(new_n567), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n630), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT96), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n638), .B(new_n640), .ZN(G6));
  OR2_X1    g455(.A1(new_n520), .A2(KEYINPUT97), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n524), .A2(G475), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n520), .A2(KEYINPUT97), .A3(new_n522), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n564), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n620), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n636), .A3(new_n637), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  OR3_X1    g465(.A1(new_n246), .A2(KEYINPUT36), .A3(new_n247), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(new_n239), .A3(new_n228), .A4(new_n241), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n652), .B(KEYINPUT98), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n242), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n657), .A3(new_n267), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n261), .A2(new_n659), .A3(new_n263), .ZN(new_n660));
  NOR4_X1   g474(.A1(new_n615), .A2(new_n632), .A3(new_n634), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT37), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G110), .ZN(G12));
  INV_X1    g477(.A(new_n382), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n381), .B1(new_n380), .B2(new_n374), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n398), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n482), .A2(new_n568), .A3(new_n614), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n530), .A2(G900), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT100), .Z(new_n669));
  XOR2_X1   g483(.A(new_n529), .B(KEYINPUT101), .Z(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n667), .A2(new_n647), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n660), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XOR2_X1   g491(.A(new_n672), .B(KEYINPUT39), .Z(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n614), .A2(new_n568), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT40), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n520), .A2(new_n522), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n643), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n646), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n675), .A2(new_n401), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n476), .A2(new_n481), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n389), .A2(new_n387), .A3(new_n385), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n347), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(G472), .A3(new_n369), .ZN(new_n690));
  NAND2_X1  g504(.A1(G472), .A2(G902), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n690), .A2(KEYINPUT102), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT102), .B1(new_n690), .B2(new_n691), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n664), .B2(new_n665), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n681), .A2(new_n685), .A3(new_n687), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  INV_X1    g511(.A(new_n627), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n683), .A2(new_n698), .A3(new_n672), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n628), .A2(KEYINPUT103), .A3(new_n672), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n667), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n666), .A2(new_n704), .A3(new_n675), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n599), .A2(new_n590), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n609), .A2(new_n604), .B1(new_n707), .B2(new_n602), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n708), .B2(new_n251), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n568), .A3(new_n601), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n601), .A3(KEYINPUT104), .A4(new_n568), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n399), .A2(new_n630), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT41), .B(G113), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND3_X1  g531(.A1(new_n399), .A2(new_n648), .A3(new_n714), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G116), .ZN(G18));
  NAND3_X1  g533(.A1(new_n712), .A2(new_n482), .A3(new_n713), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n712), .A2(KEYINPUT105), .A3(new_n482), .A4(new_n713), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n660), .B1(new_n383), .B2(new_n398), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n565), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  XOR2_X1   g541(.A(KEYINPUT106), .B(G472), .Z(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n380), .B2(new_n252), .ZN(new_n729));
  INV_X1    g543(.A(new_n350), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n347), .B1(new_n390), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n375), .B1(new_n731), .B2(new_n377), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n729), .A2(new_n271), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n684), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n619), .A3(new_n734), .A4(new_n714), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR4_X1   g550(.A1(new_n703), .A2(new_n729), .A3(new_n660), .A4(new_n732), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NOR2_X1   g553(.A1(new_n686), .A2(new_n401), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n701), .A3(new_n702), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n635), .A2(new_n567), .ZN(new_n742));
  INV_X1    g556(.A(new_n271), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n666), .A2(new_n741), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n399), .A2(KEYINPUT42), .A3(new_n742), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NOR2_X1   g563(.A1(new_n647), .A2(new_n673), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n742), .A2(new_n666), .A3(new_n743), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n740), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n291), .ZN(G36));
  OR2_X1    g568(.A1(new_n610), .A2(new_n593), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n605), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n605), .B1(new_n610), .B2(new_n593), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n569), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n756), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n613), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n613), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n601), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n568), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n683), .A2(KEYINPUT43), .A3(new_n627), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n525), .B(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n698), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n769), .B1(new_n771), .B2(KEYINPUT43), .ZN(new_n772));
  OAI21_X1  g586(.A(G472), .B1(new_n373), .B2(new_n251), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n380), .A2(new_n374), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n660), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT44), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n768), .A2(new_n776), .A3(new_n678), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n772), .A2(KEYINPUT44), .A3(new_n775), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n740), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(KEYINPUT110), .A3(new_n740), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n777), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  INV_X1    g598(.A(new_n666), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n271), .A3(new_n741), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n271), .A4(new_n741), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n768), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n568), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  AND2_X1   g610(.A1(new_n772), .A2(new_n670), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n687), .A2(new_n400), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n714), .A3(new_n733), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n714), .A2(new_n740), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n743), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n529), .A3(new_n695), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n683), .A2(new_n698), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n801), .A2(new_n802), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n797), .A2(new_n803), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n729), .A2(new_n732), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n675), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n797), .A2(new_n733), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n709), .A2(new_n601), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n568), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n740), .B(new_n811), .C1(new_n794), .C2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n805), .A2(new_n628), .ZN(new_n818));
  INV_X1    g632(.A(new_n527), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n815), .B2(new_n816), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n808), .A2(new_n399), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT48), .Z(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n811), .A2(new_n724), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(KEYINPUT115), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n817), .A2(new_n820), .A3(new_n825), .A4(new_n818), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n823), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n734), .A2(new_n482), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n673), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n695), .A2(new_n742), .A3(new_n660), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n738), .A2(new_n676), .A3(new_n705), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT113), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n724), .A2(new_n737), .B1(new_n725), .B2(new_n674), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n705), .A4(new_n834), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n840), .B2(new_n835), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n661), .B1(new_n399), .B2(new_n616), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n629), .B1(new_n564), .B2(new_n683), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n636), .A2(new_n637), .A3(new_n619), .A4(new_n844), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n726), .A2(new_n843), .A3(new_n735), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n666), .A2(new_n564), .A3(new_n645), .A4(new_n672), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n809), .A2(new_n701), .A3(new_n702), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n742), .A3(new_n675), .A4(new_n740), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n746), .A2(new_n747), .B1(new_n751), .B2(new_n740), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n718), .A2(new_n715), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n842), .A2(new_n855), .A3(KEYINPUT114), .A4(KEYINPUT53), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n748), .A2(new_n752), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n843), .A2(new_n726), .A3(new_n735), .A4(new_n845), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n852), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n840), .B1(new_n836), .B2(new_n839), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n850), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n842), .A2(new_n855), .A3(KEYINPUT53), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n831), .B(new_n856), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n863), .A2(new_n864), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT53), .B1(new_n842), .B2(new_n855), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n830), .A2(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT49), .ZN(new_n874));
  INV_X1    g688(.A(new_n812), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n687), .B(new_n695), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n637), .A2(new_n400), .A3(new_n698), .A4(new_n770), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT112), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n876), .B(new_n878), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n873), .A2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n836), .A2(new_n839), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n854), .B1(new_n882), .B2(new_n841), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT114), .B1(new_n883), .B2(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n866), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n856), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n475), .A3(new_n251), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n466), .A2(new_n472), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n479), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT116), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n887), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n887), .B2(new_n888), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n488), .A2(G952), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G51));
  NAND2_X1  g711(.A1(new_n613), .A2(KEYINPUT57), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n613), .A2(KEYINPUT57), .ZN(new_n899));
  INV_X1    g713(.A(new_n868), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n831), .B1(new_n885), .B2(new_n856), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n708), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n856), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n866), .B2(new_n884), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n906), .A2(new_n252), .A3(new_n762), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n896), .B1(new_n904), .B2(new_n907), .ZN(G54));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n252), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n513), .A2(new_n518), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n896), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(new_n911), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G60));
  NAND2_X1  g730(.A1(new_n623), .A2(new_n625), .ZN(new_n917));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n919), .C1(new_n900), .C2(new_n901), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT117), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n872), .A2(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(new_n917), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n896), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n865), .A2(new_n867), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n926), .B2(new_n905), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n868), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(KEYINPUT117), .A3(new_n917), .A4(new_n919), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n922), .A2(new_n925), .A3(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT118), .Z(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n886), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n266), .A2(new_n269), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n896), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n886), .A2(new_n655), .A3(new_n657), .A4(new_n933), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n937), .C1(KEYINPUT119), .C2(KEYINPUT61), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT61), .B1(new_n937), .B2(KEYINPUT119), .ZN(new_n939));
  INV_X1    g753(.A(new_n933), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n935), .B1(new_n906), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n941), .A3(new_n914), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n943), .ZN(G66));
  INV_X1    g758(.A(new_n531), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n945), .B2(new_n410), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n859), .A2(new_n852), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT120), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n466), .B1(G898), .B2(new_n488), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(G69));
  AOI21_X1  g765(.A(new_n488), .B1(G227), .B2(G900), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n795), .A2(new_n783), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n767), .A2(new_n399), .A3(new_n568), .A4(new_n679), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n851), .B1(new_n832), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n837), .A2(new_n705), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n488), .ZN(new_n958));
  MUX2_X1   g772(.A(new_n367), .B(new_n336), .S(KEYINPUT30), .Z(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n504), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(G900), .A2(G953), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n958), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n963), .B2(KEYINPUT124), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n680), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n399), .A2(new_n966), .A3(new_n740), .A4(new_n844), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n953), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n837), .A2(new_n696), .A3(new_n705), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n968), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n488), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n975), .A2(KEYINPUT123), .A3(new_n976), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n965), .B1(new_n982), .B2(new_n963), .ZN(new_n983));
  INV_X1    g797(.A(new_n963), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n984), .B(new_n964), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G72));
  NOR2_X1   g800(.A1(new_n973), .A2(new_n974), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n947), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n691), .B(KEYINPUT63), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT125), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n393), .A3(new_n348), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n369), .A2(KEYINPUT127), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(new_n394), .Z(new_n994));
  NOR2_X1   g808(.A1(new_n994), .A2(new_n989), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n869), .B2(new_n870), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n957), .A2(new_n947), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n393), .B1(new_n997), .B2(new_n990), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n347), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT126), .B1(new_n999), .B2(new_n914), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n999), .A2(KEYINPUT126), .A3(new_n914), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n992), .B(new_n996), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(G57));
endmodule


