//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT71), .B1(new_n468), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT72), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(new_n473), .A3(G125), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n480), .A2(new_n473), .A3(KEYINPUT70), .A4(G125), .ZN(new_n484));
  NAND2_X1  g059(.A1(G113), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n477), .A2(new_n479), .B1(G2105), .B2(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n474), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT73), .Z(new_n493));
  AND4_X1   g068(.A1(G2105), .A2(new_n469), .A3(new_n471), .A4(new_n473), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n490), .B(new_n493), .C1(G124), .C2(new_n494), .ZN(G162));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n494), .B2(G126), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n469), .A2(new_n471), .A3(new_n473), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n480), .A2(new_n473), .ZN(new_n504));
  NOR3_X1   g079(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n499), .A2(new_n507), .A3(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n502), .A2(KEYINPUT4), .B1(new_n504), .B2(new_n505), .ZN(new_n510));
  INV_X1    g085(.A(new_n496), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n511), .B1(G114), .B2(new_n472), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n469), .A2(new_n471), .A3(G2105), .A4(new_n473), .ZN(new_n513));
  INV_X1    g088(.A(G126), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  INV_X1    g100(.A(new_n521), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n524), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G166));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n526), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n529), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n526), .A2(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n540), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n523), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n530), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n533), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(new_n529), .A2(G56), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n523), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n538), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n523), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n541), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n541), .A2(new_n521), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(G651), .B1(new_n577), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  OR3_X1    g155(.A1(new_n531), .A2(KEYINPUT76), .A3(new_n534), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT76), .B1(new_n531), .B2(new_n534), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  NAND2_X1  g158(.A1(new_n577), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n523), .A2(G49), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n527), .B2(new_n528), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n590), .B2(KEYINPUT77), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n577), .A2(G86), .B1(G48), .B2(new_n523), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n523), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(new_n530), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n533), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n530), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n523), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n529), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n533), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n605), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n605), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(new_n610), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n615), .A2(new_n616), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(G868), .B1(new_n628), .B2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g206(.A1(new_n494), .A2(G123), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT81), .Z(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n634), .A2(KEYINPUT82), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(KEYINPUT82), .B2(new_n634), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n474), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n504), .A2(new_n466), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT80), .B(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT16), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n650), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n669), .B2(new_n649), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  OR2_X1    g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n690), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n691), .A2(KEYINPUT20), .A3(new_n690), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n692), .B1(new_n690), .B2(new_n688), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT87), .ZN(new_n698));
  XOR2_X1   g273(.A(G1981), .B(G1986), .Z(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n698), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G33), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT97), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n491), .A2(G139), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n711), .B(new_n712), .C1(new_n472), .C2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT98), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT99), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n714), .B(KEYINPUT98), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT99), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n707), .B1(new_n722), .B2(new_n705), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2072), .ZN(new_n724));
  NAND2_X1  g299(.A1(G160), .A2(G29), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT24), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(G34), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n705), .B1(new_n726), .B2(G34), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT100), .B(G2084), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n517), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n705), .A2(G27), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2078), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n724), .A2(new_n732), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n738), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n738), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n741), .B1(G1961), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n640), .A2(G29), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G28), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n705), .B1(new_n746), .B2(G28), .ZN(new_n748));
  AND2_X1   g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  NOR2_X1   g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n740), .B2(G1966), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n744), .A2(new_n745), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT101), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n705), .A2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n466), .ZN(new_n761));
  INV_X1    g336(.A(G129), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n513), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G141), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n474), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n756), .B1(new_n767), .B2(new_n705), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT27), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1996), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n743), .A2(G1961), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n730), .B2(new_n731), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n753), .A2(new_n754), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n755), .A2(new_n770), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT102), .ZN(new_n776));
  INV_X1    g351(.A(G2072), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n777), .B(new_n707), .C1(new_n722), .C2(new_n705), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n737), .A2(new_n775), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n724), .A2(new_n778), .A3(new_n732), .A4(new_n736), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT102), .B1(new_n780), .B2(new_n774), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n738), .A2(G19), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT93), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n563), .B2(new_n738), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(G1341), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n738), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT103), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n621), .B2(new_n738), .ZN(new_n789));
  INV_X1    g364(.A(G1956), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n705), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n705), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT29), .B(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n705), .A2(G26), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT28), .Z(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n800));
  INV_X1    g375(.A(G140), .ZN(new_n801));
  INV_X1    g376(.A(G128), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n800), .B1(new_n474), .B2(new_n801), .C1(new_n802), .C2(new_n513), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT95), .B(G2067), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n738), .A2(G4), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n617), .B2(new_n738), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT92), .B(G1348), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n810), .B(new_n811), .Z(new_n812));
  NOR4_X1   g387(.A1(new_n792), .A2(new_n796), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n779), .A2(new_n781), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(G6), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G305), .B2(new_n738), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT32), .B(G1981), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT89), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n738), .A2(G23), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n587), .B2(new_n738), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT33), .B(G1976), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT90), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n823), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n738), .A2(G22), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G166), .B2(new_n738), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1971), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n820), .A2(new_n821), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(KEYINPUT34), .ZN(new_n833));
  NOR2_X1   g408(.A1(G16), .A2(G24), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n603), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT88), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n705), .A2(G25), .ZN(new_n838));
  INV_X1    g413(.A(G119), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n472), .A2(G107), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n513), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n491), .B2(G131), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n838), .B1(new_n843), .B2(new_n705), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  XOR2_X1   g420(.A(new_n844), .B(new_n845), .Z(new_n846));
  NOR2_X1   g421(.A1(new_n837), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n833), .A2(KEYINPUT91), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT91), .B1(new_n833), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n832), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(new_n832), .C1(new_n848), .C2(new_n849), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n814), .B1(new_n851), .B2(new_n853), .ZN(G311));
  INV_X1    g429(.A(new_n814), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(G150));
  NAND2_X1  g432(.A1(new_n523), .A2(G55), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(new_n530), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n533), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT105), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n617), .A2(G559), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n864), .B1(new_n561), .B2(new_n562), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n557), .A2(new_n560), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(new_n863), .C1(KEYINPUT75), .C2(new_n556), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n870), .B(new_n874), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g452(.A(G860), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n867), .B1(new_n877), .B2(new_n879), .ZN(G145));
  XNOR2_X1  g455(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n843), .B(KEYINPUT106), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n644), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n491), .A2(G142), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n494), .A2(G130), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n472), .A2(G118), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n885), .B(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n499), .A2(new_n507), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n805), .B(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(new_n767), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n767), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n716), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n721), .B1(new_n897), .B2(new_n896), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n892), .B(new_n893), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n722), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n891), .A3(new_n898), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n640), .B(G160), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(G162), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n898), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n893), .B1(new_n909), .B2(new_n892), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n883), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n891), .A4(new_n898), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n906), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT107), .B1(new_n909), .B2(new_n892), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n882), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(new_n892), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT108), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n918), .A2(new_n904), .A3(new_n907), .A4(new_n901), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n920), .A3(new_n904), .ZN(new_n921));
  INV_X1    g496(.A(new_n913), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n919), .A2(new_n923), .A3(new_n883), .A4(new_n881), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n916), .A2(new_n924), .ZN(G395));
  NAND2_X1  g500(.A1(new_n628), .A2(G299), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n617), .A2(new_n621), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(KEYINPUT110), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n628), .A2(G559), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n874), .B(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT41), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n926), .A2(new_n927), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n929), .A2(KEYINPUT111), .A3(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n587), .B(G166), .Z(new_n943));
  XOR2_X1   g518(.A(new_n603), .B(G305), .Z(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  AND3_X1   g521(.A1(new_n935), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n935), .B2(new_n942), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G868), .B2(new_n863), .ZN(G295));
  OAI21_X1  g525(.A(new_n949), .B1(G868), .B2(new_n863), .ZN(G331));
  XNOR2_X1  g526(.A(G171), .B(KEYINPUT112), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n871), .A2(new_n952), .A3(new_n873), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n871), .B2(new_n873), .ZN(new_n954));
  OAI21_X1  g529(.A(G286), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n874), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n871), .A2(new_n952), .A3(new_n873), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(G168), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(new_n941), .A3(new_n940), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n928), .B2(new_n960), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n945), .ZN(new_n963));
  INV_X1    g538(.A(new_n945), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n961), .B(new_n964), .C1(new_n928), .C2(new_n960), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n930), .A2(new_n931), .A3(new_n955), .A4(new_n959), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n936), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n938), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n960), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n938), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n945), .B(new_n967), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AND4_X1   g548(.A1(KEYINPUT43), .A2(new_n973), .A3(new_n965), .A4(new_n883), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT44), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n963), .B2(new_n965), .ZN(new_n978));
  AND4_X1   g553(.A1(new_n977), .A2(new_n973), .A3(new_n965), .A4(new_n883), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(G397));
  NAND2_X1  g556(.A1(new_n477), .A2(new_n479), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n486), .A2(G2105), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT114), .B(G40), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n510), .B2(new_n515), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2067), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n805), .B(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n766), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n843), .B(new_n845), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1986), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n999), .A3(new_n603), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n766), .B1(KEYINPUT46), .B2(new_n994), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n991), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT46), .B1(new_n991), .B2(new_n994), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT127), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n843), .A2(new_n845), .ZN(new_n1012));
  OAI22_X1  g587(.A1(new_n996), .A2(new_n1012), .B1(G2067), .B2(new_n805), .ZN(new_n1013));
  AOI211_X1 g588(.A(new_n1002), .B(new_n1011), .C1(new_n991), .C2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n581), .A2(new_n582), .A3(G8), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI221_X4 g594(.A(new_n984), .B1(new_n486), .B2(G2105), .C1(new_n477), .C2(new_n479), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n987), .C1(new_n510), .C2(new_n515), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n508), .B2(new_n516), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1020), .B(new_n1021), .C1(new_n1022), .C2(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g598(.A(G1971), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n517), .B2(new_n987), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(new_n987), .C1(new_n510), .C2(new_n515), .ZN(new_n1028));
  NAND3_X1  g603(.A1(G160), .A2(new_n985), .A3(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(new_n1029), .A3(G2090), .ZN(new_n1030));
  OAI211_X1 g605(.A(G8), .B(new_n1019), .C1(new_n1025), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n595), .B2(new_n596), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n595), .A2(new_n596), .A3(new_n1032), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1035), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n1033), .ZN(new_n1039));
  INV_X1    g614(.A(new_n988), .ZN(new_n1040));
  NAND3_X1  g615(.A1(G160), .A2(new_n1040), .A3(new_n985), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT116), .B(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1036), .A2(new_n1039), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n587), .A2(G1976), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(new_n1041), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1044), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1035), .B(KEYINPUT117), .Z(new_n1052));
  NOR2_X1   g627(.A1(G288), .A2(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1055));
  OAI22_X1  g630(.A1(new_n1031), .A2(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1051), .ZN(new_n1058));
  AOI211_X1 g633(.A(KEYINPUT50), .B(G1384), .C1(new_n508), .C2(new_n516), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(G160), .A3(new_n985), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n1059), .A2(new_n1061), .A3(G2090), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1042), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1031), .B(new_n1058), .C1(new_n1019), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1966), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n990), .A2(G160), .A3(KEYINPUT118), .A4(new_n985), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n517), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT118), .B1(new_n1020), .B2(new_n990), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1027), .A2(G2084), .A3(new_n1029), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(G168), .A3(new_n1043), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1057), .B1(new_n1065), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1074), .ZN(new_n1076));
  OAI21_X1  g651(.A(G8), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1019), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1057), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1076), .A2(new_n1079), .A3(new_n1031), .A4(new_n1058), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1056), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(new_n1043), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1073), .B2(new_n1043), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT126), .B(KEYINPUT51), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1073), .A2(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1082), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1073), .A2(G286), .A3(new_n1043), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT62), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1085), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1090), .ZN(new_n1094));
  INV_X1    g669(.A(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1082), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1086), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1093), .B(KEYINPUT62), .C1(new_n1094), .C2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1100));
  AND4_X1   g675(.A1(new_n982), .A2(new_n1028), .A3(new_n983), .A4(new_n985), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(new_n1026), .C2(new_n1022), .ZN(new_n1103));
  INV_X1    g678(.A(G1961), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1023), .B2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  INV_X1    g683(.A(new_n990), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n986), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1106), .A2(G2078), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1068), .A3(new_n1067), .A4(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1065), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1099), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1081), .B1(new_n1092), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1105), .A2(G301), .A3(new_n1107), .A4(new_n1112), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(KEYINPUT54), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1111), .A2(G40), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n990), .A2(G160), .A3(new_n1021), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1105), .A2(new_n1107), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G171), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1065), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1113), .A2(G171), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1122), .A2(G171), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1091), .A3(new_n1128), .ZN(new_n1129));
  AND4_X1   g704(.A1(new_n982), .A2(new_n1021), .A3(new_n983), .A4(new_n985), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1130), .B(new_n994), .C1(KEYINPUT45), .C2(new_n1022), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(G1341), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n986), .B2(new_n988), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1041), .A2(KEYINPUT122), .A3(new_n1133), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n563), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1130), .B(new_n1143), .C1(KEYINPUT45), .C2(new_n1022), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n790), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n573), .B2(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G299), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n573), .B(new_n578), .C1(KEYINPUT119), .C2(KEYINPUT57), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1144), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1144), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1150), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1142), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1100), .A2(new_n1103), .A3(new_n811), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1020), .A2(new_n992), .A3(new_n1040), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n628), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n628), .A2(KEYINPUT124), .A3(new_n1162), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n617), .B2(KEYINPUT60), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1138), .A2(KEYINPUT123), .A3(new_n563), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(KEYINPUT59), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1159), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n628), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1153), .B1(new_n1177), .B2(new_n1157), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1129), .B1(new_n1179), .B2(KEYINPUT125), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(new_n1181), .A3(new_n1178), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1117), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n991), .A2(G1986), .A3(G290), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1000), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT115), .Z(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n998), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1014), .B1(new_n1183), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g763(.A1(G229), .A2(new_n463), .A3(G227), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n667), .B2(new_n670), .ZN(new_n1191));
  OAI21_X1  g765(.A(new_n1191), .B1(new_n911), .B2(new_n915), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n978), .A2(new_n979), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1192), .A2(new_n1193), .ZN(G308));
  OAI221_X1 g768(.A(new_n1191), .B1(new_n911), .B2(new_n915), .C1(new_n978), .C2(new_n979), .ZN(G225));
endmodule


