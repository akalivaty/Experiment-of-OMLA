//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT64), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT65), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT65), .B1(new_n462), .B2(new_n464), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT66), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n460), .ZN(new_n476));
  OAI22_X1  g051(.A1(new_n472), .A2(new_n473), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  OR3_X1    g056(.A1(new_n476), .A2(KEYINPUT67), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(new_n476), .B2(new_n481), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n462), .A2(new_n464), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(new_n460), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n482), .A2(new_n483), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT68), .Z(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n460), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n461), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G102), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n460), .A2(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n484), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n463), .A2(G2104), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT65), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n498), .B(new_n502), .C1(KEYINPUT4), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n511), .B1(KEYINPUT6), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(KEYINPUT69), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n511), .B(G651), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AND2_X1   g097(.A1(G75), .A2(G651), .ZN(new_n523));
  OAI21_X1  g098(.A(G543), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT5), .B(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n521), .A2(G88), .ZN(new_n526));
  AND2_X1   g101(.A1(G62), .A2(G651), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n515), .B2(new_n520), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT71), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(G51), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n521), .A2(G89), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n525), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n533), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n512), .ZN(new_n545));
  INV_X1    g120(.A(new_n525), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n515), .B2(new_n520), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G90), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n543), .A2(new_n545), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n533), .A2(G43), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n512), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n547), .A2(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n547), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n546), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n532), .A2(KEYINPUT9), .A3(G53), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(KEYINPUT73), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT73), .B1(new_n571), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT74), .ZN(G299));
  NAND2_X1  g152(.A1(new_n532), .A2(G49), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n512), .B1(new_n546), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n547), .B2(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n532), .A2(KEYINPUT75), .A3(G49), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n512), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G86), .B2(new_n547), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n532), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n533), .A2(G47), .B1(G85), .B2(new_n547), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n512), .B2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n547), .A2(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n533), .A2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n525), .A2(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n512), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT76), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n604));
  AOI211_X1 g179(.A(new_n604), .B(new_n601), .C1(new_n533), .C2(G54), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n594), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n594), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(new_n568), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n612));
  INV_X1    g187(.A(new_n572), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT9), .B1(new_n532), .B2(G53), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n615), .B2(new_n573), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT74), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G868), .ZN(G297));
  XNOR2_X1  g193(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n607), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n607), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT78), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n476), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n485), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(new_n460), .B2(G111), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT80), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2096), .ZN(new_n634));
  INV_X1    g209(.A(new_n472), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n506), .A2(new_n507), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT13), .B(G2100), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2451), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(G401));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(KEYINPUT82), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT17), .Z(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n659), .B2(new_n658), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n661), .A2(new_n657), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n660), .B1(new_n667), .B2(new_n659), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n663), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2100), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(new_n682), .C2(new_n681), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n685), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT83), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  XOR2_X1   g268(.A(KEYINPUT85), .B(G16), .Z(new_n694));
  MUX2_X1   g269(.A(G24), .B(G290), .S(new_n694), .Z(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT86), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1986), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(KEYINPUT86), .ZN(new_n698));
  INV_X1    g273(.A(G1986), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(new_n460), .B2(G107), .ZN(new_n704));
  INV_X1    g279(.A(G95), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n460), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT84), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n485), .A2(G119), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n627), .A2(G131), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(G29), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n701), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n694), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT88), .B(G1971), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G6), .B(G305), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT87), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G288), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G16), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT33), .ZN(new_n729));
  OR2_X1    g304(.A1(G16), .A2(G23), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1976), .ZN(new_n734));
  INV_X1    g309(.A(G1976), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n731), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n722), .B(new_n726), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT34), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n717), .A2(new_n739), .A3(KEYINPUT89), .A4(KEYINPUT36), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n741));
  OR2_X1    g316(.A1(KEYINPUT89), .A2(KEYINPUT36), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n701), .A2(new_n715), .A3(new_n716), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n738), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n495), .A2(G103), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT91), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n627), .A2(G139), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n636), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n749), .B(new_n750), .C1(new_n460), .C2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n702), .ZN(new_n754));
  INV_X1    g329(.A(G33), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT93), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n758));
  INV_X1    g333(.A(new_n756), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n758), .B(new_n759), .C1(new_n753), .C2(new_n702), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n633), .A2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(G171), .A2(G16), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G5), .B2(G16), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  OR2_X1    g346(.A1(G29), .A2(G32), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n485), .A2(G129), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n627), .A2(G141), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n773), .B(new_n774), .C1(G105), .C2(new_n635), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT26), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n779), .B2(new_n702), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n627), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G128), .ZN(new_n786));
  NOR2_X1   g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n460), .B2(G116), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G29), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n702), .A2(G26), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2067), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G28), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n797), .A2(KEYINPUT98), .A3(KEYINPUT30), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(KEYINPUT30), .ZN(new_n799));
  OAI21_X1  g374(.A(KEYINPUT98), .B1(new_n797), .B2(KEYINPUT30), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n771), .A2(new_n784), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n763), .A2(new_n764), .A3(new_n770), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n780), .A2(new_n783), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n761), .A2(new_n762), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n702), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n702), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(G2090), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n807), .A2(new_n808), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n806), .A2(KEYINPUT94), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n718), .A2(G20), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G16), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n617), .B2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g397(.A1(G168), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G16), .B2(G21), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT97), .B(G1966), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n821), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n805), .A2(new_n814), .A3(new_n815), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n812), .A2(new_n813), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n767), .B2(new_n766), .ZN(new_n831));
  AND2_X1   g406(.A1(KEYINPUT24), .A2(G34), .ZN(new_n832));
  NOR2_X1   g407(.A1(KEYINPUT24), .A2(G34), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G29), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n479), .B2(G29), .ZN(new_n835));
  INV_X1    g410(.A(G2084), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n827), .A2(new_n822), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n556), .A2(new_n718), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G19), .B2(new_n718), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(G1341), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(G1341), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n844), .B(new_n845), .C1(new_n768), .C2(new_n769), .ZN(new_n846));
  NOR4_X1   g421(.A1(new_n829), .A2(new_n839), .A3(new_n840), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n819), .A2(G4), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n607), .B2(new_n819), .ZN(new_n849));
  INV_X1    g424(.A(G1348), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n702), .A2(G27), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G164), .B2(new_n702), .ZN(new_n853));
  INV_X1    g428(.A(G2078), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n746), .A2(new_n847), .A3(new_n851), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n824), .A2(new_n826), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(G311));
  NOR2_X1   g433(.A1(new_n829), .A2(new_n846), .ZN(new_n859));
  INV_X1    g434(.A(new_n839), .ZN(new_n860));
  INV_X1    g435(.A(new_n840), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n745), .ZN(new_n863));
  INV_X1    g438(.A(new_n857), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n851), .A4(new_n855), .ZN(G150));
  AOI22_X1  g440(.A1(new_n533), .A2(G55), .B1(G93), .B2(new_n547), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(new_n512), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n556), .A2(new_n869), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n555), .A2(new_n868), .A3(new_n866), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n606), .A2(new_n620), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n878), .B2(G860), .ZN(G145));
  XNOR2_X1  g454(.A(new_n633), .B(G160), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G162), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n753), .B(new_n789), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT103), .B1(new_n494), .B2(new_n497), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  INV_X1    g459(.A(new_n493), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n475), .B2(G126), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n496), .C1(new_n886), .C2(new_n460), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(G138), .B(new_n460), .C1(new_n465), .C2(new_n466), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n501), .B1(new_n889), .B2(new_n499), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n779), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n882), .B(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n639), .B(new_n710), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n627), .A2(G142), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n485), .A2(G130), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT105), .ZN(new_n898));
  NOR2_X1   g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  OAI21_X1  g474(.A(G2104), .B1(new_n460), .B2(G118), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n896), .B(new_n898), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n894), .B(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n893), .B1(KEYINPUT107), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n882), .B(new_n892), .Z(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n902), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n881), .B(new_n904), .C1(new_n906), .C2(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n893), .A2(KEYINPUT107), .A3(new_n903), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n909), .A2(new_n904), .A3(new_n910), .A4(new_n881), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n906), .A2(KEYINPUT106), .ZN(new_n913));
  INV_X1    g488(.A(new_n881), .ZN(new_n914));
  INV_X1    g489(.A(new_n906), .ZN(new_n915));
  OAI21_X1  g490(.A(KEYINPUT106), .B1(new_n905), .B2(new_n902), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n912), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(G395));
  INV_X1    g497(.A(G868), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n869), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G290), .B(G288), .ZN(new_n925));
  XNOR2_X1  g500(.A(G303), .B(G305), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n925), .B(new_n926), .Z(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n928), .B2(KEYINPUT110), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(KEYINPUT42), .C1(KEYINPUT109), .C2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(KEYINPUT42), .B2(new_n929), .ZN(new_n931));
  NAND2_X1  g506(.A1(G299), .A2(new_n607), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n617), .A2(new_n606), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n622), .B(new_n874), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n934), .B2(new_n937), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n931), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n924), .B1(new_n941), .B2(new_n923), .ZN(G295));
  OAI21_X1  g517(.A(new_n924), .B1(new_n941), .B2(new_n923), .ZN(G331));
  XOR2_X1   g518(.A(G286), .B(G301), .Z(new_n944));
  OR2_X1    g519(.A1(new_n944), .A2(new_n874), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n874), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n936), .A2(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n934), .A3(new_n946), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n927), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n945), .A2(new_n946), .ZN(new_n952));
  INV_X1    g527(.A(new_n938), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT41), .B1(new_n932), .B2(new_n933), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n928), .A3(new_n948), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n950), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n950), .A2(new_n960), .A3(new_n956), .A4(new_n951), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n958), .A2(KEYINPUT111), .A3(new_n961), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n957), .A2(new_n967), .A3(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n969), .ZN(G397));
  OR2_X1    g545(.A1(G290), .A2(G1986), .ZN(new_n971));
  AOI21_X1  g546(.A(G1384), .B1(new_n888), .B2(new_n890), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT113), .B(G40), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n636), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n478), .B(new_n975), .C1(new_n976), .C2(new_n460), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n971), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT48), .Z(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n779), .B(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n789), .B(G2067), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n710), .A2(new_n713), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n710), .A2(new_n713), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n979), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n979), .B2(G1996), .ZN(new_n991));
  INV_X1    g566(.A(new_n984), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n978), .B1(new_n779), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n982), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  INV_X1    g571(.A(new_n987), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n985), .A2(new_n997), .B1(G2067), .B2(new_n789), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n978), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n989), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT127), .Z(new_n1001));
  INV_X1    g576(.A(KEYINPUT126), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n977), .B1(new_n972), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n890), .B2(new_n498), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT114), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n502), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n496), .B1(new_n886), .B2(new_n460), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT50), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1006), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n972), .A2(KEYINPUT45), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n469), .A2(new_n477), .A3(new_n974), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1014), .A2(new_n854), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1013), .A2(new_n767), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n1007), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n509), .A2(KEYINPUT119), .A3(KEYINPUT45), .A4(new_n1007), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1015), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1019), .A2(G2078), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1020), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G171), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n479), .B1(new_n972), .B2(KEYINPUT45), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n973), .A2(new_n1032), .A3(G40), .A4(new_n1028), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(G301), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT54), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n972), .A2(new_n1015), .ZN(new_n1036));
  XOR2_X1   g611(.A(KEYINPUT58), .B(G1341), .Z(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(G1996), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n556), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1042), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n556), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT60), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1036), .A2(G2067), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1046), .B(new_n1047), .C1(new_n1013), .C2(new_n850), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1043), .A2(new_n1045), .B1(new_n1048), .B2(new_n606), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n1013), .B2(new_n850), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n606), .B1(new_n1050), .B2(KEYINPUT60), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1051), .B1(KEYINPUT60), .B2(new_n1050), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n576), .A2(KEYINPUT57), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n568), .A2(new_n1054), .A3(new_n571), .A4(new_n572), .ZN(new_n1055));
  INV_X1    g630(.A(G1956), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n972), .A2(new_n1003), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1015), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1053), .A2(new_n1055), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(KEYINPUT61), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1053), .A2(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(KEYINPUT61), .B2(new_n1062), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1049), .A2(new_n1052), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1013), .A2(new_n850), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n607), .B(KEYINPUT120), .C1(new_n1067), .C2(new_n1047), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1055), .B1(new_n616), .B2(new_n1054), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1053), .A2(KEYINPUT121), .A3(new_n1055), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1050), .B2(new_n606), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1068), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1062), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1035), .B1(new_n1066), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n826), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1004), .A2(new_n1006), .A3(new_n836), .A4(new_n1012), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(G168), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1082), .A2(new_n1088), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT123), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1083), .A2(KEYINPUT124), .A3(new_n1084), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G168), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1020), .A2(G301), .A3(new_n1029), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1020), .B2(new_n1033), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1101), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT54), .A4(new_n1099), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1079), .A2(new_n1098), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1031), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1091), .A2(new_n1089), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT124), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1086), .B(KEYINPUT51), .C1(new_n1082), .C2(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1096), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1093), .A2(new_n1114), .A3(new_n1097), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G8), .ZN(new_n1118));
  NOR3_X1   g693(.A1(G166), .A2(KEYINPUT55), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT55), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(G303), .B2(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1971), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1039), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n977), .B1(new_n1005), .B2(new_n1003), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n813), .C1(new_n1003), .C2(new_n972), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1127), .A3(KEYINPUT117), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT117), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1123), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1125), .B1(G2090), .B2(new_n1013), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(new_n1122), .A3(G8), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT115), .B1(new_n1036), .B2(G8), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1137), .B(new_n1118), .C1(new_n972), .C2(new_n1015), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT49), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G305), .A2(G1981), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(G305), .A2(G1981), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1142), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1139), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g721(.A1(new_n1136), .A2(new_n1138), .B1(new_n735), .B2(G288), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT52), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT52), .B1(G288), .B2(new_n735), .ZN(new_n1149));
  OAI221_X1 g724(.A(new_n1149), .B1(new_n735), .B2(G288), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1150));
  AND4_X1   g725(.A1(new_n1135), .A2(new_n1146), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT118), .B(new_n1123), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1133), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1117), .A2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1095), .A2(G286), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1133), .A2(new_n1151), .A3(new_n1152), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1134), .A2(G8), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1159), .B2(new_n1123), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1151), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1139), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1146), .A2(new_n735), .A3(new_n727), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1164), .B2(new_n1142), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1166), .A2(new_n1135), .ZN(new_n1167));
  OR3_X1    g742(.A1(new_n1165), .A2(new_n1167), .A3(KEYINPUT116), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT116), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1162), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1154), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n988), .A2(new_n971), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(G290), .A2(G1986), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n979), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1002), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1171), .B1(new_n1117), .B2(new_n1153), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1180), .A2(KEYINPUT126), .A3(new_n1177), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1001), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g757(.A1(new_n918), .A2(G319), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G401), .A2(G227), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n965), .A2(new_n692), .A3(new_n968), .A4(new_n1185), .ZN(new_n1186));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1186), .ZN(G308));
  INV_X1    g761(.A(G319), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n912), .B2(new_n917), .ZN(new_n1189));
  AND2_X1   g763(.A1(new_n965), .A2(new_n968), .ZN(new_n1190));
  NAND4_X1  g764(.A1(new_n1189), .A2(new_n1190), .A3(new_n692), .A4(new_n1185), .ZN(G225));
endmodule


