//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  XOR2_X1   g001(.A(G141gat), .B(G148gat), .Z(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n206), .C1(new_n211), .C2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT29), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217));
  INV_X1    g016(.A(G211gat), .ZN(new_n218));
  INV_X1    g017(.A(G218gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT79), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n222), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G211gat), .B(G218gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n228), .A2(new_n221), .A3(new_n223), .A4(new_n224), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT80), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT80), .B1(new_n227), .B2(new_n229), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n216), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT88), .ZN(new_n234));
  INV_X1    g033(.A(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n230), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n216), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n227), .A2(new_n229), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n213), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n212), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n234), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G228gat), .A2(G233gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n231), .B2(new_n232), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(KEYINPUT81), .A3(new_n230), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n216), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n244), .B1(new_n240), .B2(new_n241), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT31), .B(G50gat), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G78gat), .B(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G22gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n255), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n245), .B(new_n259), .C1(new_n252), .C2(new_n253), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n256), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n256), .B2(new_n260), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G127gat), .ZN(new_n267));
  INV_X1    g066(.A(G127gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G113gat), .ZN(new_n271));
  INV_X1    g070(.A(G120gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G113gat), .A2(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI22_X1  g074(.A1(new_n270), .A2(KEYINPUT71), .B1(new_n275), .B2(KEYINPUT1), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(G113gat), .A2(G120gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(G113gat), .A2(G120gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n273), .A2(new_n283), .A3(new_n274), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(KEYINPUT1), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT74), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n279), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n241), .A2(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n214), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n265), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT5), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n270), .A2(KEYINPUT71), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n297), .B(new_n277), .C1(KEYINPUT1), .C2(new_n275), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT74), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT74), .B1(new_n285), .B2(new_n287), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  INV_X1    g103(.A(new_n241), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n298), .B(KEYINPUT75), .C1(new_n299), .C2(new_n300), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT4), .B1(new_n301), .B2(new_n241), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n296), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313));
  AND4_X1   g112(.A1(KEYINPUT4), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n314));
  INV_X1    g113(.A(new_n265), .ZN(new_n315));
  INV_X1    g114(.A(new_n214), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n213), .B1(new_n210), .B2(new_n212), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n318), .B2(new_n301), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n304), .B1(new_n301), .B2(new_n241), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT83), .B1(new_n314), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT4), .B1(new_n292), .B2(new_n305), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n295), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n303), .A2(KEYINPUT4), .A3(new_n305), .A4(new_n306), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n301), .B(new_n305), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT5), .B1(new_n329), .B2(new_n265), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n313), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  AOI211_X1 g131(.A(KEYINPUT84), .B(new_n330), .C1(new_n322), .C2(new_n327), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n312), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT0), .ZN(new_n336));
  XNOR2_X1  g135(.A(G57gat), .B(G85gat), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n334), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT87), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n334), .A2(new_n344), .A3(new_n339), .A4(new_n341), .ZN(new_n345));
  AND4_X1   g144(.A1(new_n325), .A2(new_n326), .A3(new_n319), .A4(new_n320), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n331), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT84), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n313), .A3(new_n331), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n338), .A3(new_n312), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n334), .B2(new_n339), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n343), .A2(new_n345), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  NAND3_X1  g154(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT65), .B(G169gat), .ZN(new_n365));
  INV_X1    g164(.A(G176gat), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n366), .A2(KEYINPUT23), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT23), .ZN(new_n370));
  NOR2_X1   g169(.A1(G169gat), .A2(G176gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n355), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT66), .B(new_n355), .C1(new_n364), .C2(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n356), .ZN(new_n379));
  INV_X1    g178(.A(G169gat), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n355), .B1(new_n367), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n373), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G183gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT28), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n387), .A2(new_n388), .A3(G190gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT27), .B1(new_n360), .B2(KEYINPUT67), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n390), .B(new_n361), .C1(KEYINPUT67), .C2(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT68), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OR3_X1    g192(.A1(new_n360), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(KEYINPUT68), .A3(new_n361), .A4(new_n390), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n393), .A2(KEYINPUT69), .A3(new_n388), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n389), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n372), .A2(KEYINPUT26), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n401), .B(KEYINPUT70), .Z(new_n402));
  OAI21_X1  g201(.A(new_n369), .B1(new_n372), .B2(KEYINPUT26), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n402), .A2(new_n403), .B1(new_n360), .B2(new_n361), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n383), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G226gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  OAI221_X1 g210(.A(new_n383), .B1(new_n406), .B2(new_n407), .C1(new_n400), .C2(new_n404), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n247), .A2(new_n248), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n412), .A3(new_n236), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n418), .B(new_n419), .Z(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n420), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n416), .ZN(new_n427));
  INV_X1    g226(.A(new_n414), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n411), .B2(new_n412), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n420), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n423), .A3(KEYINPUT82), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n264), .B1(new_n354), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n236), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n436), .B1(new_n411), .B2(new_n412), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n438));
  OAI22_X1  g237(.A1(new_n437), .A2(new_n438), .B1(new_n413), .B2(new_n428), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n438), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT37), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n420), .B1(new_n417), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n427), .B2(new_n429), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n415), .A2(KEYINPUT37), .A3(new_n416), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n422), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT38), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n445), .A2(new_n430), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n353), .A2(new_n352), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n338), .B1(new_n351), .B2(new_n312), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n344), .B1(new_n452), .B2(new_n341), .ZN(new_n453));
  INV_X1    g252(.A(new_n345), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n334), .A2(new_n339), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT40), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n310), .A2(new_n311), .B1(new_n292), .B2(new_n294), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT39), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n315), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n338), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n329), .A2(new_n265), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT39), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n463), .B1(new_n458), .B2(new_n315), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n457), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(new_n315), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n329), .B2(new_n265), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n338), .A4(new_n460), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n432), .A2(new_n421), .A3(new_n423), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n456), .A2(new_n465), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n471), .A2(new_n263), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n303), .A2(new_n306), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n405), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n405), .A2(new_n474), .ZN(new_n476));
  OAI211_X1 g275(.A(G227gat), .B(G233gat), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT76), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G227gat), .A2(G233gat), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n400), .A2(new_n404), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n303), .A2(new_n306), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n383), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n405), .A2(new_n474), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT76), .B1(new_n486), .B2(KEYINPUT33), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G43gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(G71gat), .B(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n484), .A2(new_n497), .A3(new_n485), .A4(new_n481), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT78), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n491), .A2(new_n479), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n481), .A3(new_n485), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT34), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT77), .A3(KEYINPUT34), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n496), .A2(new_n499), .A3(new_n503), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n499), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n494), .B1(new_n480), .B2(new_n487), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n502), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n510), .B2(new_n513), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n435), .A2(new_n473), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n519));
  INV_X1    g318(.A(new_n434), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n510), .A2(new_n513), .A3(new_n263), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n343), .A2(new_n345), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n451), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n513), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n526), .A2(new_n264), .A3(new_n470), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n522), .A2(KEYINPUT35), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n518), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT14), .B(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n532), .A2(KEYINPUT15), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT94), .Z(new_n537));
  AND2_X1   g336(.A1(new_n532), .A2(new_n535), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n533), .B(KEYINPUT15), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT95), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(KEYINPUT95), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT96), .B(KEYINPUT17), .Z(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(G8gat), .Z(new_n549));
  OAI211_X1 g348(.A(new_n537), .B(KEYINPUT17), .C1(new_n538), .C2(new_n539), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n540), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(KEYINPUT18), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n553), .B(new_n554), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n557), .B(KEYINPUT13), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n551), .A2(new_n557), .A3(new_n555), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT93), .B(KEYINPUT12), .Z(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n574), .A3(new_n561), .A4(new_n564), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n202), .B1(new_n529), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n435), .A2(new_n473), .A3(new_n517), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT35), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n354), .A2(new_n434), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n521), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n525), .A2(new_n527), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT97), .A3(new_n576), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  AND2_X1   g387(.A1(G71gat), .A2(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(KEYINPUT9), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n591), .B(new_n593), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n268), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n554), .B1(KEYINPUT21), .B2(new_n595), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G232gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n407), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n609), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT7), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT99), .Z(new_n619));
  NOR2_X1   g418(.A1(new_n617), .A2(KEYINPUT7), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT100), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n616), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n623), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(KEYINPUT101), .A3(new_n623), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n544), .A2(new_n550), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n553), .A2(new_n631), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n612), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n633), .B2(new_n635), .ZN(new_n642));
  AOI211_X1 g441(.A(new_n634), .B(new_n637), .C1(new_n630), .C2(new_n632), .ZN(new_n643));
  INV_X1    g442(.A(new_n612), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n606), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648));
  INV_X1    g447(.A(G230gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n407), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n624), .A2(new_n595), .A3(new_n626), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n629), .A2(KEYINPUT103), .A3(new_n594), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n627), .A2(new_n594), .A3(new_n628), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n595), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n650), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n656), .A2(new_n649), .A3(new_n407), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n648), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n647), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n586), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n354), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n470), .ZN(new_n676));
  OAI21_X1  g475(.A(G8gat), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n470), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n680), .A2(KEYINPUT105), .A3(new_n678), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT105), .B1(new_n680), .B2(new_n678), .ZN(new_n682));
  OAI221_X1 g481(.A(new_n677), .B1(new_n678), .B2(new_n680), .C1(new_n681), .C2(new_n682), .ZN(G1325gat));
  NOR3_X1   g482(.A1(new_n672), .A2(G15gat), .A3(new_n526), .ZN(new_n684));
  INV_X1    g483(.A(new_n517), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n673), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(G15gat), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n263), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  INV_X1    g491(.A(new_n669), .ZN(new_n693));
  INV_X1    g492(.A(new_n606), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n646), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n578), .B2(new_n585), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n534), .A3(new_n354), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n698), .B(new_n699), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n695), .A2(new_n576), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n518), .B2(new_n528), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n579), .B(KEYINPUT108), .C1(new_n582), .C2(new_n583), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n638), .A2(new_n612), .A3(new_n640), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n644), .B1(new_n642), .B2(new_n643), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT109), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n705), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT44), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(new_n704), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n703), .A2(KEYINPUT110), .A3(new_n704), .A4(new_n710), .ZN(new_n715));
  INV_X1    g514(.A(new_n646), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT44), .B1(new_n529), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n519), .B(new_n701), .C1(new_n714), .C2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n700), .B1(new_n534), .B2(new_n720), .ZN(G1328gat));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n531), .A3(new_n470), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT46), .Z(new_n723));
  AOI211_X1 g522(.A(new_n676), .B(new_n701), .C1(new_n714), .C2(new_n719), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n531), .B2(new_n724), .ZN(G1329gat));
  NOR2_X1   g524(.A1(KEYINPUT112), .A2(KEYINPUT47), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n526), .A2(G43gat), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n697), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n697), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n701), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n685), .B(new_n735), .C1(new_n713), .C2(new_n718), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n726), .B(new_n729), .C1(new_n734), .C2(new_n737), .ZN(new_n738));
  AND4_X1   g537(.A1(new_n727), .A2(new_n734), .A3(new_n737), .A4(new_n728), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n263), .A2(G50gat), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n697), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n743), .B2(KEYINPUT114), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n264), .B(new_n735), .C1(new_n713), .C2(new_n718), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n744), .B(new_n746), .C1(KEYINPUT114), .C2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  INV_X1    g547(.A(new_n743), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n748), .B1(new_n750), .B2(new_n741), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n743), .B1(new_n745), .B2(G50gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(KEYINPUT113), .A3(KEYINPUT48), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n747), .B1(new_n751), .B2(new_n753), .ZN(G1331gat));
  AND2_X1   g553(.A1(new_n703), .A2(new_n704), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n669), .A2(new_n576), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n756), .A2(new_n647), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n354), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n758), .A2(new_n676), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n758), .B2(new_n517), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n526), .A2(G71gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n759), .A2(new_n264), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  OAI211_X1 g571(.A(new_n606), .B(new_n756), .C1(new_n713), .C2(new_n718), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n519), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n694), .A2(new_n576), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n584), .A2(new_n646), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n776), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n669), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n614), .A3(new_n354), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n774), .A2(new_n783), .ZN(G1336gat));
  NOR2_X1   g583(.A1(new_n676), .A2(G92gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n782), .A2(new_n785), .B1(new_n786), .B2(KEYINPUT52), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g587(.A(G92gat), .B1(new_n773), .B2(new_n676), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(G1337gat));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n773), .A2(new_n793), .A3(new_n517), .ZN(new_n794));
  INV_X1    g593(.A(new_n526), .ZN(new_n795));
  AOI21_X1  g594(.A(G99gat), .B1(new_n782), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(G1338gat));
  OAI21_X1  g596(.A(G106gat), .B1(new_n773), .B2(new_n263), .ZN(new_n798));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n799), .A3(new_n264), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n641), .B2(new_n645), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n705), .A2(new_n706), .A3(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g608(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n810));
  AOI21_X1  g609(.A(new_n665), .B1(new_n660), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g610(.A(KEYINPUT10), .B(new_n651), .C1(new_n652), .C2(new_n655), .ZN(new_n812));
  INV_X1    g611(.A(new_n659), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n812), .A2(new_n813), .B1(new_n649), .B2(new_n407), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n658), .A2(new_n650), .A3(new_n659), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT54), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n816), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n576), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n556), .A2(new_n557), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n559), .A2(new_n560), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n570), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n575), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n667), .A3(new_n668), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n809), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n819), .A2(new_n826), .A3(new_n820), .A4(new_n821), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n709), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n606), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n671), .A2(new_n577), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n521), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n519), .A2(new_n470), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n577), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n519), .B1(new_n831), .B2(new_n832), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n527), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n576), .A2(new_n271), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n842), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n836), .A2(new_n272), .A3(new_n669), .ZN(new_n844));
  AOI21_X1  g643(.A(G120gat), .B1(new_n839), .B2(new_n693), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n836), .B2(new_n606), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n839), .A2(new_n268), .A3(new_n694), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  NAND3_X1  g648(.A1(new_n839), .A2(new_n266), .A3(new_n646), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n836), .B2(new_n716), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  AND2_X1   g653(.A1(new_n835), .A2(new_n517), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n646), .B1(new_n822), .B2(new_n827), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n830), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n832), .B1(new_n857), .B2(new_n694), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n264), .A2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n833), .B2(new_n264), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(KEYINPUT119), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(KEYINPUT57), .C1(new_n833), .C2(new_n264), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n576), .B(new_n855), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G141gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n517), .A2(new_n264), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n470), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n838), .A2(new_n868), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n869), .A2(G141gat), .A3(new_n577), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n866), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(new_n869), .ZN(new_n876));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n693), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n855), .B1(new_n862), .B2(new_n864), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n669), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(KEYINPUT59), .A3(new_n877), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n833), .A2(new_n859), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n829), .A2(new_n716), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n606), .B1(new_n856), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n832), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n885), .B2(new_n264), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n855), .A2(new_n693), .ZN(new_n888));
  OAI21_X1  g687(.A(G148gat), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(KEYINPUT59), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n878), .B1(new_n881), .B2(new_n890), .ZN(G1345gat));
  NOR3_X1   g690(.A1(new_n879), .A2(new_n204), .A3(new_n606), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n869), .A2(new_n606), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT120), .ZN(new_n894));
  AOI21_X1  g693(.A(G155gat), .B1(new_n893), .B2(KEYINPUT120), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1346gat));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n205), .A3(new_n709), .ZN(new_n897));
  AOI21_X1  g696(.A(G162gat), .B1(new_n876), .B2(new_n646), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n354), .A2(new_n676), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT121), .Z(new_n901));
  NAND3_X1  g700(.A1(new_n833), .A2(new_n521), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n833), .A2(KEYINPUT122), .A3(new_n521), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n577), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n834), .A2(new_n900), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n365), .A3(new_n576), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n906), .B2(new_n669), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n366), .A3(new_n693), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n694), .A3(new_n905), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n606), .A2(new_n387), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n914), .A2(G183gat), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT60), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n921), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n908), .A2(new_n361), .A3(new_n809), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n646), .A3(new_n905), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(G190gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n924), .B2(G190gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  XOR2_X1   g727(.A(KEYINPUT124), .B(G197gat), .Z(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n517), .B(new_n901), .C1(new_n882), .C2(new_n886), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n577), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n867), .A2(new_n354), .A3(new_n676), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n833), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n576), .A3(new_n929), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n936), .ZN(G1352gat));
  AND2_X1   g736(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n938));
  NOR2_X1   g737(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g739(.A(KEYINPUT125), .B(G204gat), .Z(new_n941));
  NOR3_X1   g740(.A1(new_n934), .A2(new_n669), .A3(new_n941), .ZN(new_n942));
  MUX2_X1   g741(.A(new_n940), .B(new_n938), .S(new_n942), .Z(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n931), .B2(new_n669), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1353gat));
  NAND3_X1  g748(.A1(new_n935), .A2(new_n218), .A3(new_n694), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n931), .A2(new_n606), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n931), .B2(new_n716), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n219), .A3(new_n809), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1355gat));
endmodule


