//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT68), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n472), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n469), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n482), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(KEYINPUT69), .A2(G138), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n462), .B(new_n489), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n469), .A2(G126), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n491), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n500), .A2(KEYINPUT72), .A3(KEYINPUT5), .A4(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(new_n509), .A3(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n509), .B2(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n506), .A2(KEYINPUT70), .A3(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n505), .A2(new_n516), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n511), .A2(new_n515), .A3(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n503), .A2(new_n504), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n499), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n507), .A2(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n520), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n524), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n521), .A2(new_n506), .ZN(new_n530));
  NOR3_X1   g105(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT74), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n525), .A2(G51), .A3(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n525), .A2(G89), .A3(new_n520), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n520), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n534), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n534), .A2(new_n535), .A3(new_n540), .A4(KEYINPUT75), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(new_n518), .A2(G52), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n525), .A2(G90), .A3(new_n520), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n546), .B(new_n547), .C1(new_n506), .C2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND4_X1  g125(.A1(new_n520), .A2(G81), .A3(new_n515), .A4(new_n511), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n511), .A2(new_n515), .A3(G43), .A4(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n503), .B2(new_n504), .ZN(new_n559));
  INV_X1    g134(.A(G68), .ZN(new_n560));
  INV_X1    g135(.A(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT76), .B1(new_n563), .B2(new_n506), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n565), .B(G651), .C1(new_n559), .C2(new_n562), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n557), .A2(KEYINPUT78), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT78), .B1(new_n557), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(new_n571));
  XOR2_X1   g146(.A(new_n571), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n577));
  AND4_X1   g152(.A1(G53), .A2(new_n511), .A3(new_n515), .A4(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n511), .A2(new_n515), .A3(G53), .A4(G543), .ZN(new_n581));
  NOR3_X1   g156(.A1(new_n581), .A2(KEYINPUT81), .A3(KEYINPUT9), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n581), .A2(KEYINPUT80), .A3(KEYINPUT9), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT80), .B1(new_n581), .B2(KEYINPUT9), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n580), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n520), .A2(G65), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT82), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n517), .A2(G91), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n585), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G168), .ZN(G286));
  INV_X1    g168(.A(KEYINPUT83), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n523), .B2(new_n531), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT74), .B1(new_n529), .B2(new_n530), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n519), .A2(new_n522), .A3(new_n499), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT83), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n598), .ZN(G303));
  NAND3_X1  g174(.A1(new_n525), .A2(G49), .A3(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT84), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n520), .A2(G74), .ZN(new_n602));
  AOI22_X1  g177(.A1(G87), .A2(new_n517), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(G288));
  AOI22_X1  g179(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n506), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n517), .A2(G86), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n518), .A2(G48), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(G305));
  AOI22_X1  g184(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n610), .A2(new_n506), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n518), .A2(G47), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n517), .A2(G85), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(G290));
  NAND2_X1  g189(.A1(G301), .A2(G868), .ZN(new_n615));
  AND4_X1   g190(.A1(G54), .A2(new_n511), .A3(new_n515), .A4(G543), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n505), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n619), .B2(G651), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n520), .A2(G92), .A3(new_n515), .A4(new_n511), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g198(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .A4(new_n520), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n615), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n615), .B1(new_n627), .B2(G868), .ZN(G321));
  MUX2_X1   g204(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g205(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n627), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n570), .B2(G868), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n481), .A2(G135), .ZN(new_n638));
  INV_X1    g213(.A(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n462), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI221_X1 g216(.A(new_n638), .B1(new_n486), .B2(new_n639), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT85), .B(G2100), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT86), .ZN(G401));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2100), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n681), .B2(new_n686), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(KEYINPUT87), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n681), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n688), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  XOR2_X1   g276(.A(KEYINPUT89), .B(G29), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(G27), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G164), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G2078), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT31), .B(G11), .Z(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G28), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(KEYINPUT96), .B1(new_n710), .B2(G28), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT26), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(KEYINPUT26), .ZN(new_n718));
  INV_X1    g293(.A(G129), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n717), .B(new_n718), .C1(new_n486), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G141), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n709), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n709), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n715), .B1(new_n642), .B2(new_n702), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n709), .A2(G33), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n469), .A2(G127), .ZN(new_n732));
  AND2_X1   g307(.A1(G115), .A2(G2104), .ZN(new_n733));
  OAI21_X1  g308(.A(G2105), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT25), .ZN(new_n735));
  NAND2_X1  g310(.A1(G103), .A2(G2104), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n481), .A2(G139), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n731), .B1(new_n740), .B2(G29), .ZN(new_n741));
  INV_X1    g316(.A(G2072), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n729), .A2(new_n730), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G34), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n703), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n479), .B2(new_n709), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2084), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n752), .ZN(new_n754));
  INV_X1    g329(.A(G1961), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  AND4_X1   g331(.A1(new_n707), .A2(new_n745), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n752), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n752), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G1966), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT97), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(G1966), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n702), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT93), .Z(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n481), .A2(G140), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n770));
  INV_X1    g345(.A(G128), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n770), .C1(new_n771), .C2(new_n486), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n766), .A2(KEYINPUT28), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n767), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n703), .A2(G35), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G162), .B2(new_n703), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n779), .B2(G2090), .ZN(new_n780));
  NOR2_X1   g355(.A1(G4), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n627), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT92), .B(G1348), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n782), .A2(new_n784), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n780), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n779), .A2(G2090), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n752), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n787), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n763), .A2(KEYINPUT98), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n752), .A2(G19), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n570), .B2(new_n752), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1341), .Z(new_n799));
  NAND4_X1  g374(.A1(new_n764), .A2(new_n795), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G290), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G16), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G1986), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n481), .A2(G131), .ZN(new_n805));
  INV_X1    g380(.A(G119), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n462), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n805), .B1(new_n486), .B2(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G25), .B(new_n809), .S(new_n703), .Z(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n803), .A2(G1986), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G6), .A2(G16), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT32), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1981), .Z(new_n820));
  MUX2_X1   g395(.A(G23), .B(G288), .S(G16), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT33), .B(G1976), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n752), .A2(G22), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT90), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n752), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n823), .B1(G1971), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n820), .B(new_n827), .C1(G1971), .C2(new_n826), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n804), .B(new_n815), .C1(new_n828), .C2(KEYINPUT34), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(KEYINPUT34), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n800), .B1(new_n832), .B2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  INV_X1    g410(.A(new_n800), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(G150));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n838), .A2(new_n526), .B1(new_n527), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n506), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n568), .B2(new_n569), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n505), .A2(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n565), .B1(new_n846), .B2(G651), .ZN(new_n847));
  INV_X1    g422(.A(new_n566), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n555), .B1(new_n551), .B2(new_n552), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n847), .A2(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT38), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n626), .A2(new_n632), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n844), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n462), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n486), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G142), .B2(new_n481), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n645), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n725), .B(new_n740), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n772), .B(new_n497), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n809), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n479), .B(G162), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n642), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n874), .B(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(KEYINPUT100), .B(G37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g455(.A(new_n634), .B(KEYINPUT101), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n854), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  INV_X1    g458(.A(new_n584), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n581), .A2(KEYINPUT80), .A3(KEYINPUT9), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n518), .A2(new_n577), .A3(new_n579), .A4(G53), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT81), .B1(new_n581), .B2(KEYINPUT9), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n884), .A2(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n589), .A2(new_n590), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n626), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(new_n585), .A2(new_n591), .B1(new_n625), .B2(new_n620), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n627), .A2(new_n585), .A3(new_n591), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n626), .B1(new_n888), .B2(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n882), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n890), .A2(new_n891), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n532), .A2(G290), .ZN(new_n901));
  AOI21_X1  g476(.A(G290), .B1(new_n596), .B2(new_n597), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G288), .A2(new_n817), .ZN(new_n904));
  NAND3_X1  g479(.A1(G305), .A2(new_n601), .A3(new_n603), .ZN(new_n905));
  AND4_X1   g480(.A1(new_n901), .A2(new_n903), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n901), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n900), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n900), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g488(.A(new_n912), .B1(G868), .B2(new_n843), .ZN(G331));
  XOR2_X1   g489(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n915));
  AND2_X1   g490(.A1(new_n892), .A2(new_n895), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT78), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n851), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n557), .A2(KEYINPUT78), .A3(new_n567), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n843), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G301), .B1(new_n543), .B2(new_n544), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n543), .A2(G301), .A3(new_n544), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n920), .A2(new_n924), .A3(new_n852), .ZN(new_n925));
  INV_X1    g500(.A(new_n923), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(new_n921), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n845), .B2(new_n853), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n916), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n906), .A2(new_n907), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n920), .B2(new_n852), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n845), .A2(new_n853), .A3(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n898), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n878), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n933), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n938), .B2(new_n908), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n938), .B2(new_n908), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n941), .B2(new_n934), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(KEYINPUT103), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n944), .B(new_n935), .C1(new_n941), .C2(new_n934), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n915), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n936), .B2(new_n941), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n931), .A2(new_n898), .A3(new_n932), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n896), .B1(new_n932), .B2(new_n931), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n908), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n934), .A4(new_n878), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n939), .B2(new_n934), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n948), .B(KEYINPUT105), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(new_n878), .A3(new_n934), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT104), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT105), .B1(new_n960), .B2(new_n948), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n946), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n946), .B(KEYINPUT106), .C1(new_n957), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G397));
  AND3_X1   g541(.A1(new_n468), .A2(new_n478), .A3(G40), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n497), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n772), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT108), .ZN(new_n974));
  INV_X1    g549(.A(new_n725), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1996), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(KEYINPUT46), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n970), .B2(G1996), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n772), .A2(G2067), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n974), .A2(new_n971), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n985), .B(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n725), .B(new_n977), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n971), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(KEYINPUT110), .A3(new_n989), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n809), .A2(new_n812), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n983), .B1(new_n995), .B2(new_n970), .ZN(new_n996));
  NOR2_X1   g571(.A1(G290), .A2(G1986), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(new_n970), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n809), .B(new_n811), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT111), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n971), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n993), .A2(KEYINPUT127), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n991), .A2(new_n992), .A3(new_n1003), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1000), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n996), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n1010));
  AND3_X1   g585(.A1(G290), .A2(new_n1010), .A3(G1986), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(G290), .B2(G1986), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n970), .B(new_n1011), .C1(new_n998), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1005), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n468), .A2(new_n478), .A3(G40), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n969), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n497), .A2(new_n968), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1971), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n967), .A2(new_n1025), .A3(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n497), .B2(new_n968), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1015), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1022), .B1(new_n1031), .B2(G2090), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(G8), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n596), .A2(new_n597), .A3(KEYINPUT83), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT83), .B1(new_n596), .B2(new_n597), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT55), .B(G8), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  NAND4_X1  g616(.A1(G303), .A2(new_n1041), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1033), .A2(new_n1037), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1042), .A3(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n497), .A2(new_n968), .A3(new_n1023), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n967), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2090), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1049), .B1(new_n1022), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1020), .A2(KEYINPUT112), .A3(new_n1021), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(new_n1045), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1056), .B(new_n1058), .C1(new_n1057), .C2(G288), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n967), .A2(new_n1018), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G288), .A2(new_n1057), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT115), .B(G1981), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n817), .A2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(G305), .B2(G1981), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1064), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(new_n1020), .B2(G2078), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1048), .A2(new_n755), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1017), .A2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(new_n1015), .A3(new_n969), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1079), .A2(KEYINPUT53), .A3(new_n706), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(G301), .ZN(new_n1083));
  AND4_X1   g658(.A1(new_n1043), .A2(new_n1054), .A3(new_n1073), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  INV_X1    g660(.A(G2084), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n967), .A2(new_n1046), .A3(new_n1086), .A4(new_n1047), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1079), .B2(G1966), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(KEYINPUT123), .B2(G286), .ZN(new_n1089));
  OAI211_X1 g664(.A(G168), .B(new_n1087), .C1(new_n1079), .C2(G1966), .ZN(new_n1090));
  NOR2_X1   g665(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT123), .B1(new_n1090), .B2(G8), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1095), .B2(KEYINPUT122), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1085), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1085), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1084), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(G1976), .B(G288), .C1(new_n1072), .C2(new_n1071), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1066), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1056), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1073), .A2(new_n1044), .A3(new_n1053), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n1020), .B2(G1996), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1079), .A2(new_n1108), .A3(new_n977), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1060), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n570), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1115), .A3(new_n570), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT61), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT56), .B(G2072), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1031), .A2(new_n793), .B1(new_n1079), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n585), .B2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(G299), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1048), .A2(new_n783), .B1(new_n1055), .B2(new_n972), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(new_n626), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n626), .A2(KEYINPUT60), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1129), .A2(KEYINPUT60), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT61), .A3(new_n1124), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1117), .A2(new_n1127), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1128), .A2(new_n626), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1126), .B1(new_n1124), .B2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1054), .A2(new_n1073), .A3(new_n1043), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1082), .A2(KEYINPUT124), .A3(G301), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1081), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(KEYINPUT54), .A3(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1138), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1100), .B(new_n1106), .C1(new_n1137), .C2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT118), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1088), .A2(new_n1150), .A3(G8), .A4(G168), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1054), .A2(new_n1043), .A3(new_n1073), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1155), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1054), .A3(new_n1073), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1154), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1157), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT125), .B(new_n1014), .C1(new_n1147), .C2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1099), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(new_n1097), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1105), .B1(new_n1169), .B2(new_n1084), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1171), .A2(new_n1138), .A3(new_n1143), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1167), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n1174), .B2(new_n1014), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1009), .B1(new_n1165), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g751(.A1(new_n943), .A2(new_n945), .ZN(new_n1178));
  NOR4_X1   g752(.A1(G229), .A2(new_n460), .A3(new_n665), .A4(G227), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n1178), .A2(new_n879), .A3(new_n1179), .ZN(G225));
  INV_X1    g754(.A(G225), .ZN(G308));
endmodule


