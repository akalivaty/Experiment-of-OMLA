//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n206));
  OR2_X1    g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT77), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G155gat), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n209), .A2(new_n213), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(KEYINPUT78), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT78), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G155gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n215), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n219), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT78), .B(G155gat), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT79), .B(KEYINPUT2), .C1(new_n226), .C2(new_n215), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(new_n205), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(new_n207), .A3(new_n208), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n218), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G211gat), .B(G218gat), .Z(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  INV_X1    g036(.A(G218gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT29), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n233), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n232), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT75), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n242), .B1(new_n246), .B2(new_n234), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(KEYINPUT75), .A3(new_n233), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n230), .B1(new_n225), .B2(new_n227), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n251), .A2(KEYINPUT3), .A3(new_n218), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n245), .B1(new_n253), .B2(KEYINPUT85), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n231), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n217), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT29), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n204), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(new_n252), .B2(KEYINPUT29), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n257), .A2(KEYINPUT86), .A3(new_n258), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n250), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n249), .B(new_n258), .C1(new_n218), .C2(new_n251), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(new_n251), .B2(new_n218), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n267), .A2(new_n268), .A3(new_n204), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n266), .A2(KEYINPUT87), .A3(new_n269), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n262), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT88), .ZN(new_n275));
  INV_X1    g074(.A(G22gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n245), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n259), .B2(new_n260), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n253), .A2(KEYINPUT85), .ZN(new_n279));
  OAI22_X1  g078(.A1(new_n278), .A2(new_n279), .B1(new_n202), .B2(new_n203), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n266), .A2(KEYINPUT87), .A3(new_n269), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT87), .B1(new_n266), .B2(new_n269), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT31), .B(G50gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT84), .ZN(new_n287));
  XOR2_X1   g086(.A(G78gat), .B(G106gat), .Z(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  AOI21_X1  g088(.A(new_n276), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  AOI211_X1 g090(.A(G22gat), .B(new_n291), .C1(new_n283), .C2(new_n284), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n275), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n274), .B2(KEYINPUT88), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G22gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n275), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n276), .A3(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G113gat), .ZN(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  INV_X1    g107(.A(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(KEYINPUT1), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT69), .B(G127gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n309), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n307), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n257), .A2(new_n268), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n217), .B(new_n307), .C1(new_n314), .C2(new_n312), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n255), .A3(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT80), .B1(new_n251), .B2(new_n317), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n255), .A2(new_n217), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n306), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G127gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n328));
  OAI21_X1  g127(.A(G134gat), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n329), .A3(new_n310), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n324), .B1(new_n330), .B2(new_n307), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n307), .B(new_n324), .C1(new_n312), .C2(new_n314), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n323), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n316), .B(new_n322), .C1(new_n334), .C2(KEYINPUT4), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT39), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  AND2_X1   g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n319), .B1(new_n318), .B2(new_n255), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n251), .A2(new_n317), .A3(KEYINPUT80), .ZN(new_n346));
  INV_X1    g145(.A(new_n315), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n345), .A2(new_n346), .B1(new_n232), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT39), .B1(new_n348), .B2(new_n338), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT89), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT89), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(KEYINPUT39), .C1(new_n348), .C2(new_n338), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n338), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n344), .A2(KEYINPUT40), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT40), .B1(new_n344), .B2(new_n354), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n334), .A2(KEYINPUT4), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n316), .A2(new_n337), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .A4(new_n322), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n320), .A2(new_n321), .B1(new_n323), .B2(new_n315), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(new_n337), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n348), .A2(KEYINPUT82), .A3(new_n338), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(KEYINPUT5), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT4), .B1(new_n320), .B2(new_n321), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n315), .A2(KEYINPUT70), .ZN(new_n369));
  AND4_X1   g168(.A1(KEYINPUT4), .A2(new_n232), .A3(new_n369), .A4(new_n332), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT81), .B1(new_n371), .B2(new_n360), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n316), .A2(new_n337), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  NOR4_X1   g173(.A1(new_n373), .A2(new_n368), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n367), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n348), .A2(new_n338), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n359), .B1(new_n377), .B2(new_n362), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n366), .B1(new_n378), .B2(new_n365), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n361), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n343), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT24), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G183gat), .ZN(new_n386));
  INV_X1    g185(.A(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G169gat), .ZN(new_n392));
  INV_X1    g191(.A(G176gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT64), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G176gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G169gat), .A2(G176gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT23), .ZN(new_n399));
  INV_X1    g198(.A(G169gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n393), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n390), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT65), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT65), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT66), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n383), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n384), .A2(KEYINPUT67), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT24), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n388), .A2(new_n389), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n393), .A3(KEYINPUT23), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n417), .A2(KEYINPUT25), .A3(new_n402), .A4(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n406), .A2(new_n408), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT28), .ZN(new_n421));
  XNOR2_X1  g220(.A(KEYINPUT27), .B(G183gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(KEYINPUT68), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT68), .B1(new_n386), .B2(KEYINPUT27), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n387), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(KEYINPUT28), .A3(new_n387), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT26), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n401), .A2(new_n429), .A3(new_n398), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n383), .B1(new_n401), .B2(new_n429), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT29), .B1(new_n420), .B2(new_n433), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n250), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n436), .B(new_n249), .C1(new_n435), .C2(new_n437), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G64gat), .B(G92gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT30), .A4(new_n444), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(new_n440), .A3(new_n444), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n357), .A2(new_n382), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n299), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n343), .A2(KEYINPUT6), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n381), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n380), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n371), .A2(new_n360), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n374), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n371), .A2(new_n360), .A3(KEYINPUT81), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n364), .A2(KEYINPUT5), .ZN(new_n464));
  INV_X1    g263(.A(new_n365), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT83), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n466), .A3(new_n367), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n467), .A2(new_n457), .A3(new_n361), .A4(new_n381), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT90), .B(KEYINPUT37), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n439), .A2(new_n440), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT91), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n439), .A2(new_n440), .A3(new_n472), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT38), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n444), .B1(new_n441), .B2(KEYINPUT37), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n459), .A2(new_n468), .A3(new_n450), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT92), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT38), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n478), .B2(KEYINPUT92), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n455), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT74), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n333), .A2(new_n331), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n391), .B1(G169gat), .B2(G176gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(G169gat), .A2(G176gat), .ZN(new_n491));
  OAI211_X1 g290(.A(KEYINPUT25), .B(new_n418), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n416), .B2(new_n415), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n430), .B(new_n431), .C1(new_n426), .C2(new_n427), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT71), .B(new_n487), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n333), .B2(new_n331), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n369), .A2(KEYINPUT71), .A3(new_n332), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n498), .A2(new_n433), .A3(new_n499), .A4(new_n420), .ZN(new_n500));
  NAND2_X1  g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT32), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n506), .A3(KEYINPUT32), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n503), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n505), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n503), .B(KEYINPUT32), .C1(new_n511), .C2(new_n510), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n502), .B1(new_n496), .B2(new_n500), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n513), .A2(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n496), .A2(new_n500), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n501), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT34), .B1(new_n524), .B2(KEYINPUT73), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n518), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n513), .A3(new_n514), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n486), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n514), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n486), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n485), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n527), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n533), .A2(new_n485), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n459), .A2(new_n468), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n448), .A2(KEYINPUT76), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n446), .A2(new_n538), .A3(new_n447), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n536), .A2(new_n452), .A3(new_n537), .A4(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n532), .A2(new_n535), .B1(new_n540), .B2(new_n299), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n484), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n536), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n543), .A2(new_n531), .A3(new_n528), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n299), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n526), .A2(new_n514), .A3(new_n513), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(new_n521), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n293), .A2(new_n298), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT35), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G197gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT11), .B(G169gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT12), .Z(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G15gat), .B(G22gat), .Z(new_n562));
  INV_X1    g361(.A(G1gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n565), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G8gat), .ZN(new_n569));
  INV_X1    g368(.A(G8gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n564), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G43gat), .B(G50gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n575));
  INV_X1    g374(.A(G29gat), .ZN(new_n576));
  INV_X1    g375(.A(G36gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n574), .A2(KEYINPUT15), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n581));
  INV_X1    g380(.A(G43gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(G50gat), .ZN(new_n583));
  INV_X1    g382(.A(G50gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(G43gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G29gat), .A2(G36gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(G29gat), .A3(G36gat), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n588), .A2(new_n590), .A3(KEYINPUT96), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT96), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n580), .B(new_n586), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(KEYINPUT94), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n578), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n588), .A2(new_n590), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n584), .A2(G43gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n582), .A2(G50gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT15), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n593), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n593), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n573), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n569), .A2(new_n571), .B1(new_n593), .B2(new_n604), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT18), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n608), .A2(new_n609), .A3(new_n611), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n609), .B(KEYINPUT13), .Z(new_n616));
  NOR2_X1   g415(.A1(new_n591), .A2(new_n592), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n578), .A2(new_n579), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n586), .A2(new_n602), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n588), .A2(new_n590), .ZN(new_n620));
  NOR2_X1   g419(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n579), .A2(new_n594), .B1(new_n621), .B2(new_n577), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n622), .B2(new_n596), .ZN(new_n623));
  OAI22_X1  g422(.A1(new_n617), .A2(new_n619), .B1(new_n623), .B2(new_n602), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n572), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n616), .B1(new_n625), .B2(new_n610), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n615), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(KEYINPUT17), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n593), .A2(new_n604), .A3(new_n605), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n610), .B1(new_n630), .B2(new_n573), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n614), .B1(new_n631), .B2(new_n609), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n555), .B(new_n561), .C1(new_n627), .C2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n613), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n636), .A2(new_n626), .A3(new_n615), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n561), .B1(new_n637), .B2(new_n555), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n554), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(G57gat), .A2(G64gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(G57gat), .A2(G64gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(G71gat), .A2(G78gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(G71gat), .A2(G78gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT99), .B1(new_n645), .B2(KEYINPUT9), .ZN(new_n649));
  NAND2_X1  g448(.A1(G71gat), .A2(G78gat), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT9), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G71gat), .B(G78gat), .ZN(new_n657));
  AND2_X1   g456(.A1(G57gat), .A2(G64gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(G57gat), .A2(G64gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n652), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT98), .B1(new_n658), .B2(new_n659), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n651), .B1(new_n650), .B2(new_n652), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n660), .A2(new_n657), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT100), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n656), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n572), .B1(new_n670), .B2(KEYINPUT21), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n214), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n673), .B(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(G231gat), .B(G233gat), .C1(new_n670), .C2(KEYINPUT21), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n655), .B1(new_n648), .B2(new_n654), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n642), .A2(new_n661), .A3(new_n643), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n663), .A3(KEYINPUT9), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n647), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT21), .ZN(new_n684));
  NAND2_X1  g483(.A1(G231gat), .A2(G233gat), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n656), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n308), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(G127gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G183gat), .B(G211gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n691), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n677), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n694), .A3(new_n676), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(G99gat), .ZN(new_n701));
  INV_X1    g500(.A(G106gat), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT8), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(G85gat), .A2(G92gat), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT7), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G85gat), .ZN(new_n708));
  INV_X1    g507(.A(G92gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(G99gat), .B(G106gat), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n704), .A2(new_n705), .ZN(new_n716));
  NAND3_X1  g515(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(KEYINPUT7), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n712), .A2(new_n714), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  OAI211_X1 g519(.A(KEYINPUT104), .B(new_n713), .C1(new_n720), .C2(new_n711), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n628), .B2(new_n629), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n624), .ZN(new_n724));
  AND2_X1   g523(.A1(G232gat), .A2(G233gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT41), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(G190gat), .B(G218gat), .Z(new_n728));
  OR3_X1    g527(.A1(new_n723), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n723), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n725), .A2(KEYINPUT41), .ZN(new_n732));
  XNOR2_X1  g531(.A(G134gat), .B(G162gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n734), .A3(new_n730), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(G120gat), .B(G148gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(G176gat), .B(G204gat), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n739), .B(new_n740), .Z(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(G230gat), .A2(G233gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n670), .A2(new_n722), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n683), .A2(new_n656), .A3(new_n721), .A4(new_n719), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT10), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n670), .A2(KEYINPUT10), .A3(new_n722), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n745), .A2(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n744), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n742), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n748), .A2(new_n749), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n743), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT105), .B(new_n744), .C1(new_n748), .C2(new_n749), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n752), .A2(new_n741), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT106), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n757), .A2(new_n758), .A3(new_n763), .A4(new_n760), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n754), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n700), .A2(new_n738), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n641), .A2(new_n543), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G1gat), .ZN(G1324gat));
  NOR3_X1   g569(.A1(new_n554), .A2(new_n640), .A3(new_n767), .ZN(new_n771));
  XNOR2_X1  g570(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G8gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n453), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n641), .A2(new_n768), .ZN(new_n775));
  INV_X1    g574(.A(new_n453), .ZN(new_n776));
  OAI21_X1  g575(.A(G8gat), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n774), .ZN(new_n778));
  MUX2_X1   g577(.A(new_n774), .B(new_n778), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g578(.A1(new_n528), .A2(new_n531), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n775), .A2(G15gat), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n532), .A2(new_n535), .ZN(new_n783));
  OAI21_X1  g582(.A(G15gat), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1326gat));
  NAND2_X1  g584(.A1(new_n771), .A2(new_n299), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT43), .B(G22gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1327gat));
  NOR3_X1   g587(.A1(new_n700), .A2(new_n738), .A3(new_n765), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n536), .A2(G29gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n553), .A2(new_n639), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(KEYINPUT108), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(KEYINPUT108), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(KEYINPUT45), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n792), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n738), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n738), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n804), .B1(new_n542), .B2(new_n552), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n293), .A2(new_n298), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n537), .A2(new_n452), .A3(new_n539), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n468), .B2(new_n459), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT74), .B1(new_n548), .B2(new_n521), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT36), .B1(new_n809), .B2(new_n530), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n806), .A2(new_n808), .B1(new_n810), .B2(new_n534), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n478), .A2(KEYINPUT92), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n479), .A3(new_n482), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n455), .ZN(new_n814));
  INV_X1    g613(.A(new_n550), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n808), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n816), .A2(KEYINPUT35), .B1(new_n544), .B2(new_n546), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n797), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n805), .B1(new_n818), .B2(KEYINPUT44), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n634), .B2(new_n638), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n555), .B1(new_n627), .B2(new_n632), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n560), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(KEYINPUT109), .A3(new_n633), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n700), .A2(new_n765), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT111), .B1(new_n819), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n803), .B1(new_n553), .B2(new_n797), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n830), .B(new_n826), .C1(new_n831), .C2(new_n805), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n829), .A2(new_n833), .A3(new_n536), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n796), .B1(new_n834), .B2(new_n576), .ZN(G1328gat));
  AND2_X1   g634(.A1(new_n641), .A2(new_n789), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n837));
  AOI211_X1 g636(.A(G36gat), .B(new_n776), .C1(new_n837), .C2(KEYINPUT46), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n837), .B2(KEYINPUT46), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n837), .A2(KEYINPUT46), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n841), .A3(new_n838), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n829), .A2(new_n833), .A3(new_n776), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n840), .B(new_n842), .C1(new_n843), .C2(new_n577), .ZN(G1329gat));
  NAND3_X1  g643(.A1(new_n836), .A2(new_n582), .A3(new_n780), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n819), .A2(new_n783), .A3(new_n827), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n845), .B(KEYINPUT47), .C1(new_n582), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n641), .A2(new_n789), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(G43gat), .A3(new_n781), .ZN(new_n849));
  INV_X1    g648(.A(new_n783), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n850), .A3(new_n832), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(G43gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n852), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n584), .A3(new_n299), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n819), .A2(new_n806), .A3(new_n827), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n854), .B(KEYINPUT48), .C1(new_n584), .C2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n848), .A2(G50gat), .A3(new_n806), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n828), .A2(new_n299), .A3(new_n832), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G50gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n859), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g659(.A1(new_n700), .A2(new_n738), .A3(new_n765), .A4(new_n825), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n554), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n543), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT113), .B(G57gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1332gat));
  NOR3_X1   g664(.A1(new_n554), .A2(new_n776), .A3(new_n861), .ZN(new_n866));
  NOR2_X1   g665(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n867));
  AND2_X1   g666(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n866), .B2(new_n867), .ZN(G1333gat));
  AOI21_X1  g669(.A(KEYINPUT114), .B1(new_n862), .B2(new_n780), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n554), .A2(new_n872), .A3(new_n781), .A4(new_n861), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n871), .A2(G71gat), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n862), .A2(G71gat), .A3(new_n850), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n871), .A2(G71gat), .A3(new_n873), .ZN(new_n878));
  INV_X1    g677(.A(new_n876), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT50), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(G1334gat));
  NAND2_X1  g680(.A1(new_n862), .A2(new_n299), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(G78gat), .ZN(G1335gat));
  INV_X1    g682(.A(new_n825), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n700), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n553), .A2(new_n797), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n766), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n708), .A3(new_n543), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n885), .A2(new_n765), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n819), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G85gat), .B1(new_n894), .B2(new_n536), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(new_n895), .ZN(G1336gat));
  AOI21_X1  g695(.A(new_n709), .B1(new_n893), .B2(new_n453), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n776), .A2(G92gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT52), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  AOI211_X1 g702(.A(new_n766), .B(new_n903), .C1(new_n888), .C2(new_n889), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT52), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1337gat));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n701), .A3(new_n780), .ZN(new_n907));
  OAI21_X1  g706(.A(G99gat), .B1(new_n894), .B2(new_n783), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1338gat));
  AOI21_X1  g708(.A(new_n702), .B1(new_n893), .B2(new_n299), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n299), .A2(new_n702), .A3(new_n765), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT115), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n915), .B1(new_n888), .B2(new_n889), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n912), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT53), .B1(new_n910), .B2(new_n916), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1339gat));
  NAND2_X1  g719(.A1(new_n756), .A2(new_n743), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n750), .A2(new_n755), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n761), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n763), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n759), .A2(KEYINPUT106), .A3(new_n761), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT54), .B1(new_n756), .B2(new_n743), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n757), .A3(new_n758), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n742), .B1(new_n921), .B2(KEYINPUT54), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n931), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n922), .A2(new_n923), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n933), .B(KEYINPUT55), .C1(new_n934), .C2(new_n929), .ZN(new_n935));
  INV_X1    g734(.A(new_n637), .ZN(new_n936));
  OR3_X1    g735(.A1(new_n625), .A2(new_n610), .A3(new_n616), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n631), .B2(new_n609), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n936), .A2(new_n561), .B1(new_n938), .B2(new_n559), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n927), .A2(new_n932), .A3(new_n935), .A4(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n801), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n765), .A2(new_n939), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n825), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n801), .B2(new_n944), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n945), .A2(new_n700), .B1(new_n767), .B2(new_n884), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(new_n806), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n536), .A2(new_n453), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n780), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G113gat), .B1(new_n951), .B2(new_n640), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n946), .A2(new_n948), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(new_n815), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT116), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n884), .A2(new_n302), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1340gat));
  OAI21_X1  g756(.A(G120gat), .B1(new_n951), .B2(new_n766), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n765), .A2(new_n300), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n955), .B2(new_n959), .ZN(G1341gat));
  OAI211_X1 g759(.A(new_n950), .B(new_n700), .C1(new_n327), .C2(new_n328), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT117), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n954), .A2(new_n700), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n963), .B(new_n964), .C1(new_n313), .C2(new_n965), .ZN(G1342gat));
  NAND3_X1  g765(.A1(new_n954), .A2(new_n309), .A3(new_n797), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n967), .A2(KEYINPUT56), .ZN(new_n968));
  OAI21_X1  g767(.A(G134gat), .B1(new_n951), .B2(new_n738), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(KEYINPUT56), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G1343gat));
  AND2_X1   g770(.A1(new_n783), .A2(new_n948), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n946), .A2(new_n299), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n973), .A2(KEYINPUT57), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n767), .A2(new_n884), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n942), .B1(new_n943), .B2(new_n640), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n738), .ZN(new_n977));
  INV_X1    g776(.A(new_n941), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n700), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT57), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n806), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n972), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(G141gat), .B1(new_n984), .B2(new_n640), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n850), .A2(new_n806), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n953), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n987), .A2(G141gat), .A3(new_n640), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n988), .A2(KEYINPUT58), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n984), .A2(new_n825), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n988), .B1(new_n991), .B2(G141gat), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT58), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1344gat));
  INV_X1    g793(.A(new_n987), .ZN(new_n995));
  INV_X1    g794(.A(G148gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n995), .A2(new_n996), .A3(new_n765), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT59), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n944), .A2(new_n801), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n700), .B1(new_n999), .B2(new_n978), .ZN(new_n1000));
  OAI211_X1 g799(.A(KEYINPUT57), .B(new_n299), .C1(new_n1000), .C2(new_n975), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(KEYINPUT120), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT120), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n946), .A2(new_n1003), .A3(KEYINPUT57), .A4(new_n299), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n940), .A2(new_n738), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n700), .B1(new_n977), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n767), .A2(new_n639), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n299), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(new_n982), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1002), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n766), .B1(new_n972), .B2(KEYINPUT119), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1011), .B1(KEYINPUT119), .B2(new_n972), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n996), .B1(new_n1013), .B2(KEYINPUT121), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT121), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1015), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n998), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n765), .B(new_n972), .C1(new_n974), .C2(new_n983), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n996), .A2(KEYINPUT59), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n1018), .A2(KEYINPUT118), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(KEYINPUT118), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n997), .B1(new_n1017), .B2(new_n1022), .ZN(G1345gat));
  INV_X1    g822(.A(new_n226), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1024), .B1(new_n984), .B2(new_n980), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n995), .A2(new_n226), .A3(new_n700), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1346gat));
  OR3_X1    g826(.A1(new_n984), .A2(new_n215), .A3(new_n801), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n215), .B1(new_n987), .B2(new_n738), .ZN(new_n1029));
  AND2_X1   g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1347gat));
  NOR2_X1   g829(.A1(new_n543), .A2(new_n776), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n946), .A2(new_n815), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1032), .A2(new_n400), .A3(new_n884), .ZN(new_n1033));
  XNOR2_X1  g832(.A(new_n1033), .B(KEYINPUT122), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n544), .A2(new_n453), .ZN(new_n1035));
  XNOR2_X1  g834(.A(new_n1035), .B(KEYINPUT123), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1036), .A2(new_n947), .ZN(new_n1037));
  OAI21_X1  g836(.A(G169gat), .B1(new_n1037), .B2(new_n640), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1034), .A2(new_n1038), .ZN(G1348gat));
  AOI21_X1  g838(.A(G176gat), .B1(new_n1032), .B2(new_n765), .ZN(new_n1040));
  XOR2_X1   g839(.A(new_n1040), .B(KEYINPUT124), .Z(new_n1041));
  AOI211_X1 g840(.A(new_n766), .B(new_n1037), .C1(new_n394), .C2(new_n396), .ZN(new_n1042));
  NOR2_X1   g841(.A1(new_n1041), .A2(new_n1042), .ZN(G1349gat));
  NAND3_X1  g842(.A1(new_n1032), .A2(new_n422), .A3(new_n700), .ZN(new_n1044));
  XNOR2_X1  g843(.A(new_n1044), .B(KEYINPUT125), .ZN(new_n1045));
  OAI21_X1  g844(.A(G183gat), .B1(new_n1037), .B2(new_n980), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g846(.A(new_n1047), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g847(.A1(new_n1032), .A2(new_n387), .A3(new_n802), .ZN(new_n1049));
  OAI21_X1  g848(.A(G190gat), .B1(new_n1037), .B2(new_n738), .ZN(new_n1050));
  AND2_X1   g849(.A1(new_n1050), .A2(KEYINPUT61), .ZN(new_n1051));
  NOR2_X1   g850(.A1(new_n1050), .A2(KEYINPUT61), .ZN(new_n1052));
  OAI21_X1  g851(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(G1351gat));
  AND2_X1   g852(.A1(new_n783), .A2(new_n1031), .ZN(new_n1054));
  NAND2_X1  g853(.A1(new_n973), .A2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g854(.A1(new_n1055), .A2(G197gat), .A3(new_n825), .ZN(new_n1056));
  XOR2_X1   g855(.A(new_n1056), .B(KEYINPUT126), .Z(new_n1057));
  NAND3_X1  g856(.A1(new_n1002), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1058));
  NAND2_X1  g857(.A1(new_n1058), .A2(new_n1054), .ZN(new_n1059));
  OAI21_X1  g858(.A(G197gat), .B1(new_n1059), .B2(new_n640), .ZN(new_n1060));
  NAND2_X1  g859(.A1(new_n1057), .A2(new_n1060), .ZN(G1352gat));
  NOR3_X1   g860(.A1(new_n1055), .A2(G204gat), .A3(new_n766), .ZN(new_n1062));
  XNOR2_X1  g861(.A(new_n1062), .B(KEYINPUT62), .ZN(new_n1063));
  OAI21_X1  g862(.A(G204gat), .B1(new_n1059), .B2(new_n766), .ZN(new_n1064));
  NAND2_X1  g863(.A1(new_n1063), .A2(new_n1064), .ZN(G1353gat));
  INV_X1    g864(.A(new_n1055), .ZN(new_n1066));
  NAND3_X1  g865(.A1(new_n1066), .A2(new_n237), .A3(new_n700), .ZN(new_n1067));
  NAND3_X1  g866(.A1(new_n1058), .A2(new_n700), .A3(new_n1054), .ZN(new_n1068));
  AND3_X1   g867(.A1(new_n1068), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1069));
  AOI21_X1  g868(.A(KEYINPUT63), .B1(new_n1068), .B2(G211gat), .ZN(new_n1070));
  OAI21_X1  g869(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g870(.A(KEYINPUT127), .ZN(new_n1072));
  NAND2_X1  g871(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g872(.A(KEYINPUT127), .B(new_n1067), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g873(.A1(new_n1073), .A2(new_n1074), .ZN(G1354gat));
  OAI21_X1  g874(.A(G218gat), .B1(new_n1059), .B2(new_n738), .ZN(new_n1076));
  NAND3_X1  g875(.A1(new_n1066), .A2(new_n238), .A3(new_n802), .ZN(new_n1077));
  NAND2_X1  g876(.A1(new_n1076), .A2(new_n1077), .ZN(G1355gat));
endmodule


