//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT68), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n188), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(G128), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n198), .B(new_n200), .C1(new_n201), .C2(KEYINPUT23), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT74), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n199), .B2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n197), .A2(KEYINPUT74), .A3(G119), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n200), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n211));
  INV_X1    g025(.A(G125), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n212), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n211), .A2(G146), .A3(new_n213), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n203), .B(new_n209), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n216), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n207), .A2(KEYINPUT75), .A3(new_n208), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(G110), .B2(new_n202), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT75), .B1(new_n207), .B2(new_n208), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n218), .B(new_n220), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT76), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n217), .A2(new_n227), .A3(new_n224), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n196), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n196), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G234), .ZN(new_n235));
  OAI21_X1  g049(.A(G217), .B1(new_n235), .B2(G902), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT79), .B1(new_n229), .B2(new_n231), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n234), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n228), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n227), .B1(new_n217), .B2(new_n224), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n195), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n244), .B2(new_n230), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT25), .B1(new_n245), .B2(KEYINPUT78), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT78), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n247), .B(new_n248), .C1(new_n232), .C2(G902), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(new_n236), .B(KEYINPUT73), .Z(new_n251));
  AOI21_X1  g065(.A(new_n241), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n254));
  INV_X1    g068(.A(G237), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n193), .A2(G210), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n199), .A2(G116), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G119), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT2), .B(G113), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT0), .A3(G128), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT64), .A2(G134), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(G137), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT65), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n276), .A2(new_n280), .A3(G137), .A4(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n283), .A2(new_n275), .A3(G137), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G137), .B1(new_n276), .B2(new_n277), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n285), .B1(new_n286), .B2(KEYINPUT11), .ZN(new_n287));
  OAI21_X1  g101(.A(G131), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G137), .ZN(new_n289));
  AND2_X1   g103(.A1(KEYINPUT64), .A2(G134), .ZN(new_n290));
  NOR2_X1   g104(.A1(KEYINPUT64), .A2(G134), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n284), .B1(new_n292), .B2(new_n283), .ZN(new_n293));
  INV_X1    g107(.A(G131), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n279), .A4(new_n281), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n273), .B1(new_n288), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n275), .A2(G137), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(G143), .B2(new_n219), .ZN(new_n300));
  INV_X1    g114(.A(G143), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(G146), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n219), .A2(G143), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n300), .A2(new_n197), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n219), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n301), .A2(G146), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n299), .A4(G128), .ZN(new_n307));
  AOI22_X1  g121(.A1(G131), .A2(new_n298), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT66), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n295), .A3(KEYINPUT66), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n269), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n288), .A2(new_n295), .ZN(new_n313));
  INV_X1    g127(.A(new_n273), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(new_n295), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n268), .B(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n260), .B1(new_n312), .B2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n308), .A2(new_n295), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n296), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n259), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n296), .A2(new_n321), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n316), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n315), .A2(new_n311), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n329), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n319), .B1(new_n333), .B2(new_n268), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT31), .B1(new_n334), .B2(new_n259), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n315), .A2(KEYINPUT30), .A3(new_n316), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n308), .A2(new_n295), .A3(KEYINPUT66), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n296), .A2(new_n337), .A3(new_n309), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n268), .B(new_n336), .C1(new_n338), .C2(KEYINPUT30), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT31), .A3(new_n259), .A4(new_n323), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n327), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G472), .A2(G902), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(KEYINPUT32), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n339), .A2(new_n259), .A3(new_n323), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT31), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n326), .B1(new_n349), .B2(new_n340), .ZN(new_n350));
  INV_X1    g164(.A(new_n343), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G472), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT71), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n334), .B2(new_n259), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n339), .A2(new_n323), .ZN(new_n358));
  INV_X1    g172(.A(new_n259), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT71), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n332), .A2(new_n268), .B1(new_n322), .B2(new_n318), .ZN(new_n361));
  INV_X1    g175(.A(new_n260), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n259), .B(new_n325), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n356), .A2(new_n357), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n325), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n322), .B(new_n318), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(KEYINPUT28), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n359), .A2(new_n357), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n354), .B1(new_n364), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n254), .B1(new_n353), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n369), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G472), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT72), .A3(new_n344), .A4(new_n352), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n253), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G210), .B1(G237), .B2(G902), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT86), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G104), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT80), .A3(G104), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(KEYINPUT3), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n384), .A3(KEYINPUT80), .A4(G104), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g207(.A(new_n385), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n383), .A4(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n392), .B(new_n268), .C1(new_n390), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G104), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  OAI21_X1  g213(.A(G101), .B1(new_n399), .B2(new_n385), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n199), .A3(G116), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(G113), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n404), .B(new_n405), .C1(new_n402), .C2(new_n264), .ZN(new_n406));
  OAI211_X1 g220(.A(G113), .B(new_n403), .C1(new_n264), .C2(new_n402), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT84), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n401), .A2(new_n406), .A3(new_n266), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n397), .A2(new_n409), .A3(new_n411), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n304), .A2(new_n307), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n212), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n212), .B2(new_n273), .ZN(new_n418));
  INV_X1    g232(.A(G224), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(G953), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n420), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n410), .A2(new_n424), .A3(new_n412), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n415), .A2(KEYINPUT85), .A3(new_n423), .A4(new_n425), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n421), .A2(new_n422), .A3(new_n431), .ZN(new_n432));
  OR3_X1    g246(.A1(new_n418), .A2(KEYINPUT7), .A3(new_n420), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n266), .A2(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n401), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n411), .B(KEYINPUT8), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n408), .A2(new_n266), .A3(new_n406), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n435), .B(new_n436), .C1(new_n437), .C2(new_n401), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n432), .A2(new_n433), .A3(new_n414), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n237), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n382), .B1(new_n430), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n428), .B2(new_n429), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n381), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n378), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT9), .B(G234), .ZN(new_n445));
  OAI21_X1  g259(.A(G221), .B1(new_n445), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n401), .A2(KEYINPUT10), .A3(new_n416), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n392), .B1(new_n390), .B2(new_n396), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n273), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n401), .A2(new_n451), .A3(new_n416), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n304), .A2(new_n307), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n395), .A2(new_n400), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT81), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n452), .A2(new_n455), .A3(new_n459), .A4(new_n456), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n450), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n313), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n452), .B(new_n455), .C1(new_n416), .C2(new_n401), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n313), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(KEYINPUT12), .A3(new_n313), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n193), .A2(G227), .ZN(new_n471));
  XOR2_X1   g285(.A(G110), .B(G140), .Z(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n461), .A2(new_n462), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n461), .B2(new_n462), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n470), .A2(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G469), .B1(new_n476), .B2(G902), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n461), .A2(new_n462), .ZN(new_n478));
  AOI211_X1 g292(.A(new_n313), .B(new_n450), .C1(new_n458), .C2(new_n460), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G469), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n237), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n447), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(G128), .B(G143), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n276), .A2(new_n277), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G116), .B(G122), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n384), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n262), .A2(KEYINPUT14), .A3(G122), .ZN(new_n491));
  XOR2_X1   g305(.A(G116), .B(G122), .Z(new_n492));
  OAI211_X1 g306(.A(G107), .B(new_n491), .C1(new_n492), .C2(KEYINPUT14), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(G107), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n490), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n301), .A3(G128), .ZN(new_n498));
  OAI211_X1 g312(.A(G134), .B(new_n498), .C1(new_n486), .C2(new_n497), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n499), .C1(new_n487), .C2(new_n486), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G217), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n445), .A2(new_n502), .A3(G953), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n500), .A3(new_n503), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n237), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT90), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n505), .B2(new_n506), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G478), .ZN(new_n514));
  NOR2_X1   g328(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n519), .B1(new_n508), .B2(new_n520), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  XNOR2_X1  g339(.A(G113), .B(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n398), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n193), .A2(G214), .A3(new_n255), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n301), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n193), .A2(G143), .A3(G214), .A4(new_n255), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(KEYINPUT87), .A2(KEYINPUT18), .A3(G131), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n210), .A2(new_n219), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n220), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT88), .A3(new_n220), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n534), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n294), .B1(new_n529), .B2(new_n530), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n529), .A2(new_n294), .A3(new_n530), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n215), .A2(new_n216), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n544), .B2(new_n545), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n527), .B(new_n542), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n527), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n534), .A2(new_n540), .A3(new_n541), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n210), .B(KEYINPUT19), .Z(new_n553));
  OAI21_X1  g367(.A(new_n218), .B1(G146), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n544), .B2(new_n546), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT89), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n525), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT20), .B(new_n559), .C1(new_n550), .C2(new_n556), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n542), .B1(new_n547), .B2(new_n549), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n551), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n564), .B2(new_n550), .ZN(new_n565));
  INV_X1    g379(.A(G475), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n561), .A2(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n189), .A2(G952), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n235), .B2(new_n255), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n237), .B(new_n193), .C1(G234), .C2(G237), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT21), .B(G898), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n524), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n444), .A2(new_n485), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n376), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT93), .B(G101), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G3));
  NAND2_X1  g392(.A1(new_n342), .A2(new_n237), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n342), .A2(new_n343), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n485), .A2(new_n252), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n377), .B1(new_n442), .B2(new_n380), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n379), .B(new_n440), .C1(new_n428), .C2(new_n429), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n573), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n514), .A2(G902), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n507), .A2(KEYINPUT33), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n505), .B2(new_n506), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT94), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n509), .A2(new_n514), .A3(new_n512), .ZN(new_n596));
  OAI211_X1 g410(.A(KEYINPUT94), .B(new_n589), .C1(new_n590), .C2(new_n592), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n567), .A2(new_n588), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n584), .A2(new_n587), .A3(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT34), .B(G104), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G6));
  NAND2_X1  g416(.A1(new_n557), .A2(new_n560), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT20), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n557), .A2(new_n525), .A3(new_n560), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(KEYINPUT95), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(KEYINPUT95), .B2(new_n605), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n565), .A2(new_n566), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n524), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n588), .A3(new_n587), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n610), .A2(new_n587), .A3(KEYINPUT96), .A4(new_n588), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n584), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  INV_X1    g432(.A(new_n575), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n580), .A2(new_n581), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n250), .A2(new_n251), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n242), .A2(new_n243), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n195), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n239), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n619), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT37), .B(G110), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G12));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n587), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n570), .B1(new_n571), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n607), .A2(new_n609), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n634), .A2(new_n485), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n345), .B1(new_n342), .B2(new_n343), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT32), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n350), .A2(new_n637), .A3(new_n351), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT72), .B1(new_n639), .B2(new_n373), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n353), .A2(new_n254), .A3(new_n370), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n631), .B(new_n635), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  INV_X1    g457(.A(new_n626), .ZN(new_n644));
  INV_X1    g458(.A(new_n567), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n522), .A2(new_n523), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n647), .A3(new_n377), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n441), .A2(new_n443), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n633), .B(KEYINPUT39), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n485), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n648), .B(new_n651), .C1(KEYINPUT40), .C2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(KEYINPUT40), .B2(new_n653), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n366), .A2(new_n359), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT97), .Z(new_n657));
  INV_X1    g471(.A(new_n347), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n237), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n639), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT98), .Z(new_n662));
  OR2_X1    g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT99), .B(G143), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G45));
  INV_X1    g479(.A(new_n598), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n645), .A2(new_n666), .A3(new_n633), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n485), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n631), .B(new_n668), .C1(new_n640), .C2(new_n641), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT100), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n630), .B1(new_n371), .B2(new_n374), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(new_n668), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  AOI21_X1  g489(.A(new_n483), .B1(new_n482), .B2(new_n237), .ZN(new_n676));
  AOI211_X1 g490(.A(G469), .B(G902), .C1(new_n480), .C2(new_n481), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n678), .A2(new_n587), .A3(new_n599), .A4(new_n446), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n376), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT101), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G15));
  INV_X1    g497(.A(new_n676), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n446), .A3(new_n484), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n613), .B2(new_n614), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n375), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n585), .A2(new_n586), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n689), .B1(new_n685), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n678), .A2(new_n587), .A3(KEYINPUT102), .A4(new_n446), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n691), .A2(new_n574), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n644), .B1(new_n371), .B2(new_n374), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT103), .B(G119), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G21));
  XNOR2_X1  g511(.A(KEYINPUT104), .B(G472), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n579), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g513(.A1(new_n335), .A2(new_n341), .B1(new_n259), .B2(new_n367), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n343), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n253), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n647), .A2(new_n587), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n685), .A2(new_n573), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n703), .A2(new_n708), .A3(new_n704), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND4_X1  g525(.A1(new_n667), .A2(new_n699), .A3(new_n626), .A4(new_n701), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n691), .A3(new_n692), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  NAND3_X1  g529(.A1(new_n441), .A2(new_n377), .A3(new_n443), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n485), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n645), .A2(new_n666), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(KEYINPUT42), .A3(new_n633), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n375), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n668), .A2(new_n717), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n581), .A2(new_n637), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n373), .A3(new_n344), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n252), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT106), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n723), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(G131), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G33));
  NOR2_X1   g549(.A1(new_n376), .A2(new_n718), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n634), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  NAND2_X1  g552(.A1(new_n470), .A2(new_n473), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n474), .A2(new_n475), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n476), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(G469), .A2(G902), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n677), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n447), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n652), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n666), .A2(new_n567), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT43), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n582), .A3(new_n626), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n716), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n752), .B(new_n757), .C1(new_n756), .C2(new_n755), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT108), .B(G137), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G39));
  XNOR2_X1  g574(.A(new_n751), .B(KEYINPUT47), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n717), .A2(new_n253), .A3(new_n667), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n371), .A3(new_n374), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT109), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G140), .ZN(G42));
  INV_X1    g579(.A(new_n678), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n651), .B1(KEYINPUT49), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n377), .A3(new_n446), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n768), .B(new_n253), .C1(KEYINPUT49), .C2(new_n766), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n662), .C1(new_n770), .C2(new_n769), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n685), .A2(new_n569), .A3(new_n716), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n662), .A2(new_n252), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n567), .A2(new_n598), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(KEYINPUT116), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n773), .A2(new_n754), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n644), .A3(new_n702), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n651), .A2(new_n378), .A3(new_n446), .A4(new_n678), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n703), .A2(new_n570), .A3(new_n754), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n785), .B1(new_n783), .B2(new_n784), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n780), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n784), .A2(new_n716), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n766), .A2(new_n446), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT115), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n761), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n761), .B2(new_n792), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n774), .A2(new_n720), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n691), .A2(new_n692), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n784), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n568), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n801), .A2(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(KEYINPUT117), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n781), .A2(new_n727), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT48), .Z(new_n805));
  NAND4_X1  g619(.A1(new_n797), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n626), .A2(new_n633), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n661), .A2(new_n485), .A3(new_n704), .A4(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n642), .A2(new_n714), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n674), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n808), .B1(new_n674), .B2(new_n811), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT114), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n730), .A2(new_n732), .A3(new_n737), .ZN(new_n815));
  AOI221_X4 g629(.A(new_n253), .B1(new_n575), .B2(new_n679), .C1(new_n371), .C2(new_n374), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n567), .A2(new_n646), .A3(new_n573), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n444), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT111), .ZN(new_n819));
  INV_X1    g633(.A(new_n583), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n444), .A2(new_n821), .A3(new_n817), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n620), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n620), .A3(new_n444), .A4(new_n599), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n627), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n816), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n686), .A2(new_n375), .B1(new_n693), .B2(new_n694), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n712), .A2(new_n718), .A3(KEYINPUT112), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT112), .B1(new_n712), .B2(new_n718), .ZN(new_n829));
  INV_X1    g643(.A(new_n633), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n608), .A2(new_n646), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n718), .A2(new_n607), .A3(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n828), .A2(new_n829), .B1(new_n694), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n826), .A2(new_n710), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n671), .A2(new_n672), .A3(new_n668), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n672), .B1(new_n671), .B2(new_n668), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n642), .A2(new_n714), .A3(new_n810), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT52), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n674), .A2(new_n811), .A3(new_n808), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n814), .A2(new_n835), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n642), .A2(new_n714), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT113), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT113), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n642), .A2(new_n847), .A3(new_n714), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n846), .A2(new_n674), .A3(new_n810), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n812), .B1(KEYINPUT52), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n815), .A2(new_n834), .A3(KEYINPUT53), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n844), .A2(KEYINPUT53), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n737), .A2(KEYINPUT53), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n834), .A2(new_n857), .A3(new_n729), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n807), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n861), .A2(new_n862), .B1(G952), .B2(G953), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n772), .B1(new_n863), .B2(new_n864), .ZN(G75));
  NOR2_X1   g679(.A1(new_n193), .A2(G952), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT120), .Z(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n415), .A2(new_n425), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n423), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n237), .B1(new_n855), .B2(new_n859), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n873), .B(new_n876), .C1(new_n874), .C2(new_n871), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n868), .B1(new_n878), .B2(new_n879), .ZN(G51));
  INV_X1    g694(.A(new_n866), .ZN(new_n881));
  INV_X1    g695(.A(new_n482), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n855), .A2(new_n859), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n860), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n746), .B(KEYINPUT57), .Z(new_n886));
  AOI21_X1  g700(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n237), .B(new_n745), .C1(new_n855), .C2(new_n859), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT121), .B(new_n881), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n890));
  AOI221_X4 g704(.A(KEYINPUT54), .B1(new_n850), .B2(new_n858), .C1(new_n844), .C2(new_n854), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n856), .B1(new_n855), .B2(new_n859), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n893), .B2(new_n482), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n890), .B1(new_n894), .B2(new_n866), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n889), .A2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n898));
  INV_X1    g712(.A(new_n557), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n881), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  NOR2_X1   g717(.A1(new_n590), .A2(new_n592), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT123), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n853), .A2(new_n860), .ZN(new_n906));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT59), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n905), .A2(new_n908), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n868), .B(new_n909), .C1(new_n885), .C2(new_n910), .ZN(G63));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT60), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n883), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n234), .A2(new_n240), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n624), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n916), .B(new_n867), .C1(new_n917), .C2(new_n914), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G66));
  OAI21_X1  g734(.A(G953), .B1(new_n572), .B2(new_n419), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n826), .A2(new_n710), .A3(new_n827), .ZN(new_n922));
  INV_X1    g736(.A(new_n193), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(G898), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n869), .B1(new_n925), .B2(new_n923), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n924), .B(new_n926), .Z(G69));
  XOR2_X1   g741(.A(new_n333), .B(new_n553), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n193), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n524), .B(new_n608), .C1(new_n561), .C2(new_n562), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n716), .B(new_n653), .C1(new_n721), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n375), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n764), .A2(new_n758), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n846), .A2(new_n674), .A3(new_n848), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n663), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n934), .A2(new_n937), .A3(KEYINPUT124), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n930), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n193), .A2(G900), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n928), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n752), .A2(new_n252), .A3(new_n704), .A4(new_n726), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n758), .A2(new_n764), .A3(new_n935), .A4(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n815), .A2(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n815), .A2(KEYINPUT126), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n952), .B2(new_n193), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n944), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n944), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n942), .B2(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(G72));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  NAND3_X1  g774(.A1(new_n356), .A2(new_n347), .A3(new_n360), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n852), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n949), .A2(new_n922), .A3(new_n950), .A4(new_n951), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n960), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n358), .B(KEYINPUT127), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(new_n259), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n881), .B(new_n962), .C1(new_n964), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n259), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n940), .A2(new_n922), .A3(new_n941), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n960), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n967), .A2(new_n970), .ZN(G57));
endmodule


