

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n641), .ZN(n607) );
  XNOR2_X1 U550 ( .A(n539), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X1 U551 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X2 U552 ( .A1(n525), .A2(G2105), .ZN(n711) );
  XNOR2_X2 U553 ( .A(n642), .B(n588), .ZN(n641) );
  INV_X1 U554 ( .A(KEYINPUT28), .ZN(n600) );
  NOR2_X1 U555 ( .A1(n646), .A2(n645), .ZN(n648) );
  NAND2_X1 U556 ( .A1(n518), .A2(n709), .ZN(n747) );
  NAND2_X1 U557 ( .A1(n708), .A2(KEYINPUT96), .ZN(n709) );
  AND2_X1 U558 ( .A1(n746), .A2(n745), .ZN(n517) );
  AND2_X1 U559 ( .A1(n701), .A2(n700), .ZN(n518) );
  INV_X1 U560 ( .A(KEYINPUT94), .ZN(n647) );
  BUF_X1 U561 ( .A(n605), .Z(n656) );
  XNOR2_X1 U562 ( .A(G2104), .B(KEYINPUT66), .ZN(n521) );
  INV_X1 U563 ( .A(n752), .ZN(n745) );
  XNOR2_X1 U564 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n724) );
  AND2_X1 U566 ( .A1(G2105), .A2(n525), .ZN(n887) );
  NOR2_X1 U567 ( .A1(G651), .A2(n570), .ZN(n788) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n792) );
  XOR2_X1 U569 ( .A(KEYINPUT81), .B(n530), .Z(G164) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n520), .B(n519), .ZN(n531) );
  NAND2_X1 U572 ( .A1(G138), .A2(n531), .ZN(n523) );
  INV_X1 U573 ( .A(n521), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n711), .A2(G102), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U576 ( .A(KEYINPUT80), .B(n524), .ZN(n529) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U578 ( .A1(G114), .A2(n886), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G126), .A2(n887), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  BUF_X1 U581 ( .A(n531), .Z(n891) );
  NAND2_X1 U582 ( .A1(n891), .A2(G137), .ZN(n538) );
  NAND2_X1 U583 ( .A1(G113), .A2(n886), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G125), .A2(n887), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U586 ( .A1(G101), .A2(n711), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT23), .B(n534), .ZN(n535) );
  NOR2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n570) );
  INV_X1 U591 ( .A(G651), .ZN(n543) );
  NOR2_X1 U592 ( .A1(n570), .A2(n543), .ZN(n791) );
  NAND2_X1 U593 ( .A1(G77), .A2(n791), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G90), .A2(n792), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U596 ( .A(KEYINPUT9), .B(n542), .ZN(n548) );
  NOR2_X1 U597 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U598 ( .A(KEYINPUT1), .B(n544), .Z(n787) );
  NAND2_X1 U599 ( .A1(G64), .A2(n787), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G52), .A2(n788), .ZN(n545) );
  AND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(G301) );
  NAND2_X1 U603 ( .A1(G63), .A2(n787), .ZN(n550) );
  NAND2_X1 U604 ( .A1(G51), .A2(n788), .ZN(n549) );
  NAND2_X1 U605 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U606 ( .A(KEYINPUT6), .B(n551), .ZN(n558) );
  NAND2_X1 U607 ( .A1(n792), .A2(G89), .ZN(n552) );
  XNOR2_X1 U608 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G76), .A2(n791), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT5), .B(n555), .ZN(n556) );
  XNOR2_X1 U612 ( .A(KEYINPUT71), .B(n556), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(n559), .Z(G168) );
  NAND2_X1 U615 ( .A1(G75), .A2(n791), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G88), .A2(n792), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U618 ( .A1(G62), .A2(n787), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G50), .A2(n788), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n565), .A2(n564), .ZN(G166) );
  XOR2_X1 U622 ( .A(KEYINPUT82), .B(G166), .Z(G303) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G49), .A2(n788), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U627 ( .A(KEYINPUT73), .B(n568), .Z(n569) );
  NOR2_X1 U628 ( .A1(n787), .A2(n569), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n570), .A2(G87), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(G288) );
  NAND2_X1 U631 ( .A1(G61), .A2(n787), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G48), .A2(n788), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G73), .A2(n791), .ZN(n575) );
  XOR2_X1 U635 ( .A(KEYINPUT2), .B(n575), .Z(n576) );
  NOR2_X1 U636 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n792), .A2(G86), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n579), .A2(n578), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G72), .A2(n791), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G85), .A2(n792), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n787), .A2(G60), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n582), .Z(n583) );
  NOR2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n788), .A2(G47), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n586), .A2(n585), .ZN(G290) );
  NAND2_X1 U647 ( .A1(G160), .A2(G40), .ZN(n723) );
  INV_X1 U648 ( .A(n723), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n587), .A2(n724), .ZN(n605) );
  INV_X2 U650 ( .A(n605), .ZN(n642) );
  INV_X1 U651 ( .A(KEYINPUT90), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G1956), .A2(n641), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G2072), .A2(n607), .ZN(n589) );
  XNOR2_X1 U654 ( .A(KEYINPUT27), .B(n589), .ZN(n590) );
  INV_X1 U655 ( .A(n590), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT91), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G65), .A2(n787), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G53), .A2(n788), .ZN(n594) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G78), .A2(n791), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G91), .A2(n792), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n975) );
  NOR2_X1 U665 ( .A1(n602), .A2(n975), .ZN(n601) );
  XNOR2_X1 U666 ( .A(n601), .B(n600), .ZN(n639) );
  NAND2_X1 U667 ( .A1(n602), .A2(n975), .ZN(n637) );
  NAND2_X1 U668 ( .A1(G1996), .A2(n642), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT26), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT64), .B(n604), .ZN(n618) );
  NAND2_X1 U671 ( .A1(G1348), .A2(n656), .ZN(n606) );
  XOR2_X1 U672 ( .A(KEYINPUT93), .B(n606), .Z(n609) );
  NAND2_X1 U673 ( .A1(G2067), .A2(n607), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n633) );
  NAND2_X1 U675 ( .A1(G79), .A2(n791), .ZN(n611) );
  NAND2_X1 U676 ( .A1(G54), .A2(n788), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U678 ( .A1(G66), .A2(n787), .ZN(n613) );
  NAND2_X1 U679 ( .A1(G92), .A2(n792), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U681 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U682 ( .A(n616), .B(KEYINPUT15), .Z(n989) );
  INV_X1 U683 ( .A(n989), .ZN(n766) );
  NAND2_X1 U684 ( .A1(n633), .A2(n766), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n632) );
  NAND2_X1 U686 ( .A1(n656), .A2(G1341), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n619), .B(KEYINPUT92), .ZN(n630) );
  XOR2_X1 U688 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n621) );
  NAND2_X1 U689 ( .A1(G56), .A2(n787), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n621), .B(n620), .ZN(n629) );
  NAND2_X1 U691 ( .A1(n792), .A2(G81), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n622), .B(KEYINPUT12), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G68), .A2(n791), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT13), .ZN(n627) );
  NAND2_X1 U696 ( .A1(G43), .A2(n788), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n980) );
  NAND2_X1 U699 ( .A1(n630), .A2(n980), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n633), .A2(n766), .ZN(n634) );
  NOR2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U705 ( .A(n640), .B(KEYINPUT29), .ZN(n646) );
  XOR2_X1 U706 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U707 ( .A1(n929), .A2(n641), .ZN(n644) );
  NOR2_X1 U708 ( .A1(n642), .A2(G1961), .ZN(n643) );
  NOR2_X1 U709 ( .A1(n644), .A2(n643), .ZN(n649) );
  NOR2_X1 U710 ( .A1(G301), .A2(n649), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n648), .B(n647), .ZN(n669) );
  AND2_X1 U712 ( .A1(G301), .A2(n649), .ZN(n654) );
  NAND2_X1 U713 ( .A1(n656), .A2(G8), .ZN(n689) );
  NOR2_X1 U714 ( .A1(G1966), .A2(n689), .ZN(n671) );
  NOR2_X1 U715 ( .A1(G2084), .A2(n656), .ZN(n670) );
  NOR2_X1 U716 ( .A1(n671), .A2(n670), .ZN(n650) );
  NAND2_X1 U717 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U718 ( .A(KEYINPUT30), .B(n651), .ZN(n652) );
  NOR2_X1 U719 ( .A1(G168), .A2(n652), .ZN(n653) );
  NOR2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT31), .B(n655), .Z(n668) );
  INV_X1 U722 ( .A(G8), .ZN(n661) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n689), .ZN(n658) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n656), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U726 ( .A1(G303), .A2(n659), .ZN(n660) );
  OR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n663) );
  AND2_X1 U728 ( .A1(n668), .A2(n663), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n669), .A2(n662), .ZN(n666) );
  INV_X1 U730 ( .A(n663), .ZN(n664) );
  OR2_X1 U731 ( .A1(n664), .A2(G286), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT32), .ZN(n676) );
  AND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n674) );
  AND2_X1 U735 ( .A1(G8), .A2(n670), .ZN(n672) );
  OR2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  OR2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n678) );
  INV_X1 U739 ( .A(KEYINPUT95), .ZN(n677) );
  XNOR2_X2 U740 ( .A(n678), .B(n677), .ZN(n703) );
  NOR2_X1 U741 ( .A1(G2090), .A2(G303), .ZN(n679) );
  NAND2_X1 U742 ( .A1(G8), .A2(n679), .ZN(n680) );
  NAND2_X1 U743 ( .A1(n703), .A2(n680), .ZN(n681) );
  NAND2_X1 U744 ( .A1(n681), .A2(n689), .ZN(n707) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n687), .A2(n682), .ZN(n974) );
  INV_X1 U748 ( .A(KEYINPUT33), .ZN(n683) );
  AND2_X1 U749 ( .A1(n974), .A2(n683), .ZN(n702) );
  INV_X1 U750 ( .A(KEYINPUT96), .ZN(n684) );
  AND2_X1 U751 ( .A1(n702), .A2(n684), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n703), .A2(n685), .ZN(n695) );
  INV_X1 U753 ( .A(n689), .ZN(n698) );
  NAND2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n978) );
  AND2_X1 U755 ( .A1(n698), .A2(n978), .ZN(n686) );
  OR2_X1 U756 ( .A1(KEYINPUT33), .A2(n686), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  OR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n693) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n985) );
  INV_X1 U761 ( .A(n985), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n704) );
  OR2_X1 U763 ( .A1(KEYINPUT96), .A2(n704), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n707), .A2(n696), .ZN(n701) );
  NOR2_X1 U766 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n697), .B(KEYINPUT24), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U772 ( .A(G1986), .B(G290), .Z(n979) );
  XOR2_X1 U773 ( .A(G2067), .B(KEYINPUT37), .Z(n710) );
  XNOR2_X1 U774 ( .A(KEYINPUT83), .B(n710), .ZN(n748) );
  XNOR2_X1 U775 ( .A(KEYINPUT84), .B(KEYINPUT34), .ZN(n715) );
  BUF_X1 U776 ( .A(n711), .Z(n890) );
  NAND2_X1 U777 ( .A1(G104), .A2(n890), .ZN(n713) );
  NAND2_X1 U778 ( .A1(G140), .A2(n891), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(n715), .B(n714), .ZN(n720) );
  NAND2_X1 U781 ( .A1(G116), .A2(n886), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G128), .A2(n887), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U784 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(KEYINPUT36), .B(n721), .ZN(n877) );
  NOR2_X1 U787 ( .A1(n748), .A2(n877), .ZN(n722) );
  XNOR2_X1 U788 ( .A(n722), .B(KEYINPUT85), .ZN(n1011) );
  NAND2_X1 U789 ( .A1(n979), .A2(n1011), .ZN(n725) );
  NOR2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n758) );
  NAND2_X1 U791 ( .A1(n725), .A2(n758), .ZN(n746) );
  NAND2_X1 U792 ( .A1(n887), .A2(G119), .ZN(n726) );
  XNOR2_X1 U793 ( .A(n726), .B(KEYINPUT86), .ZN(n728) );
  NAND2_X1 U794 ( .A1(G107), .A2(n886), .ZN(n727) );
  NAND2_X1 U795 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U796 ( .A(KEYINPUT87), .B(n729), .ZN(n733) );
  NAND2_X1 U797 ( .A1(n890), .A2(G95), .ZN(n731) );
  NAND2_X1 U798 ( .A1(G131), .A2(n891), .ZN(n730) );
  AND2_X1 U799 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U800 ( .A1(n733), .A2(n732), .ZN(n868) );
  NAND2_X1 U801 ( .A1(G1991), .A2(n868), .ZN(n734) );
  XNOR2_X1 U802 ( .A(n734), .B(KEYINPUT88), .ZN(n743) );
  NAND2_X1 U803 ( .A1(G141), .A2(n891), .ZN(n736) );
  NAND2_X1 U804 ( .A1(G117), .A2(n886), .ZN(n735) );
  NAND2_X1 U805 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U806 ( .A1(n890), .A2(G105), .ZN(n737) );
  XOR2_X1 U807 ( .A(KEYINPUT38), .B(n737), .Z(n738) );
  NOR2_X1 U808 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U809 ( .A1(n887), .A2(G129), .ZN(n740) );
  NAND2_X1 U810 ( .A1(n741), .A2(n740), .ZN(n872) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n872), .ZN(n742) );
  NAND2_X1 U812 ( .A1(n743), .A2(n742), .ZN(n1013) );
  NAND2_X1 U813 ( .A1(n758), .A2(n1013), .ZN(n744) );
  XNOR2_X1 U814 ( .A(KEYINPUT89), .B(n744), .ZN(n752) );
  NAND2_X1 U815 ( .A1(n747), .A2(n517), .ZN(n761) );
  NAND2_X1 U816 ( .A1(n877), .A2(n748), .ZN(n1010) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n872), .ZN(n1019) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n868), .ZN(n749) );
  XOR2_X1 U820 ( .A(KEYINPUT97), .B(n749), .Z(n1006) );
  NOR2_X1 U821 ( .A1(n750), .A2(n1006), .ZN(n751) );
  NOR2_X1 U822 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U823 ( .A1(n1019), .A2(n753), .ZN(n754) );
  XNOR2_X1 U824 ( .A(KEYINPUT39), .B(n754), .ZN(n755) );
  XNOR2_X1 U825 ( .A(n755), .B(KEYINPUT98), .ZN(n756) );
  NAND2_X1 U826 ( .A1(n756), .A2(n1011), .ZN(n757) );
  NAND2_X1 U827 ( .A1(n1010), .A2(n757), .ZN(n759) );
  NAND2_X1 U828 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U829 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U830 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(n975), .ZN(G299) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  INV_X1 U834 ( .A(G132), .ZN(G219) );
  INV_X1 U835 ( .A(G82), .ZN(G220) );
  NAND2_X1 U836 ( .A1(G7), .A2(G661), .ZN(n763) );
  XOR2_X1 U837 ( .A(n763), .B(KEYINPUT10), .Z(n828) );
  NAND2_X1 U838 ( .A1(n828), .A2(G567), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT11), .ZN(n765) );
  XNOR2_X1 U840 ( .A(KEYINPUT69), .B(n765), .ZN(G234) );
  NAND2_X1 U841 ( .A1(n980), .A2(G860), .ZN(G153) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U843 ( .A(G868), .ZN(n776) );
  NAND2_X1 U844 ( .A1(n766), .A2(n776), .ZN(n767) );
  NAND2_X1 U845 ( .A1(n768), .A2(n767), .ZN(G284) );
  NOR2_X1 U846 ( .A1(G286), .A2(n776), .ZN(n770) );
  NOR2_X1 U847 ( .A1(G868), .A2(G299), .ZN(n769) );
  NOR2_X1 U848 ( .A1(n770), .A2(n769), .ZN(G297) );
  INV_X1 U849 ( .A(G860), .ZN(n771) );
  NAND2_X1 U850 ( .A1(n771), .A2(G559), .ZN(n772) );
  NAND2_X1 U851 ( .A1(n772), .A2(n989), .ZN(n773) );
  XNOR2_X1 U852 ( .A(n773), .B(KEYINPUT72), .ZN(n774) );
  XNOR2_X1 U853 ( .A(KEYINPUT16), .B(n774), .ZN(G148) );
  NAND2_X1 U854 ( .A1(n989), .A2(G868), .ZN(n775) );
  NOR2_X1 U855 ( .A1(G559), .A2(n775), .ZN(n778) );
  AND2_X1 U856 ( .A1(n776), .A2(n980), .ZN(n777) );
  NOR2_X1 U857 ( .A1(n778), .A2(n777), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G135), .A2(n891), .ZN(n780) );
  NAND2_X1 U859 ( .A1(G111), .A2(n886), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n780), .A2(n779), .ZN(n785) );
  NAND2_X1 U861 ( .A1(G123), .A2(n887), .ZN(n781) );
  XNOR2_X1 U862 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U863 ( .A1(n890), .A2(G99), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U865 ( .A1(n785), .A2(n784), .ZN(n1005) );
  XNOR2_X1 U866 ( .A(n1005), .B(G2096), .ZN(n786) );
  INV_X1 U867 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U868 ( .A1(n786), .A2(n852), .ZN(G156) );
  NAND2_X1 U869 ( .A1(G67), .A2(n787), .ZN(n790) );
  NAND2_X1 U870 ( .A1(G55), .A2(n788), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U872 ( .A1(G80), .A2(n791), .ZN(n794) );
  NAND2_X1 U873 ( .A1(G93), .A2(n792), .ZN(n793) );
  NAND2_X1 U874 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U875 ( .A1(n796), .A2(n795), .ZN(n811) );
  NAND2_X1 U876 ( .A1(n989), .A2(G559), .ZN(n809) );
  XOR2_X1 U877 ( .A(n980), .B(n809), .Z(n797) );
  NOR2_X1 U878 ( .A1(G860), .A2(n797), .ZN(n798) );
  XNOR2_X1 U879 ( .A(n811), .B(n798), .ZN(G145) );
  XOR2_X1 U880 ( .A(KEYINPUT19), .B(KEYINPUT74), .Z(n800) );
  XNOR2_X1 U881 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n799) );
  XNOR2_X1 U882 ( .A(n800), .B(n799), .ZN(n801) );
  XOR2_X1 U883 ( .A(n801), .B(KEYINPUT75), .Z(n803) );
  XOR2_X1 U884 ( .A(G299), .B(n811), .Z(n802) );
  XNOR2_X1 U885 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U886 ( .A(n980), .B(n804), .ZN(n806) );
  XNOR2_X1 U887 ( .A(G288), .B(G166), .ZN(n805) );
  XNOR2_X1 U888 ( .A(n806), .B(n805), .ZN(n807) );
  XOR2_X1 U889 ( .A(n807), .B(G305), .Z(n808) );
  XNOR2_X1 U890 ( .A(G290), .B(n808), .ZN(n901) );
  XNOR2_X1 U891 ( .A(n809), .B(n901), .ZN(n810) );
  NAND2_X1 U892 ( .A1(n810), .A2(G868), .ZN(n813) );
  OR2_X1 U893 ( .A1(n811), .A2(G868), .ZN(n812) );
  NAND2_X1 U894 ( .A1(n813), .A2(n812), .ZN(G295) );
  XNOR2_X1 U895 ( .A(KEYINPUT20), .B(KEYINPUT79), .ZN(n816) );
  NAND2_X1 U896 ( .A1(G2084), .A2(G2078), .ZN(n814) );
  XNOR2_X1 U897 ( .A(n814), .B(KEYINPUT78), .ZN(n815) );
  XNOR2_X1 U898 ( .A(n816), .B(n815), .ZN(n817) );
  NAND2_X1 U899 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U900 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U901 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U902 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U903 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U905 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G96), .A2(n822), .ZN(n832) );
  NAND2_X1 U907 ( .A1(n832), .A2(G2106), .ZN(n826) );
  NAND2_X1 U908 ( .A1(G69), .A2(G120), .ZN(n823) );
  NOR2_X1 U909 ( .A1(G237), .A2(n823), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G108), .A2(n824), .ZN(n833) );
  NAND2_X1 U911 ( .A1(n833), .A2(G567), .ZN(n825) );
  NAND2_X1 U912 ( .A1(n826), .A2(n825), .ZN(n834) );
  NAND2_X1 U913 ( .A1(G483), .A2(G661), .ZN(n827) );
  NOR2_X1 U914 ( .A1(n834), .A2(n827), .ZN(n831) );
  NAND2_X1 U915 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n828), .ZN(G217) );
  INV_X1 U917 ( .A(n828), .ZN(G223) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n834), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT41), .B(G1991), .Z(n836) );
  XNOR2_X1 U930 ( .A(G1981), .B(G1996), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U932 ( .A(n837), .B(KEYINPUT103), .Z(n839) );
  XNOR2_X1 U933 ( .A(G1971), .B(G1986), .ZN(n838) );
  XNOR2_X1 U934 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U935 ( .A(G1956), .B(G1961), .Z(n841) );
  XNOR2_X1 U936 ( .A(G1976), .B(G1966), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U938 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U939 ( .A(KEYINPUT104), .B(G2474), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2678), .Z(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(KEYINPUT101), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U944 ( .A(KEYINPUT102), .B(G2090), .Z(n849) );
  XNOR2_X1 U945 ( .A(G2072), .B(G2067), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U947 ( .A(n851), .B(n850), .Z(n854) );
  XOR2_X1 U948 ( .A(G2096), .B(n852), .Z(n853) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U950 ( .A(G2084), .B(G2078), .Z(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U952 ( .A1(G100), .A2(n890), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G112), .A2(n886), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U955 ( .A1(n887), .A2(G124), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G136), .A2(n891), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U959 ( .A(KEYINPUT105), .B(n862), .Z(n863) );
  NOR2_X1 U960 ( .A1(n864), .A2(n863), .ZN(G162) );
  XOR2_X1 U961 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n866) );
  XNOR2_X1 U962 ( .A(n1005), .B(KEYINPUT109), .ZN(n865) );
  XNOR2_X1 U963 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U964 ( .A(KEYINPUT48), .B(n867), .ZN(n870) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT106), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n872), .B(n871), .ZN(n874) );
  XNOR2_X1 U968 ( .A(G160), .B(G164), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U970 ( .A(G162), .B(n875), .Z(n876) );
  XNOR2_X1 U971 ( .A(n877), .B(n876), .ZN(n899) );
  NAND2_X1 U972 ( .A1(G103), .A2(n890), .ZN(n879) );
  NAND2_X1 U973 ( .A1(G139), .A2(n891), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U975 ( .A(KEYINPUT107), .B(n880), .Z(n885) );
  NAND2_X1 U976 ( .A1(G115), .A2(n886), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G127), .A2(n887), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n1014) );
  NAND2_X1 U981 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U982 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U983 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U984 ( .A1(G106), .A2(n890), .ZN(n893) );
  NAND2_X1 U985 ( .A1(G142), .A2(n891), .ZN(n892) );
  NAND2_X1 U986 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U987 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U988 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U989 ( .A(n1014), .B(n897), .Z(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U991 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U992 ( .A(G286), .B(n989), .Z(n902) );
  XNOR2_X1 U993 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U994 ( .A(n903), .B(G301), .Z(n904) );
  NOR2_X1 U995 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U996 ( .A(KEYINPUT110), .B(n905), .ZN(G397) );
  XNOR2_X1 U997 ( .A(G2451), .B(G2427), .ZN(n915) );
  XOR2_X1 U998 ( .A(G2430), .B(G2443), .Z(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT99), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1001 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1004 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2446), .B(KEYINPUT100), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n915), .B(n914), .ZN(n916) );
  NAND2_X1 U1008 ( .A1(n916), .A2(G14), .ZN(n922) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G301), .ZN(G171) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n922), .ZN(G401) );
  XOR2_X1 U1019 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n1035) );
  INV_X1 U1020 ( .A(KEYINPUT55), .ZN(n1028) );
  XOR2_X1 U1021 ( .A(G1996), .B(G32), .Z(n928) );
  XOR2_X1 U1022 ( .A(G2072), .B(G33), .Z(n923) );
  XNOR2_X1 U1023 ( .A(KEYINPUT115), .B(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G26), .B(G2067), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT116), .B(n926), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n932) );
  XOR2_X1 U1028 ( .A(G27), .B(n929), .Z(n930) );
  XNOR2_X1 U1029 ( .A(KEYINPUT117), .B(n930), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(KEYINPUT118), .B(n933), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n934), .A2(G28), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(G25), .B(G1991), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT114), .B(n935), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1036 ( .A(KEYINPUT53), .B(n938), .Z(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n939), .B(G34), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(G2084), .B(n940), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G35), .B(G2090), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1043 ( .A(n1028), .B(n945), .Z(n947) );
  INV_X1 U1044 ( .A(G29), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(G11), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n949), .ZN(n1003) );
  XOR2_X1 U1048 ( .A(G4), .B(KEYINPUT124), .Z(n951) );
  XNOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT59), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(n951), .B(n950), .ZN(n958) );
  XOR2_X1 U1051 ( .A(G1981), .B(G6), .Z(n955) );
  XNOR2_X1 U1052 ( .A(G1956), .B(G20), .ZN(n953) );
  XNOR2_X1 U1053 ( .A(G19), .B(G1341), .ZN(n952) );
  NOR2_X1 U1054 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1056 ( .A(KEYINPUT123), .B(n956), .Z(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(KEYINPUT60), .B(n959), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n961) );
  XNOR2_X1 U1060 ( .A(G5), .B(G1961), .ZN(n960) );
  NOR2_X1 U1061 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G1976), .B(G23), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n964) );
  NOR2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n966) );
  NAND2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n968), .ZN(n969) );
  NOR2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1070 ( .A(KEYINPUT61), .B(n971), .Z(n972) );
  NOR2_X1 U1071 ( .A1(G16), .A2(n972), .ZN(n1000) );
  XOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .Z(n998) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1075 ( .A(G1956), .B(n975), .Z(n976) );
  NOR2_X1 U1076 ( .A1(n977), .A2(n976), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1078 ( .A(n980), .B(G1341), .Z(n981) );
  NOR2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(n987), .B(KEYINPUT57), .ZN(n993) );
  XOR2_X1 U1084 ( .A(G301), .B(G1961), .Z(n988) );
  XNOR2_X1 U1085 ( .A(n988), .B(KEYINPUT121), .ZN(n991) );
  XOR2_X1 U1086 ( .A(G1348), .B(n989), .Z(n990) );
  NOR2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(n996), .B(KEYINPUT122), .ZN(n997) );
  NOR2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1093 ( .A(n1001), .B(KEYINPUT125), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1033) );
  XOR2_X1 U1095 ( .A(G160), .B(G2084), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(KEYINPUT111), .B(n1004), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT112), .B(n1009), .ZN(n1026) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1024) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1014), .Z(n1016) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1017), .Z(n1022) );
  XOR2_X1 U1106 ( .A(G2090), .B(G162), .Z(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT51), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT113), .B(n1031), .Z(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(n1035), .B(n1034), .ZN(n1036) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

