//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n632, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  XOR2_X1   g043(.A(new_n468), .B(KEYINPUT67), .Z(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n462), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT68), .B1(new_n462), .B2(G2104), .ZN(new_n472));
  OR2_X1    g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n471), .A2(new_n472), .ZN(new_n478));
  INV_X1    g053(.A(G101), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n475), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n470), .B1(new_n476), .B2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n465), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n465), .A2(new_n462), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n462), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT70), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n493));
  OAI211_X1 g068(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(KEYINPUT72), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(G88), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT71), .B(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n506), .B(new_n507), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n515));
  OAI221_X1 g090(.A(new_n512), .B1(new_n513), .B2(new_n508), .C1(new_n514), .C2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  AOI211_X1 g092(.A(KEYINPUT74), .B(new_n501), .C1(new_n504), .C2(new_n505), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(new_n505), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n515), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n506), .B1(new_n510), .B2(new_n511), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n524), .A2(new_n526), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n508), .ZN(new_n535));
  OAI211_X1 g110(.A(G52), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n536));
  OAI211_X1 g111(.A(G90), .B(new_n506), .C1(new_n510), .C2(new_n511), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n538), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  OAI211_X1 g118(.A(G43), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n544));
  OAI211_X1 g119(.A(G81), .B(new_n506), .C1(new_n510), .C2(new_n511), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n500), .A2(KEYINPUT72), .A3(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT72), .B1(new_n500), .B2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n521), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT74), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n506), .A2(new_n519), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(G56), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n508), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI211_X1 g131(.A(KEYINPUT76), .B(new_n508), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT77), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n553), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n523), .B2(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT76), .B1(new_n560), .B2(new_n508), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n554), .A2(new_n555), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n546), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(new_n528), .A2(G91), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(KEYINPUT78), .B2(KEYINPUT9), .ZN(new_n573));
  OAI211_X1 g148(.A(G543), .B(new_n573), .C1(new_n510), .C2(new_n511), .ZN(new_n574));
  NOR2_X1   g149(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(G78), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G65), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n549), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(G651), .A3(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n574), .A2(new_n575), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(G299));
  INV_X1    g160(.A(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n550), .A2(new_n551), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G49), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n515), .B1(new_n527), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n549), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n508), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n528), .A2(G86), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n596), .A2(KEYINPUT80), .A3(new_n597), .ZN(new_n602));
  OAI211_X1 g177(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(G305));
  AOI22_X1  g179(.A1(G47), .A2(new_n525), .B1(new_n528), .B2(G85), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n606), .B(new_n607), .C1(new_n587), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(new_n597), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n523), .A2(G60), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n606), .B1(new_n611), .B2(new_n607), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n610), .B2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n527), .A2(KEYINPUT82), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT82), .B1(new_n527), .B2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n586), .B1(new_n621), .B2(KEYINPUT83), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n622), .A2(new_n623), .B1(G54), .B2(new_n525), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n625));
  AND3_X1   g200(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n614), .B1(new_n626), .B2(G868), .ZN(G321));
  XNOR2_X1  g202(.A(G321), .B(KEYINPUT84), .ZN(G284));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n581), .A2(G651), .A3(new_n582), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n584), .A2(new_n571), .A3(new_n576), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n629), .B1(new_n632), .B2(G868), .ZN(G297));
  OAI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(G868), .ZN(G280));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n626), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n626), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g215(.A1(new_n478), .A2(new_n465), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT85), .B(KEYINPUT13), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n484), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n486), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n462), .A2(G111), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n646), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2427), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT15), .B(G2435), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n658), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n671), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n678), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(new_n687), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n689), .B(new_n692), .C1(new_n684), .C2(new_n688), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT89), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G35), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n704), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2090), .ZN(new_n708));
  INV_X1    g283(.A(new_n704), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G26), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT28), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n484), .A2(G140), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT93), .ZN(new_n713));
  OAI21_X1  g288(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n714));
  INV_X1    g289(.A(G116), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G2105), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n486), .B2(G128), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT24), .B(G34), .ZN(new_n723));
  AOI22_X1  g298(.A1(G160), .A2(G29), .B1(new_n709), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n721), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n704), .A2(G27), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G164), .B2(new_n704), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2078), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G2084), .B2(new_n724), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NOR2_X1   g306(.A1(G5), .A2(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n733), .B(new_n734), .C1(G301), .C2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n726), .B(new_n730), .C1(new_n731), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n701), .A2(G33), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n484), .A2(G139), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT94), .Z(new_n740));
  NAND2_X1  g315(.A1(G115), .A2(G2104), .ZN(new_n741));
  INV_X1    g316(.A(G127), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n465), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  NAND2_X1  g319(.A1(G103), .A2(G2104), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G2105), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n743), .A2(G2105), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n738), .B1(new_n750), .B2(new_n701), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  NOR2_X1   g327(.A1(G168), .A2(new_n735), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n735), .B2(G21), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n473), .A2(G105), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n484), .A2(G141), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n486), .A2(G129), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND4_X1  g336(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(new_n701), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n701), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT31), .B(G11), .Z(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n701), .B1(new_n770), .B2(G28), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT95), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n772), .A2(KEYINPUT95), .B1(new_n770), .B2(G28), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n651), .B2(new_n709), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n767), .A2(new_n768), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n752), .A2(new_n756), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n754), .A2(new_n755), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n737), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n708), .B(new_n780), .C1(new_n731), .C2(new_n736), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n735), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n565), .B2(new_n735), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G1341), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G1341), .ZN(new_n785));
  NOR2_X1   g360(.A1(G4), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n626), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1348), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n735), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT23), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT97), .B(G1956), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n781), .A2(new_n784), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n735), .A2(G24), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT90), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G290), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT91), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1986), .Z(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT92), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n735), .A2(G22), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n735), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n735), .A2(G23), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n589), .A2(new_n592), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n735), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT33), .B(G1976), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n804), .A2(new_n808), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n484), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n486), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(new_n704), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n823), .B(new_n824), .Z(new_n825));
  NAND4_X1  g400(.A1(new_n800), .A2(new_n816), .A3(new_n817), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT36), .Z(new_n827));
  NOR2_X1   g402(.A1(new_n795), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n626), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT99), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(KEYINPUT38), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n836), .A2(new_n515), .B1(new_n527), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n587), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n841), .B2(new_n597), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n556), .B2(new_n557), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g420(.A(KEYINPUT98), .B(new_n842), .C1(new_n556), .C2(new_n557), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n842), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n558), .A2(new_n564), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n834), .A2(new_n835), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n834), .B2(new_n835), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n831), .ZN(new_n855));
  AOI211_X1 g430(.A(KEYINPUT100), .B(KEYINPUT39), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n830), .B1(new_n831), .B2(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n842), .A2(new_n830), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n718), .B(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n497), .A2(new_n498), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n495), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT101), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n762), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n861), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n749), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n749), .A2(KEYINPUT103), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n871), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n486), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n462), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G142), .B2(new_n484), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n642), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n822), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT104), .ZN(new_n883));
  XOR2_X1   g458(.A(G162), .B(G160), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n651), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n886), .B2(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n873), .A2(new_n881), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(new_n882), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n888), .B(new_n889), .C1(new_n885), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g468(.A(new_n810), .B(G303), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n610), .A2(new_n612), .ZN(new_n895));
  AOI21_X1  g470(.A(G305), .B1(new_n895), .B2(new_n605), .ZN(new_n896));
  OAI211_X1 g471(.A(G305), .B(new_n605), .C1(new_n610), .C2(new_n612), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n894), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G166), .B(new_n810), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n901));
  NAND3_X1  g476(.A1(G290), .A2(new_n600), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n902), .A3(new_n897), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT105), .A3(KEYINPUT106), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT105), .B1(new_n899), .B2(new_n903), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  MUX2_X1   g485(.A(new_n906), .B(new_n910), .S(KEYINPUT42), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n850), .B(new_n637), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n620), .A2(new_n624), .A3(new_n625), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G299), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n632), .A2(new_n624), .A3(new_n625), .A4(new_n620), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n916), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n911), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(G868), .B2(new_n842), .ZN(G295));
  OAI21_X1  g501(.A(new_n925), .B1(G868), .B2(new_n842), .ZN(G331));
  NAND3_X1  g502(.A1(G168), .A2(new_n535), .A3(new_n541), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n534), .A2(new_n508), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n539), .A2(new_n540), .ZN(new_n930));
  OAI21_X1  g505(.A(G286), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n850), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n561), .A2(new_n563), .A3(new_n546), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT98), .B1(new_n935), .B2(new_n842), .ZN(new_n936));
  INV_X1    g511(.A(new_n846), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n849), .B(new_n932), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n917), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n932), .B1(new_n847), .B2(new_n849), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n847), .A2(new_n942), .A3(new_n849), .A4(new_n932), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n939), .B1(new_n944), .B2(new_n920), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n899), .A2(KEYINPUT105), .A3(new_n903), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n908), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT108), .B1(new_n949), .B2(G37), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n947), .B(new_n939), .C1(new_n944), .C2(new_n920), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G37), .B1(new_n945), .B2(new_n948), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n941), .A2(new_n943), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n940), .A2(new_n916), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n934), .A2(new_n938), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n916), .B(KEYINPUT41), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n958), .A2(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n889), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n963), .B2(new_n952), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n958), .A2(new_n959), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n920), .B1(new_n934), .B2(new_n938), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n948), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n889), .A4(new_n951), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n957), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n956), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n957), .B1(new_n950), .B2(new_n955), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n963), .A2(new_n952), .A3(KEYINPUT43), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n971), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n866), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(G40), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(new_n470), .C1(new_n476), .C2(new_n482), .ZN(new_n981));
  NOR2_X1   g556(.A1(G164), .A2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1956), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT57), .B1(new_n630), .B2(new_n631), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n577), .A2(new_n583), .A3(new_n989), .A4(new_n584), .ZN(new_n990));
  INV_X1    g565(.A(new_n495), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n862), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n977), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n866), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT56), .B(G2072), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n995), .A2(new_n981), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n987), .A2(new_n988), .A3(new_n990), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n470), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT69), .B1(new_n474), .B2(new_n475), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n480), .A2(new_n477), .A3(new_n481), .ZN(new_n1002));
  OAI211_X1 g577(.A(G40), .B(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1003), .A2(new_n978), .A3(G2067), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n866), .A2(new_n983), .A3(new_n977), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n981), .B(new_n1005), .C1(new_n983), .C2(new_n982), .ZN(new_n1006));
  INV_X1    g581(.A(G1348), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n913), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n987), .A2(new_n998), .B1(new_n988), .B2(new_n990), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n999), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n995), .A2(new_n981), .A3(new_n996), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1003), .A2(new_n978), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT58), .B(G1341), .ZN(new_n1014));
  OAI22_X1  g589(.A1(new_n1012), .A2(G1996), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n565), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT59), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n565), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1010), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1021), .A2(new_n999), .A3(KEYINPUT61), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT61), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1003), .B1(new_n983), .B2(new_n982), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1956), .B1(new_n1024), .B2(new_n979), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n988), .A2(new_n990), .ZN(new_n1026));
  INV_X1    g601(.A(new_n998), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1023), .B1(new_n1028), .B2(new_n1010), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1020), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n626), .B1(new_n1008), .B2(KEYINPUT60), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT121), .B1(new_n1008), .B2(KEYINPUT60), .ZN(new_n1032));
  OAI211_X1 g607(.A(G160), .B(G40), .C1(new_n982), .C2(new_n983), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1005), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1007), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1004), .ZN(new_n1036));
  AND4_X1   g611(.A1(KEYINPUT121), .A2(new_n1035), .A3(new_n1036), .A4(KEYINPUT60), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n913), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1008), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1011), .B1(new_n1030), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n995), .A2(new_n981), .A3(new_n996), .A4(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(new_n1006), .B2(new_n731), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n866), .B2(new_n977), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1003), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n992), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1049), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1052), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1054), .A2(KEYINPUT53), .A3(new_n1049), .A4(new_n996), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1052), .A2(G301), .A3(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT126), .B(new_n1048), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1063), .B1(new_n1060), .B2(G171), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(KEYINPUT54), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT127), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1052), .A2(new_n1068), .A3(new_n1062), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1052), .B2(new_n1062), .ZN(new_n1070));
  OAI21_X1  g645(.A(G171), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(KEYINPUT54), .C1(G171), .C2(new_n1060), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1047), .A2(new_n1064), .A3(new_n1067), .A4(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT118), .B1(new_n1006), .B2(G2084), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n755), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1033), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(new_n722), .A4(new_n1005), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(G8), .A3(G286), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(KEYINPUT122), .A3(G8), .A4(G286), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1074), .A2(new_n1076), .A3(new_n1079), .A4(G168), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT51), .B1(new_n1085), .B2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1086), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1088), .A2(new_n1091), .B1(new_n1092), .B2(new_n1061), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1061), .A2(KEYINPUT62), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(G303), .A2(G8), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1097), .B(KEYINPUT55), .Z(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1012), .A2(new_n807), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT111), .B(G2090), .Z(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1102), .B1(new_n985), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1024), .A2(KEYINPUT115), .A3(new_n979), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1106), .B2(KEYINPUT116), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1108), .B(new_n1100), .C1(new_n1105), .C2(new_n1104), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1099), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT49), .ZN(new_n1112));
  INV_X1    g687(.A(G1981), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n901), .B2(new_n600), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G305), .A2(G1981), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G8), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n866), .A2(new_n977), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n981), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n901), .A2(new_n1113), .A3(new_n600), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G305), .A2(G1981), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(KEYINPUT49), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1116), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1976), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT52), .B1(G288), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(new_n1119), .C1(new_n1124), .C2(G288), .ZN(new_n1126));
  NOR2_X1   g701(.A1(G288), .A2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n1003), .B2(new_n978), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT52), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1111), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1116), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(KEYINPUT117), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1012), .A2(new_n807), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1102), .B2(new_n1006), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(G8), .A3(new_n1098), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT112), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(KEYINPUT112), .A3(G8), .A4(new_n1098), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1131), .A2(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1096), .A2(new_n1110), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1094), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1141), .A2(new_n1110), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1151), .A2(KEYINPUT63), .A3(new_n1144), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT113), .B1(new_n1123), .B2(new_n1130), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT113), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1132), .A2(new_n1154), .A3(new_n1133), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(G8), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1099), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1156), .A2(KEYINPUT120), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT120), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1148), .A2(new_n1150), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1151), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n810), .A2(new_n1124), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT114), .Z(new_n1166));
  OR2_X1    g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1128), .B1(new_n1167), .B2(new_n1120), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1143), .A2(new_n1162), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n981), .A2(new_n1053), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1172), .A2(G1996), .A3(new_n762), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT110), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n718), .B(new_n720), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(G1996), .B2(new_n762), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n822), .B(new_n824), .Z(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(G290), .B(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1171), .B1(new_n1175), .B2(new_n763), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT46), .B1(new_n1171), .B2(G1996), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1171), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT47), .Z(new_n1187));
  NOR3_X1   g762(.A1(G290), .A2(new_n1171), .A3(G1986), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT48), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1179), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n822), .A2(new_n824), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1177), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n713), .A2(new_n720), .A3(new_n717), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1171), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1182), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g771(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n699), .A2(new_n1198), .ZN(new_n1199));
  OAI211_X1 g773(.A(new_n892), .B(new_n1199), .C1(new_n973), .C2(new_n974), .ZN(G225));
  INV_X1    g774(.A(G225), .ZN(G308));
endmodule


