//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n202), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n216), .B1(new_n209), .B2(new_n208), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT66), .B(G77), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n220), .A2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G87), .A2(G250), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT67), .Z(new_n229));
  AOI211_X1 g0029(.A(new_n218), .B(new_n229), .C1(KEYINPUT1), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G97), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  AOI21_X1  g0045(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G226), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n248), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G232), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n246), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT13), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n259), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(G238), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n256), .A2(new_n257), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n257), .B1(new_n256), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g0069(.A(G169), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT14), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT14), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n272), .B(G169), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n268), .A2(new_n269), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n214), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G68), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n278), .A2(G77), .B1(G20), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G50), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(new_n286), .B1(G1), .B2(G13), .ZN(new_n287));
  NAND4_X1  g0087(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n290), .A2(KEYINPUT11), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n279), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT12), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n214), .A2(G1), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G68), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n284), .A2(KEYINPUT11), .A3(new_n289), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n291), .A2(new_n295), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n274), .B2(G190), .ZN(new_n302));
  OAI21_X1  g0102(.A(G200), .B1(new_n268), .B2(new_n269), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT71), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n307));
  INV_X1    g0107(.A(KEYINPUT16), .ZN(new_n308));
  AND2_X1   g0108(.A1(G58), .A2(G68), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n309), .B2(new_n202), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n282), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(KEYINPUT72), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT7), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n248), .B2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n279), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n308), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n310), .A2(KEYINPUT72), .A3(new_n311), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT72), .B1(new_n310), .B2(new_n311), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n322), .B2(new_n214), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n317), .B(G20), .C1(new_n319), .C2(new_n321), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n332), .A3(new_n289), .ZN(new_n333));
  INV_X1    g0133(.A(G58), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(KEYINPUT8), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT69), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT69), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT8), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G58), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n336), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT70), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT70), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n336), .B(new_n342), .C1(new_n335), .C2(new_n339), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n292), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n341), .A2(new_n343), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n297), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n333), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT75), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n319), .A2(new_n321), .A3(G226), .A4(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT73), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n248), .A2(new_n351), .A3(G226), .A4(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n248), .A2(G223), .A3(new_n249), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n350), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n246), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n265), .A2(new_n254), .B1(new_n260), .B2(new_n259), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(G200), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AOI211_X1 g0159(.A(G190), .B(new_n357), .C1(new_n355), .C2(new_n246), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n348), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n362), .A3(new_n358), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n357), .B1(new_n355), .B2(new_n246), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(KEYINPUT75), .C1(G200), .C2(new_n364), .ZN(new_n365));
  AOI211_X1 g0165(.A(new_n307), .B(new_n347), .C1(new_n361), .C2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n361), .A2(new_n365), .ZN(new_n368));
  INV_X1    g0168(.A(new_n347), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n356), .A2(new_n358), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT74), .B1(new_n371), .B2(G179), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  INV_X1    g0175(.A(G179), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n347), .A2(new_n373), .A3(new_n374), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n375), .B1(new_n364), .B2(new_n376), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n333), .A2(new_n346), .B1(new_n372), .B2(new_n371), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT18), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n366), .A2(new_n370), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n388));
  INV_X1    g0188(.A(G223), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n388), .B1(new_n219), .B2(new_n248), .C1(new_n253), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n246), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n261), .B1(new_n266), .B2(G226), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n372), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(G179), .B2(new_n393), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n287), .A2(new_n288), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n341), .A2(new_n278), .A3(new_n343), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n282), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n297), .A2(G50), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G50), .B2(new_n292), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G200), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n391), .B2(new_n392), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n391), .A2(new_n392), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(G190), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(KEYINPUT9), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n399), .B2(new_n401), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT10), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n407), .A2(new_n408), .A3(new_n413), .A4(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n403), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n297), .A2(G77), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n338), .A2(G58), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n335), .A2(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n418), .A2(new_n283), .B1(new_n214), .B2(new_n219), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n278), .B2(new_n420), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n416), .B1(new_n220), .B2(new_n292), .C1(new_n421), .C2(new_n396), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n423), .B1(new_n424), .B2(new_n248), .C1(new_n250), .C2(new_n254), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n246), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n261), .B1(new_n266), .B2(G244), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n422), .B1(G190), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n376), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n372), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n422), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n387), .A2(new_n415), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n306), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n293), .A2(new_n424), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT84), .B(KEYINPUT25), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n292), .B1(G1), .B2(new_n262), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n289), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(G107), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT79), .A2(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT79), .A2(G116), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT23), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n448), .A2(new_n214), .A3(G107), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT23), .B1(new_n424), .B2(G20), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n447), .A2(new_n277), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n248), .A2(new_n214), .A3(G87), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n248), .A2(new_n454), .A3(new_n214), .A4(G87), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n289), .B1(new_n456), .B2(KEYINPUT24), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n444), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n248), .A2(G250), .A3(new_n249), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n248), .A2(G257), .A3(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G294), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n246), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n258), .B(G45), .C1(new_n263), .C2(KEYINPUT5), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n467), .A2(G264), .A3(new_n264), .ZN(new_n468));
  OR3_X1    g0268(.A1(new_n465), .A2(new_n466), .A3(new_n260), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n372), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(G179), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n459), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n248), .A2(G257), .A3(new_n249), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n248), .A2(G264), .A3(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n322), .A2(G303), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n474), .A2(new_n475), .A3(KEYINPUT81), .A4(new_n476), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n246), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n467), .A2(G270), .A3(new_n264), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n443), .A2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  XOR2_X1   g0287(.A(KEYINPUT79), .B(G116), .Z(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n488), .B2(new_n292), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n447), .A2(new_n293), .A3(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n287), .A2(new_n288), .B1(new_n447), .B2(G20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G283), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n214), .C1(G33), .C2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT83), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n262), .A2(G97), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(KEYINPUT83), .A3(new_n214), .A4(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT20), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT20), .B1(new_n492), .B2(new_n500), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n486), .B(new_n491), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n485), .A2(new_n503), .A3(G169), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n485), .A2(new_n503), .A3(KEYINPUT21), .A4(G169), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n264), .B1(new_n477), .B2(new_n478), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n483), .B1(new_n508), .B2(new_n480), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n509), .A3(G179), .ZN(new_n510));
  AND4_X1   g0310(.A1(new_n473), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n319), .A2(new_n321), .A3(G250), .A4(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n493), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(new_n249), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT77), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(KEYINPUT4), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n264), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n467), .A2(G257), .A3(new_n264), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n469), .ZN(new_n522));
  OAI21_X1  g0322(.A(G169), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(KEYINPUT4), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n524), .A2(new_n493), .A3(new_n519), .A4(new_n512), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n246), .ZN(new_n526));
  INV_X1    g0326(.A(new_n522), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(G179), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n329), .B2(new_n330), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n424), .A2(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n494), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n424), .A2(KEYINPUT6), .A3(G97), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n396), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n292), .A2(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n442), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n396), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(new_n494), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT78), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n282), .A2(G77), .ZN(new_n544));
  INV_X1    g0344(.A(new_n534), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n532), .B2(new_n243), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(new_n214), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n424), .B1(new_n318), .B2(new_n323), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n289), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT78), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n443), .B2(G97), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n523), .A2(new_n528), .B1(new_n543), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n526), .A2(G190), .A3(new_n527), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n549), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n526), .A2(new_n527), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(G200), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n553), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n319), .A2(new_n321), .A3(G238), .A4(new_n249), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(G1698), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n445), .A2(G33), .A3(new_n446), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n246), .ZN(new_n563));
  INV_X1    g0363(.A(G45), .ZN(new_n564));
  OAI21_X1  g0364(.A(G250), .B1(new_n564), .B2(G1), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n258), .A2(G45), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n246), .A2(new_n565), .B1(new_n260), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G200), .ZN(new_n570));
  NAND3_X1  g0370(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n214), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n214), .A2(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT80), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n319), .A2(new_n321), .A3(new_n214), .A4(G68), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n277), .B2(new_n494), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n577), .A2(new_n580), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n420), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n584), .A2(new_n289), .B1(new_n293), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n443), .A2(G87), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n567), .B1(new_n562), .B2(new_n246), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G190), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n570), .A2(new_n586), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(G169), .ZN(new_n591));
  AOI211_X1 g0391(.A(G179), .B(new_n567), .C1(new_n246), .C2(new_n562), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n581), .B(new_n583), .C1(new_n578), .C2(new_n579), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n289), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n585), .A2(new_n293), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n443), .A2(new_n420), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n470), .A2(G200), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n464), .A2(new_n468), .A3(G190), .A4(new_n469), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n590), .B(new_n600), .C1(new_n459), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n491), .B1(new_n541), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n502), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n492), .A2(new_n500), .A3(KEYINPUT20), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n485), .B2(new_n362), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n509), .A2(new_n404), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n437), .A2(new_n511), .A3(new_n558), .A4(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n412), .A2(new_n414), .ZN(new_n615));
  INV_X1    g0415(.A(new_n307), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n368), .A2(new_n369), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n347), .B1(new_n361), .B2(new_n365), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n618), .B2(new_n367), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n435), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n304), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n620), .B1(new_n301), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n378), .A2(new_n379), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n615), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n403), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n437), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n569), .A2(KEYINPUT85), .A3(new_n372), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n588), .B2(G169), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n588), .A2(new_n376), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n632), .A2(new_n599), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n523), .A2(new_n528), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n638), .A2(new_n555), .A3(new_n590), .A4(new_n636), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n543), .A2(new_n552), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n600), .A2(new_n590), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT26), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n636), .A2(new_n590), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n459), .A2(new_n603), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n473), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n558), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n630), .B1(new_n631), .B2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n214), .A2(G13), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n258), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n503), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n612), .B1(new_n656), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n656), .B2(new_n664), .ZN(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n663), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n656), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n473), .A2(new_n663), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n649), .B1(new_n459), .B2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(new_n473), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n674), .ZN(G399));
  INV_X1    g0480(.A(new_n207), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n575), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n211), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n653), .A2(new_n670), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n690), .A2(KEYINPUT87), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n569), .A2(new_n362), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n588), .A2(new_n404), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n596), .A2(new_n597), .A3(new_n587), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n694), .A2(new_n695), .B1(new_n593), .B2(new_n599), .ZN(new_n696));
  AOI211_X1 g0496(.A(KEYINPUT87), .B(KEYINPUT26), .C1(new_n553), .C2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n637), .B1(new_n691), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n652), .B1(new_n699), .B2(KEYINPUT88), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n647), .A2(KEYINPUT26), .A3(new_n638), .A4(new_n555), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT26), .B1(new_n553), .B2(new_n696), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT87), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT88), .B(new_n636), .C1(new_n704), .C2(new_n697), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n670), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n689), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n511), .A2(new_n613), .A3(new_n558), .A4(new_n670), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT31), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n588), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n556), .A2(new_n485), .A3(new_n470), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT86), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n464), .A2(new_n588), .A3(new_n468), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n509), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n715), .B1(new_n717), .B2(new_n528), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n520), .A2(new_n376), .A3(new_n522), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n716), .A3(KEYINPUT30), .A4(new_n509), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n670), .B1(new_n714), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n710), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n721), .A2(new_n712), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n667), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n708), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n687), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n213), .B1(G20), .B2(new_n372), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n376), .A2(new_n404), .A3(KEYINPUT91), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT91), .B1(new_n376), .B2(new_n404), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n214), .A2(G190), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G159), .ZN(new_n740));
  OR3_X1    g0540(.A1(new_n739), .A2(KEYINPUT32), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n735), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n214), .B1(new_n742), .B2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT32), .B1(new_n739), .B2(new_n740), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n214), .A2(new_n362), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n749), .A2(new_n404), .A3(G179), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n322), .B1(new_n750), .B2(G87), .ZN(new_n751));
  XOR2_X1   g0551(.A(new_n751), .B(KEYINPUT92), .Z(new_n752));
  NOR2_X1   g0552(.A1(new_n376), .A2(new_n404), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n736), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n376), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n736), .A2(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n279), .B1(new_n756), .B2(new_n219), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n748), .A2(new_n755), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G58), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT90), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n748), .A2(new_n753), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n748), .B2(new_n753), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n752), .B(new_n760), .C1(new_n281), .C2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n737), .A2(G179), .A3(new_n404), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT94), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n747), .B(new_n765), .C1(G107), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n754), .ZN(new_n773));
  NOR2_X1   g0573(.A1(KEYINPUT33), .A2(G317), .ZN(new_n774));
  AND2_X1   g0574(.A1(KEYINPUT33), .A2(G317), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n758), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G303), .B2(new_n750), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n744), .A2(G294), .ZN(new_n780));
  INV_X1    g0580(.A(new_n756), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n248), .B1(new_n781), .B2(G311), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G326), .B1(new_n738), .B2(G329), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n771), .B2(G283), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n732), .B1(new_n772), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n258), .B1(new_n657), .B2(G45), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n682), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n241), .A2(G45), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n681), .A2(new_n248), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n792), .B(new_n793), .C1(G45), .C2(new_n211), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n248), .A2(new_n207), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n605), .B2(new_n681), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n732), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n791), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n787), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n666), .B2(new_n801), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n668), .A2(new_n790), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n666), .A2(new_n667), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  NOR2_X1   g0609(.A1(new_n435), .A2(new_n663), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n430), .A2(new_n431), .B1(new_n422), .B2(new_n663), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n621), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n688), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n663), .B1(new_n646), .B2(new_n652), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n790), .B1(new_n818), .B2(new_n728), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n814), .A2(new_n727), .A3(new_n817), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G77), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n732), .A2(new_n799), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n791), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n816), .A2(new_n800), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n770), .A2(new_n279), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G143), .A2(new_n759), .B1(new_n781), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n754), .C1(new_n764), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n827), .B1(KEYINPUT34), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n750), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n248), .B1(new_n834), .B2(new_n281), .C1(new_n739), .C2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G58), .B2(new_n744), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n833), .B(new_n837), .C1(KEYINPUT34), .C2(new_n832), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n771), .A2(G87), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n322), .B1(new_n754), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n834), .A2(new_n424), .B1(new_n447), .B2(new_n756), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(G294), .C2(new_n759), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n783), .A2(G303), .B1(new_n738), .B2(G311), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n839), .A2(new_n745), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n838), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT95), .ZN(new_n847));
  INV_X1    g0647(.A(new_n732), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n846), .B2(KEYINPUT95), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n825), .B(new_n826), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n821), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  OAI211_X1 g0652(.A(G116), .B(new_n215), .C1(new_n535), .C2(KEYINPUT35), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(KEYINPUT35), .B2(new_n535), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT36), .ZN(new_n855));
  OR3_X1    g0655(.A1(new_n211), .A2(new_n219), .A3(new_n309), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n201), .A2(G68), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n258), .B(G13), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n722), .B1(new_n709), .B2(KEYINPUT31), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT31), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n861), .B(new_n670), .C1(new_n714), .C2(new_n721), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n437), .B(G330), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n300), .A2(new_n663), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n301), .A2(new_n304), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n276), .A2(new_n300), .A3(new_n663), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n816), .ZN(new_n869));
  INV_X1    g0669(.A(new_n862), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n869), .B1(new_n724), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n661), .B1(new_n333), .B2(new_n346), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n386), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n661), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n347), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n378), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n872), .B2(KEYINPUT96), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n877), .A3(new_n618), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n383), .B2(new_n384), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n368), .A2(new_n369), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT96), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n875), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n880), .B1(new_n882), .B2(KEYINPUT37), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n873), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n875), .B1(new_n619), .B2(new_n626), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n876), .B2(new_n618), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n886), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n871), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n877), .B1(new_n876), .B2(new_n618), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n886), .B1(new_n887), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT40), .B1(new_n885), .B2(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n894), .A2(KEYINPUT40), .B1(new_n871), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n863), .B1(new_n900), .B2(new_n667), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n437), .B1(new_n860), .B2(new_n862), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n630), .B1(new_n708), .B2(new_n631), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n903), .B(new_n904), .Z(new_n905));
  AOI21_X1  g0705(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n906));
  INV_X1    g0706(.A(new_n868), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n885), .A2(new_n898), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n908), .A2(new_n909), .B1(new_n627), .B2(new_n661), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n301), .A2(new_n663), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n885), .A2(new_n892), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n885), .B2(new_n898), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT97), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT97), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n893), .B2(KEYINPUT39), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n258), .B2(new_n657), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n905), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n859), .B1(new_n923), .B2(new_n924), .ZN(G367));
  NOR2_X1   g0725(.A1(new_n695), .A2(new_n670), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n636), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n647), .B2(new_n926), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT98), .Z(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n668), .A2(new_n678), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n555), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n558), .B1(new_n934), .B2(new_n670), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT99), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n638), .A2(new_n555), .A3(new_n663), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT100), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(KEYINPUT100), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n943), .A3(new_n929), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n938), .A2(new_n656), .A3(new_n670), .A4(new_n678), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n553), .B1(new_n938), .B2(new_n676), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n946), .B(new_n947), .C1(new_n663), .C2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n940), .B(new_n941), .C1(KEYINPUT43), .C2(new_n930), .ZN(new_n950));
  AND4_X1   g0750(.A1(new_n931), .A2(new_n944), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n944), .A2(new_n950), .B1(new_n949), .B2(new_n931), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n938), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n674), .B1(new_n677), .B2(new_n671), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT44), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT44), .ZN(new_n957));
  INV_X1    g0757(.A(new_n955), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n938), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n954), .A2(new_n960), .A3(new_n955), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT45), .B1(new_n938), .B2(new_n958), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n932), .B1(new_n956), .B2(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n672), .B(new_n677), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n729), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n682), .B(KEYINPUT41), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n788), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n929), .A2(new_n801), .ZN(new_n969));
  INV_X1    g0769(.A(new_n793), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n237), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n802), .B1(new_n207), .B2(new_n585), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n790), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n769), .A2(new_n494), .B1(new_n974), .B2(new_n739), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G311), .B2(new_n783), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n750), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  INV_X1    g0777(.A(G303), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n977), .B1(new_n840), .B2(new_n756), .C1(new_n978), .C2(new_n758), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT46), .B1(new_n750), .B2(new_n488), .ZN(new_n980));
  INV_X1    g0780(.A(G294), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n322), .B1(new_n754), .B2(new_n981), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n976), .B(new_n983), .C1(new_n424), .C2(new_n743), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n744), .A2(G68), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n829), .B2(new_n758), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT101), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(KEYINPUT101), .ZN(new_n988));
  INV_X1    g0788(.A(new_n201), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n781), .A2(new_n989), .B1(new_n773), .B2(G159), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n248), .C1(new_n334), .C2(new_n834), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G137), .B2(new_n738), .ZN(new_n992));
  INV_X1    g0792(.A(new_n769), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(new_n220), .B1(G143), .B2(new_n783), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n984), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT47), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n848), .B1(new_n996), .B2(new_n997), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n973), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n953), .A2(new_n968), .B1(new_n969), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1001), .A2(KEYINPUT102), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(KEYINPUT102), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(new_n1003), .ZN(G387));
  AOI21_X1  g0804(.A(new_n683), .B1(new_n730), .B2(new_n964), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n730), .B2(new_n964), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n684), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n564), .B1(new_n279), .B2(new_n822), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n418), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n281), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1007), .B(new_n1008), .C1(new_n1010), .C2(KEYINPUT50), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT50), .B2(new_n1010), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n793), .C1(new_n564), .C2(new_n234), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n796), .A2(new_n1007), .B1(new_n424), .B2(new_n681), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT103), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n802), .B1(new_n1015), .B2(KEYINPUT103), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n790), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n744), .A2(G283), .B1(G294), .B2(new_n750), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n783), .A2(G322), .B1(G311), .B2(new_n773), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n758), .A2(new_n974), .B1(new_n756), .B2(new_n978), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT106), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT107), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n322), .B1(new_n769), .B2(new_n447), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G326), .B2(new_n738), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n248), .B1(new_n834), .B2(new_n219), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT104), .B(G150), .Z(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n738), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n770), .B2(new_n494), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(KEYINPUT105), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT105), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n744), .A2(new_n420), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G50), .A2(new_n759), .B1(new_n781), .B2(G68), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n740), .C2(new_n764), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n345), .B2(new_n773), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1030), .A2(new_n1033), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1018), .B1(new_n1045), .B2(new_n732), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1046), .A2(KEYINPUT109), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1046), .A2(KEYINPUT109), .B1(new_n677), .B2(new_n801), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n789), .A2(new_n964), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT110), .B1(new_n1006), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1006), .A2(KEYINPUT110), .A3(new_n1049), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(G393));
  OAI22_X1  g0853(.A1(new_n961), .A2(new_n962), .B1(new_n956), .B2(new_n959), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n933), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n963), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n788), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n954), .A2(new_n801), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n750), .A2(G68), .B1(new_n1009), .B2(new_n781), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n738), .A2(G143), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n322), .B1(new_n989), .B2(new_n773), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G77), .B2(new_n744), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n764), .A2(new_n829), .B1(new_n740), .B2(new_n758), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT51), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n839), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n783), .A2(G317), .B1(G311), .B2(new_n759), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  AOI21_X1  g0870(.A(new_n248), .B1(new_n750), .B2(G283), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G303), .A2(new_n773), .B1(new_n781), .B2(G294), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n739), .C2(new_n777), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n488), .B2(new_n744), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1070), .B(new_n1074), .C1(new_n424), .C2(new_n770), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n848), .B1(new_n1068), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n244), .A2(new_n970), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n802), .B1(new_n494), .B2(new_n207), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n790), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR4_X1   g0879(.A1(new_n1059), .A2(new_n1060), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1057), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n730), .A2(new_n964), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1056), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n963), .A2(new_n730), .A3(new_n964), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n682), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1085), .ZN(G390));
  XOR2_X1   g0886(.A(new_n912), .B(KEYINPUT112), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n893), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n652), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n636), .B1(new_n704), .B2(new_n697), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT88), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n663), .B1(new_n1093), .B2(new_n705), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n812), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n435), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n810), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1089), .B1(new_n1097), .B2(new_n907), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n913), .B1(new_n906), .B2(new_n907), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n917), .A2(new_n919), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n813), .B1(new_n866), .B2(new_n867), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n727), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(KEYINPUT113), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT113), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1098), .A2(new_n1100), .A3(new_n1105), .A4(new_n1102), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1101), .B(G330), .C1(new_n860), .C2(new_n862), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n917), .A2(new_n919), .A3(new_n1099), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n670), .B(new_n1096), .C1(new_n700), .C2(new_n706), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n811), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1088), .B1(new_n1111), .B2(new_n868), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1108), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1104), .A2(new_n789), .A3(new_n1106), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n917), .A2(new_n799), .A3(new_n919), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n823), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n790), .B1(new_n345), .B2(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n424), .A2(new_n754), .B1(new_n758), .B2(new_n605), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n322), .B1(new_n834), .B2(new_n574), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(G97), .C2(new_n781), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n783), .A2(G283), .B1(new_n738), .B2(G294), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n822), .C2(new_n743), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n750), .A2(new_n1035), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT53), .Z(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1124), .B1(new_n1125), .B2(new_n739), .C1(new_n1126), .C2(new_n764), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n835), .A2(new_n758), .B1(new_n754), .B2(new_n830), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT54), .B(G143), .Z(new_n1129));
  AOI211_X1 g0929(.A(new_n322), .B(new_n1128), .C1(new_n781), .C2(new_n1129), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1130), .B1(new_n740), .B2(new_n743), .C1(new_n201), .C2(new_n769), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1122), .A2(new_n827), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1117), .B1(new_n1132), .B2(new_n732), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1115), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1114), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1107), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(KEYINPUT113), .B2(new_n1103), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n630), .B(new_n863), .C1(new_n708), .C2(new_n631), .ZN(new_n1138));
  OAI211_X1 g0938(.A(G330), .B(new_n816), .C1(new_n860), .C2(new_n862), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n727), .A2(new_n1101), .B1(new_n1139), .B2(new_n907), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n726), .ZN(new_n1141));
  OAI211_X1 g0941(.A(G330), .B(new_n816), .C1(new_n860), .C2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n907), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1107), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n906), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1097), .A2(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT114), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT114), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1137), .A2(new_n1106), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1104), .A2(new_n1106), .A3(new_n1113), .A4(new_n1147), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n682), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1135), .B1(new_n1151), .B2(new_n1153), .ZN(G378));
  NOR2_X1   g0954(.A1(new_n248), .A2(G41), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G50), .B(new_n1155), .C1(new_n262), .C2(new_n263), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n494), .A2(new_n754), .B1(new_n758), .B2(new_n424), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1155), .B1(new_n834), .B2(new_n219), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1157), .B(new_n1158), .C1(new_n420), .C2(new_n781), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n783), .A2(G116), .B1(new_n738), .B2(G283), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n993), .A2(G58), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n985), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n758), .A2(new_n1126), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n754), .A2(new_n835), .B1(new_n756), .B2(new_n830), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n750), .C2(new_n1129), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n764), .B2(new_n1125), .C1(new_n743), .C2(new_n829), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n262), .B(new_n263), .C1(new_n769), .C2(new_n740), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G124), .B2(new_n738), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1174), .A2(new_n732), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n790), .B1(new_n989), .B2(new_n1116), .C1(new_n1175), .C2(KEYINPUT115), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n615), .A2(new_n629), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n402), .A2(new_n661), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1178), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n415), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT116), .B(KEYINPUT117), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1179), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n415), .A2(new_n1180), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n403), .B(new_n1178), .C1(new_n412), .C2(new_n414), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1184), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n800), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1176), .B(new_n1191), .C1(KEYINPUT115), .C2(new_n1175), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT118), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n900), .A2(new_n1194), .A3(new_n667), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1190), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1184), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1196), .A2(KEYINPUT118), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n871), .A2(new_n899), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1101), .B1(new_n860), .B2(new_n862), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n885), .B2(new_n892), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT40), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1199), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1198), .B1(new_n1203), .B2(G330), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1195), .A2(new_n1204), .B1(new_n920), .B2(new_n911), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1194), .B1(new_n900), .B2(new_n667), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n920), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(G330), .A3(new_n1198), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n910), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1192), .B1(new_n1210), .B2(new_n789), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1138), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1152), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n682), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1152), .A2(new_n1212), .B1(new_n1209), .B2(new_n1205), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1216), .A2(KEYINPUT57), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1211), .B1(new_n1215), .B2(new_n1217), .ZN(G375));
  XOR2_X1   g1018(.A(new_n966), .B(KEYINPUT119), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n790), .B1(new_n1116), .B2(G68), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n248), .B1(new_n773), .B2(new_n488), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n424), .B2(new_n756), .C1(new_n834), .C2(new_n494), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G294), .B2(new_n783), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n978), .B2(new_n739), .C1(new_n770), .C2(new_n822), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1040), .B1(new_n840), .B2(new_n758), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT120), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G137), .A2(new_n759), .B1(new_n773), .B2(new_n1129), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n829), .B2(new_n756), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n322), .B(new_n1231), .C1(G159), .C2(new_n750), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n281), .B2(new_n743), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1161), .B1(new_n1126), .B2(new_n739), .C1(new_n835), .C2(new_n764), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n1227), .A2(new_n1229), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1223), .B1(new_n1235), .B2(new_n732), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n868), .B2(new_n800), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(new_n1146), .B2(new_n788), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1222), .A2(new_n1238), .ZN(G381));
  NAND3_X1  g1039(.A1(new_n1051), .A2(new_n808), .A3(new_n1052), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G384), .A2(G381), .A3(new_n1240), .A4(G390), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n683), .B1(new_n1216), .B2(KEYINPUT57), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1213), .A2(new_n1210), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G378), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1211), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1241), .A2(G387), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(G407));
  OAI211_X1 g1050(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  INV_X1    g1051(.A(KEYINPUT125), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G375), .A2(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n662), .A2(G213), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1135), .B(new_n1211), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1219), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1213), .A2(new_n1210), .A3(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1258), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n682), .C1(new_n1221), .C2(KEYINPUT60), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1220), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1221), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1261), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n851), .B1(new_n1266), .B2(new_n1238), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1264), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1269), .A2(new_n1147), .A3(new_n683), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1238), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(G384), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1267), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT123), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1254), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(G378), .B2(G375), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1274), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT63), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(G390), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1052), .ZN(new_n1284));
  OAI21_X1  g1084(.A(G396), .B1(new_n1284), .B2(new_n1050), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1285), .A2(new_n1240), .B1(new_n1001), .B2(G390), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1001), .B(G390), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1285), .A2(new_n1240), .A3(KEYINPUT124), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT124), .B1(new_n1285), .B2(new_n1240), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1288), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1267), .A2(new_n1273), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n851), .B(new_n1238), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1247), .B1(new_n1246), .B2(new_n1211), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1295), .B(new_n1299), .C1(new_n1300), .C2(new_n1276), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1301), .A4(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1252), .B1(new_n1281), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1292), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1299), .A2(new_n1295), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1302), .B1(new_n1277), .B2(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1278), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1310));
  NOR4_X1   g1110(.A1(new_n1300), .A2(KEYINPUT123), .A3(new_n1276), .A4(new_n1274), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1308), .A2(KEYINPUT125), .A3(new_n1312), .A4(new_n1293), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1304), .A2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1307), .B(KEYINPUT126), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1259), .A2(new_n1316), .A3(new_n1274), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1316), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(KEYINPUT127), .B(new_n1316), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1315), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1322), .B2(new_n1292), .ZN(G405));
  NAND2_X1  g1123(.A1(new_n1253), .A2(new_n1248), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1324), .B(new_n1274), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1325), .B(new_n1305), .ZN(G402));
endmodule


