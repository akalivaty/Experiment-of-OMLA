//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n552, new_n553,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT68), .Z(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n461), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n466), .B(KEYINPUT69), .ZN(G160));
  NAND2_X1  g042(.A1(new_n461), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G124), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n470), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND4_X1  g056(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n458), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT71), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n461), .A2(new_n484), .A3(G138), .A4(new_n458), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n472), .A2(new_n474), .A3(G126), .A4(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n461), .A2(KEYINPUT70), .A3(G126), .A4(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n482), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n458), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n486), .A2(new_n491), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n496), .B1(new_n489), .B2(new_n490), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n500), .A2(new_n486), .A3(new_n501), .A4(new_n493), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n504), .A2(KEYINPUT6), .A3(G651), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT6), .B1(new_n504), .B2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(G62), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n511), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NOR2_X1   g098(.A1(new_n507), .A2(new_n512), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT74), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n505), .A2(new_n506), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n528), .B(new_n530), .C1(new_n516), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n516), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n524), .A2(G52), .B1(G651), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n507), .A2(new_n516), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n516), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n524), .A2(G43), .B1(G651), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n539), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g126(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n552));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(G188));
  NAND2_X1  g131(.A1(new_n531), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT77), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n524), .A2(new_n560), .A3(G53), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  OAI211_X1 g138(.A(KEYINPUT77), .B(new_n563), .C1(new_n557), .C2(new_n558), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n516), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n539), .A2(G91), .B1(G651), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n524), .A2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n539), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n516), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(G48), .A2(new_n524), .B1(new_n539), .B2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n539), .A2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n524), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G651), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(G290));
  AOI22_X1  g163(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n524), .A2(G54), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n539), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT79), .B1(new_n596), .B2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  MUX2_X1   g173(.A(KEYINPUT79), .B(new_n597), .S(new_n598), .Z(G284));
  MUX2_X1   g174(.A(KEYINPUT79), .B(new_n597), .S(new_n598), .Z(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n570), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n570), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n596), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n596), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n476), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n469), .A2(G123), .B1(new_n476), .B2(G135), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n458), .A2(G111), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT81), .Z(new_n617));
  OAI21_X1  g192(.A(new_n614), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2438), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G14), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT17), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT18), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n639), .B2(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2096), .B(G2100), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G227));
  XNOR2_X1  g225(.A(G1971), .B(G1976), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT85), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XOR2_X1   g228(.A(G1956), .B(G2474), .Z(new_n654));
  XOR2_X1   g229(.A(G1961), .B(G1966), .Z(new_n655));
  AND2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT20), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n653), .A2(new_n656), .A3(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G1986), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G1981), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  NOR2_X1   g243(.A1(G16), .A2(G24), .ZN(new_n669));
  XOR2_X1   g244(.A(G290), .B(KEYINPUT87), .Z(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(G16), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(G1986), .Z(new_n672));
  OAI21_X1  g247(.A(G2104), .B1(new_n458), .B2(G107), .ZN(new_n673));
  INV_X1    g248(.A(G95), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n673), .B1(new_n674), .B2(new_n458), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G131), .B2(new_n476), .ZN(new_n677));
  INV_X1    g252(.A(G119), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n468), .ZN(new_n679));
  MUX2_X1   g254(.A(G25), .B(new_n679), .S(G29), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT35), .B(G1991), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n511), .B2(new_n521), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(G22), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n685), .A2(KEYINPUT90), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT90), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n684), .A2(G23), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n684), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT89), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n687), .A2(G1971), .A3(new_n688), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n691), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n684), .A2(G6), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G305), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT32), .B(G1981), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT88), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(KEYINPUT34), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n691), .A2(new_n697), .A3(new_n698), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n708));
  NOR3_X1   g283(.A1(new_n707), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n672), .B(new_n683), .C1(new_n706), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT36), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n699), .A2(KEYINPUT34), .A3(new_n705), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n708), .B1(new_n707), .B2(new_n704), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n714), .A2(new_n715), .A3(new_n672), .A4(new_n683), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G32), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT98), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT26), .ZN(new_n722));
  NAND2_X1  g297(.A1(G105), .A2(G2104), .ZN(new_n723));
  INV_X1    g298(.A(G141), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n475), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g300(.A1(G129), .A2(new_n469), .B1(new_n725), .B2(new_n458), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(new_n718), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT99), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n729), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G2072), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n718), .A2(G33), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT94), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G2105), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT92), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n476), .A2(G139), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n743), .A2(KEYINPUT25), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n737), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n746), .B(KEYINPUT93), .ZN(new_n752));
  AOI21_X1  g327(.A(KEYINPUT95), .B1(new_n752), .B2(new_n737), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n733), .B(new_n734), .C1(new_n754), .C2(new_n718), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n749), .A2(new_n750), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(KEYINPUT95), .A3(new_n737), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n718), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n734), .ZN(new_n759));
  OAI21_X1  g334(.A(G2072), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(KEYINPUT30), .A2(G28), .ZN(new_n761));
  NOR2_X1   g336(.A1(KEYINPUT30), .A2(G28), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n761), .A2(new_n762), .A3(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n618), .B2(G29), .ZN(new_n764));
  NAND2_X1  g339(.A1(G160), .A2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(G34), .Z(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(G29), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n732), .A2(new_n755), .A3(new_n760), .A4(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT102), .ZN(new_n772));
  INV_X1    g347(.A(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G29), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n718), .A2(KEYINPUT102), .A3(G27), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G164), .C2(new_n718), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  OR2_X1    g352(.A1(G16), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G286), .B2(new_n684), .ZN(new_n779));
  INV_X1    g354(.A(G1966), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n684), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n684), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1961), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT100), .B(KEYINPUT31), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G11), .Z(new_n787));
  NOR4_X1   g362(.A1(new_n777), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n771), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT103), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n779), .A2(new_n780), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n768), .A2(new_n769), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n718), .A2(G26), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n476), .A2(G140), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT91), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n469), .A2(G128), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n795), .B(new_n802), .S(KEYINPUT28), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n806));
  INV_X1    g381(.A(G20), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G16), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n808), .C1(new_n570), .C2(new_n684), .ZN(new_n809));
  INV_X1    g384(.A(G1956), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1341), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n549), .A2(G16), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G16), .B2(G19), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n804), .B(new_n811), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n771), .A2(new_n788), .A3(new_n793), .A4(new_n791), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(KEYINPUT103), .ZN(new_n817));
  AND3_X1   g392(.A1(new_n717), .A2(new_n794), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(G29), .A2(G35), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G162), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT29), .B(G2090), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n684), .A2(G4), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n596), .B2(new_n684), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1348), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n814), .A2(new_n812), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n818), .A2(new_n822), .A3(new_n825), .A4(new_n826), .ZN(G150));
  INV_X1    g402(.A(KEYINPUT104), .ZN(new_n828));
  NAND2_X1  g403(.A1(G150), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g404(.A1(new_n826), .A2(new_n717), .A3(new_n794), .A4(new_n817), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n830), .A2(KEYINPUT104), .A3(new_n822), .A4(new_n825), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n539), .A2(G93), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n524), .A2(G55), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n833), .B(new_n834), .C1(new_n586), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  XOR2_X1   g413(.A(new_n836), .B(new_n548), .Z(new_n839));
  XOR2_X1   g414(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n604), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n841), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n838), .B1(new_n844), .B2(G860), .ZN(G145));
  INV_X1    g420(.A(new_n801), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n754), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n480), .B(KEYINPUT105), .ZN(new_n848));
  XNOR2_X1  g423(.A(G160), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n618), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n679), .B(new_n727), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n469), .A2(G130), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n476), .A2(G142), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT106), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(KEYINPUT106), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n855), .A2(new_n857), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n851), .A2(new_n862), .A3(new_n852), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n611), .B(new_n498), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n867), .A3(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(G303), .B(G288), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(G290), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(G290), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G305), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n875), .A2(new_n582), .A3(new_n581), .A4(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n881));
  AND2_X1   g456(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n839), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n606), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n596), .A2(new_n887), .A3(new_n570), .ZN(new_n888));
  OAI21_X1  g463(.A(KEYINPUT107), .B1(new_n562), .B2(new_n569), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n559), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n890), .A2(new_n887), .A3(new_n564), .A4(new_n568), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n842), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n888), .A2(new_n892), .A3(KEYINPUT41), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n894), .B1(new_n898), .B2(new_n886), .ZN(new_n899));
  OR3_X1    g474(.A1(new_n883), .A2(new_n884), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n883), .B2(new_n884), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(G868), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G868), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT109), .B1(new_n836), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n906), .B2(new_n902), .ZN(G295));
  AOI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n902), .ZN(G331));
  INV_X1    g483(.A(KEYINPUT112), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT111), .ZN(new_n910));
  NAND3_X1  g485(.A1(G168), .A2(KEYINPUT110), .A3(G171), .ZN(new_n911));
  NAND2_X1  g486(.A1(G171), .A2(KEYINPUT110), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(G286), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n839), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n839), .B1(new_n911), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n893), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n839), .A2(new_n911), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT111), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n896), .B(new_n897), .C1(new_n917), .C2(new_n916), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n909), .B(new_n871), .C1(new_n924), .C2(new_n880), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n880), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT112), .B1(new_n926), .B2(G37), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n923), .A3(new_n880), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n893), .A2(new_n916), .A3(new_n917), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n918), .A2(new_n921), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n898), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n871), .B(new_n929), .C1(new_n933), .C2(new_n880), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(KEYINPUT44), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n925), .A2(new_n927), .A3(KEYINPUT43), .A4(new_n929), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n928), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(KEYINPUT113), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(KEYINPUT113), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(G397));
  XNOR2_X1  g518(.A(KEYINPUT114), .B(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n498), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G40), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n463), .A2(new_n465), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n679), .B(new_n682), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT117), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n801), .B(G2067), .Z(new_n954));
  NAND2_X1  g529(.A1(new_n727), .A2(G1996), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT115), .B1(G290), .B2(G1986), .ZN(new_n960));
  OR3_X1    g535(.A1(G290), .A2(KEYINPUT115), .A3(G1986), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n951), .A2(G1986), .A3(G290), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT116), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n959), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(G303), .A2(G8), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT55), .Z(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n499), .A2(new_n969), .A3(new_n502), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n946), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n944), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n972), .A2(new_n949), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT118), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(KEYINPUT118), .A3(new_n973), .ZN(new_n977));
  AOI21_X1  g552(.A(G1971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n498), .A2(new_n969), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n950), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G2090), .ZN(new_n985));
  OAI211_X1 g560(.A(G8), .B(new_n968), .C1(new_n978), .C2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT119), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n971), .A2(KEYINPUT118), .A3(new_n973), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT118), .B1(new_n971), .B2(new_n973), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n690), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n985), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(new_n968), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n950), .B1(KEYINPUT50), .B2(new_n980), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n499), .A2(new_n982), .A3(new_n969), .A4(new_n502), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G2090), .ZN(new_n1000));
  OAI21_X1  g575(.A(G8), .B1(new_n978), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n968), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G305), .B(G1981), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n950), .A2(new_n980), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n988), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1011), .B2(G288), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n693), .A2(G1976), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n1012), .A2(KEYINPUT52), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n1012), .B2(KEYINPUT52), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n1012), .A2(new_n1015), .A3(KEYINPUT52), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1010), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n980), .A2(new_n946), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n949), .B(new_n1020), .C1(new_n970), .C2(new_n946), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n780), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n979), .A2(new_n983), .A3(new_n769), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n988), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(G168), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n996), .A2(new_n1003), .A3(new_n1019), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1018), .B1(new_n987), .B2(new_n995), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n993), .A2(new_n968), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1029), .A2(KEYINPUT63), .A3(new_n1025), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n976), .A2(new_n1033), .A3(new_n977), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1961), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n984), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n465), .A2(KEYINPUT123), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1039), .A2(new_n948), .A3(new_n463), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1035), .B(G2078), .C1(new_n465), .C2(KEYINPUT123), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n947), .A2(new_n972), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1036), .A2(G301), .A3(new_n1038), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT124), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1034), .A2(new_n1035), .B1(new_n1037), .B2(new_n984), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT124), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(G301), .A4(new_n1042), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n1021), .A2(new_n1035), .A3(G2078), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n989), .A2(new_n990), .A3(G2078), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1038), .B(new_n1049), .C1(new_n1050), .C2(KEYINPUT53), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(G301), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1046), .A2(G171), .A3(new_n1042), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT54), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n986), .A2(KEYINPUT119), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n994), .B1(new_n993), .B2(new_n968), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1003), .B(new_n1019), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1022), .A2(G168), .A3(new_n1023), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n988), .A2(KEYINPUT122), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(KEYINPUT51), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT51), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1024), .A2(G286), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n570), .A2(KEYINPUT57), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n562), .B2(new_n569), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n971), .A2(new_n973), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1956), .B1(new_n997), .B2(new_n998), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n971), .A2(new_n973), .A3(new_n1074), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n979), .B2(new_n983), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n950), .A2(new_n980), .A3(G2067), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n842), .A2(KEYINPUT60), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1082), .A2(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT58), .B(G1341), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n974), .A2(G1996), .B1(new_n1008), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n549), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n549), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1086), .A2(new_n842), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1084), .A2(new_n596), .A3(new_n1085), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1077), .A2(new_n1081), .A3(KEYINPUT61), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1088), .A2(new_n1096), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1081), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1102), .A2(new_n1077), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1069), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1057), .A2(new_n1061), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n996), .A2(new_n1018), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1010), .A2(new_n1011), .A3(new_n693), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G1981), .B2(G305), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1009), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1032), .A2(new_n1105), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n1067), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1112));
  AOI21_X1  g687(.A(G301), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n1060), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n1003), .A4(new_n1029), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n966), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n954), .A2(new_n728), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT46), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1122), .A2(new_n951), .B1(KEYINPUT126), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n951), .A2(new_n956), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(KEYINPUT126), .B2(new_n1123), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1125), .A2(KEYINPUT126), .A3(new_n1123), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT47), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n962), .B(KEYINPUT48), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n959), .A2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n679), .A2(new_n681), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n958), .A2(new_n1132), .B1(G2067), .B2(new_n801), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n951), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT127), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g712(.A1(new_n937), .A2(new_n649), .A3(new_n939), .ZN(new_n1139));
  NOR2_X1   g713(.A1(G401), .A2(G229), .ZN(new_n1140));
  NAND4_X1  g714(.A1(new_n1139), .A2(new_n1140), .A3(new_n872), .A4(G319), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


