//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930;
  OR2_X1    g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT0), .A2(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  MUX2_X1   g004(.A(new_n189), .B(new_n188), .S(new_n190), .Z(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n192), .A2(new_n193), .A3(G137), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G134), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(G137), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n196), .A2(new_n197), .A3(G137), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n195), .B(new_n198), .C1(new_n199), .C2(KEYINPUT11), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT64), .A2(G134), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT64), .A2(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n194), .B1(new_n206), .B2(new_n192), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n202), .B1(new_n207), .B2(new_n198), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n191), .B1(new_n201), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n202), .A3(new_n198), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n204), .A2(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n199), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n215), .B1(new_n218), .B2(KEYINPUT66), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n220), .A3(KEYINPUT1), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n190), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n190), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .A3(new_n215), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n212), .B(new_n214), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n200), .A2(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n212), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT65), .A3(new_n191), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n209), .A2(KEYINPUT30), .A3(new_n225), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT2), .B(G113), .Z(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n231), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n240));
  NOR2_X1   g054(.A1(G237), .A2(G953), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G210), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n240), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G101), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n209), .A2(new_n237), .A3(new_n225), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT31), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT69), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n239), .A2(new_n245), .A3(new_n246), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n229), .A2(new_n238), .ZN(new_n253));
  INV_X1    g067(.A(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n245), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n247), .A2(new_n262), .A3(KEYINPUT31), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n249), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G472), .ZN(new_n265));
  INV_X1    g079(.A(G902), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT32), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n232), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n229), .B2(new_n230), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n254), .B1(new_n271), .B2(new_n238), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n245), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n258), .A2(new_n259), .ZN(new_n274));
  OR3_X1    g088(.A1(new_n273), .A2(KEYINPUT29), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n209), .ZN(new_n276));
  INV_X1    g090(.A(new_n225), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n238), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT71), .A3(new_n246), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n238), .C1(new_n276), .C2(new_n277), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT28), .A3(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT29), .A3(new_n245), .A4(new_n257), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n275), .A2(new_n266), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G472), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n264), .A2(KEYINPUT32), .A3(new_n265), .A4(new_n266), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n269), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G217), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(new_n266), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G119), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n215), .A2(G119), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n295), .B1(new_n298), .B2(new_n294), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n294), .A2(new_n296), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT24), .B(G110), .Z(new_n301));
  OAI22_X1  g115(.A1(new_n299), .A2(G110), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(G125), .B(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(G125), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n305), .A2(KEYINPUT16), .A3(G140), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(G146), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n216), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n216), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT74), .A3(new_n307), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n304), .A2(new_n313), .A3(G146), .A4(new_n306), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n300), .A2(new_n301), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n299), .A2(G110), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT73), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n309), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT22), .B(G137), .Z(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n326), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n329), .B2(new_n324), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n266), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n266), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n292), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n291), .A2(G902), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n289), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n341));
  OAI21_X1  g155(.A(G214), .B1(G237), .B2(G902), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n342), .B(KEYINPUT81), .Z(new_n343));
  AND2_X1   g157(.A1(new_n321), .A2(G952), .ZN(new_n344));
  NAND2_X1  g158(.A1(G234), .A2(G237), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n346), .B(KEYINPUT92), .Z(new_n347));
  AND3_X1   g161(.A1(new_n345), .A2(G902), .A3(G953), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT21), .B(G898), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G210), .B1(G237), .B2(G902), .ZN(new_n353));
  INV_X1    g167(.A(G104), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G107), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(G107), .ZN(new_n357));
  OAI21_X1  g171(.A(G101), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  INV_X1    g173(.A(G107), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g176(.A(G101), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n359), .A2(new_n364), .A3(new_n360), .A4(G104), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n355), .A4(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n358), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G113), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n293), .A2(G116), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n375), .A2(new_n376), .B1(new_n236), .B2(new_n233), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT79), .B(new_n358), .C1(new_n367), .C2(new_n368), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n362), .A2(new_n355), .A3(new_n365), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT4), .B(new_n381), .C1(new_n367), .C2(new_n368), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n238), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT82), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(G110), .B(G122), .Z(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n388), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n391), .A3(new_n384), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT6), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(KEYINPUT83), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT83), .B1(new_n390), .B2(new_n394), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n191), .A2(G125), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n222), .A2(new_n224), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n321), .A2(G224), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n379), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n379), .B2(new_n384), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(new_n391), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n397), .A2(new_n398), .A3(new_n403), .A4(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n406), .B2(new_n393), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n390), .A2(KEYINPUT83), .A3(new_n394), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n411), .A2(new_n403), .A3(new_n408), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT84), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n371), .A2(new_n378), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n377), .B1(new_n416), .B2(KEYINPUT85), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n388), .B(KEYINPUT8), .Z(new_n418));
  NOR2_X1   g232(.A1(new_n377), .A2(KEYINPUT85), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(KEYINPUT79), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n417), .B(new_n418), .C1(new_n369), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT86), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n422), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n402), .A2(KEYINPUT7), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n401), .B1(KEYINPUT87), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n427));
  XOR2_X1   g241(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND4_X1  g242(.A1(new_n423), .A2(new_n424), .A3(new_n392), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n266), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n353), .B1(new_n415), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n353), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n433), .B(new_n430), .C1(new_n409), .C2(new_n414), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n343), .B(new_n352), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n339), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n400), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n371), .A2(new_n378), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n382), .A2(new_n383), .A3(new_n191), .ZN(new_n443));
  INV_X1    g257(.A(new_n227), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n190), .B1(G128), .B2(new_n218), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n224), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n369), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n321), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n400), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n371), .B2(new_n378), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n369), .A2(new_n446), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n227), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT12), .B(new_n227), .C1(new_n454), .C2(new_n455), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n442), .A2(new_n447), .A3(new_n443), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n227), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n451), .B1(new_n462), .B2(new_n448), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n439), .B(new_n266), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n448), .A3(new_n451), .ZN(new_n465));
  INV_X1    g279(.A(new_n448), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n458), .B2(new_n459), .ZN(new_n467));
  OAI211_X1 g281(.A(G469), .B(new_n465), .C1(new_n467), .C2(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(G469), .A2(G902), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G221), .ZN(new_n471));
  XOR2_X1   g285(.A(KEYINPUT9), .B(G234), .Z(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(new_n266), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n312), .A2(new_n314), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n241), .A2(G214), .ZN(new_n482));
  INV_X1    g296(.A(G143), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(KEYINPUT88), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(G214), .A3(new_n241), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(KEYINPUT17), .A3(G131), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n202), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n481), .B(new_n488), .C1(new_n490), .C2(KEYINPUT17), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n303), .B(new_n216), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(new_n202), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(G131), .ZN(new_n495));
  OAI221_X1 g309(.A(new_n492), .B1(new_n487), .B2(new_n494), .C1(new_n495), .C2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n354), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n499), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n303), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n307), .B1(new_n504), .B2(G146), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n496), .B(new_n501), .C1(new_n505), .C2(new_n489), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n507), .A2(G475), .A3(G902), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n499), .A2(KEYINPUT90), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n497), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n511), .B2(new_n497), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G475), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G122), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT91), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n360), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(G116), .B2(new_n516), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n519), .B(new_n520), .Z(new_n521));
  NAND2_X1  g335(.A1(new_n203), .A2(new_n205), .ZN(new_n522));
  XNOR2_X1  g336(.A(G128), .B(G143), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n520), .B(G107), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(KEYINPUT13), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n215), .A2(KEYINPUT13), .A3(G143), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n193), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n527), .A2(new_n529), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n472), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n532), .A2(new_n290), .A3(G953), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n525), .B2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n266), .ZN(new_n539));
  INV_X1    g353(.A(G478), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n539), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n515), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n480), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n341), .A2(new_n436), .A3(new_n438), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(G101), .ZN(G3));
  NAND2_X1  g361(.A1(new_n264), .A2(new_n266), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G472), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n267), .ZN(new_n550));
  INV_X1    g364(.A(new_n338), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n480), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT93), .Z(new_n553));
  OAI211_X1 g367(.A(new_n342), .B(new_n352), .C1(new_n432), .C2(new_n434), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n510), .A2(new_n514), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n538), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n535), .A2(KEYINPUT33), .A3(new_n537), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n540), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n538), .A2(new_n540), .A3(new_n266), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n540), .A2(new_n266), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(KEYINPUT34), .B(G104), .Z(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(G6));
  AND2_X1   g382(.A1(new_n413), .A2(KEYINPUT84), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n413), .A2(KEYINPUT84), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n431), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n433), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n415), .A2(new_n353), .A3(new_n431), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n351), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n555), .A2(new_n543), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n553), .A2(new_n342), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G107), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G9));
  INV_X1    g393(.A(new_n550), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n333), .A2(new_n334), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n291), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n329), .A2(new_n583), .A3(new_n323), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n327), .B(new_n328), .C1(KEYINPUT36), .C2(new_n324), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n336), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n589), .A3(new_n336), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n582), .A2(KEYINPUT96), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(new_n335), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n436), .A2(new_n545), .A3(new_n580), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT37), .B(G110), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G12));
  AND2_X1   g413(.A1(new_n289), .A2(new_n479), .ZN(new_n600));
  INV_X1    g414(.A(new_n342), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n572), .B2(new_n573), .ZN(new_n602));
  INV_X1    g416(.A(G900), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n348), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n347), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n542), .A2(new_n510), .A3(new_n514), .A4(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT97), .Z(new_n608));
  AND4_X1   g422(.A1(new_n596), .A2(new_n600), .A3(new_n602), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n215), .ZN(G30));
  XNOR2_X1  g424(.A(new_n605), .B(KEYINPUT39), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT40), .B1(new_n480), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n593), .A2(new_n335), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n614));
  INV_X1    g428(.A(new_n611), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n479), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n342), .A2(new_n612), .A3(new_n613), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n247), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n279), .A2(new_n259), .A3(new_n281), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(KEYINPUT98), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n619), .A2(KEYINPUT98), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n622), .B2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n269), .A3(new_n288), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n623), .A2(new_n269), .A3(KEYINPUT99), .A4(new_n288), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n572), .A2(new_n573), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT38), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n515), .A2(new_n543), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n617), .A2(new_n628), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G143), .ZN(G45));
  OAI21_X1  g447(.A(new_n342), .B1(new_n432), .B2(new_n434), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n289), .A2(new_n479), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n564), .A2(new_n605), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n634), .A2(new_n635), .A3(new_n595), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n216), .ZN(G48));
  OR2_X1    g453(.A1(new_n460), .A2(new_n463), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n266), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G469), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n642), .A2(new_n474), .A3(new_n464), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n289), .A2(new_n338), .A3(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n554), .A2(new_n644), .A3(new_n564), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT41), .B(G113), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G15));
  NAND2_X1  g461(.A1(new_n515), .A2(new_n542), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n554), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(G116), .Z(G18));
  OAI211_X1 g464(.A(new_n342), .B(new_n643), .C1(new_n432), .C2(new_n434), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT100), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n629), .A2(new_n653), .A3(new_n342), .A4(new_n643), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n544), .B1(new_n591), .B2(new_n594), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n656), .A2(new_n289), .A3(new_n352), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G119), .ZN(G21));
  OAI211_X1 g473(.A(new_n342), .B(new_n631), .C1(new_n432), .C2(new_n434), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n629), .A2(KEYINPUT101), .A3(new_n342), .A4(new_n631), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n282), .A2(new_n257), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n252), .B1(new_n665), .B2(new_n245), .ZN(new_n666));
  INV_X1    g480(.A(new_n248), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n265), .B(new_n266), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n549), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n338), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n643), .A2(new_n352), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n664), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G122), .ZN(G24));
  INV_X1    g488(.A(new_n613), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n669), .A2(new_n636), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n652), .B2(new_n654), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n305), .ZN(G27));
  NAND4_X1  g492(.A1(new_n572), .A2(new_n636), .A3(new_n342), .A4(new_n573), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n475), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n289), .A2(new_n338), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n680), .A2(KEYINPUT42), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n679), .B2(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G131), .ZN(G33));
  AND2_X1   g502(.A1(new_n683), .A2(new_n608), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n572), .A2(new_n342), .A3(new_n573), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT102), .B(G134), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G36));
  OAI21_X1  g508(.A(new_n465), .B1(new_n467), .B2(new_n451), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n697));
  OR3_X1    g511(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n439), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(KEYINPUT46), .A3(new_n469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n464), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT46), .B1(new_n701), .B2(new_n469), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n474), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n615), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n515), .A2(new_n563), .ZN(new_n709));
  NAND2_X1  g523(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n712));
  OAI21_X1  g526(.A(new_n711), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n550), .A3(new_n675), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n707), .B1(new_n708), .B2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n715), .B(new_n691), .C1(new_n708), .C2(new_n714), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G137), .ZN(G39));
  XNOR2_X1  g531(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n706), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n706), .A2(new_n718), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n289), .A2(new_n338), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n680), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G140), .ZN(G42));
  NAND3_X1  g539(.A1(new_n613), .A2(new_n681), .A3(new_n606), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n626), .B2(new_n627), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n664), .A2(KEYINPUT110), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT110), .B1(new_n664), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OR3_X1    g544(.A1(new_n677), .A2(new_n609), .A3(new_n638), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT52), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n733));
  INV_X1    g547(.A(new_n645), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n673), .A3(new_n687), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n648), .B(KEYINPUT107), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n435), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n575), .B(KEYINPUT107), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n574), .A2(new_n740), .A3(KEYINPUT108), .A4(new_n343), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n552), .ZN(new_n742));
  INV_X1    g556(.A(new_n564), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n436), .A2(new_n552), .A3(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n742), .A2(new_n744), .A3(new_n546), .A4(new_n597), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n600), .A2(new_n656), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n669), .A2(new_n681), .A3(new_n743), .A4(new_n675), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n605), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n746), .B(new_n691), .C1(new_n749), .C2(new_n689), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n748), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n606), .A3(new_n691), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .A3(new_n692), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n745), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n677), .A2(new_n609), .A3(new_n638), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n756), .C1(new_n729), .C2(new_n728), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n732), .A2(new_n736), .A3(new_n754), .A4(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT53), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT54), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n762));
  INV_X1    g576(.A(new_n347), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n713), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n671), .ZN(new_n765));
  INV_X1    g579(.A(new_n630), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n601), .A4(new_n643), .ZN(new_n767));
  NAND2_X1  g581(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n767), .B(new_n768), .Z(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(KEYINPUT112), .B2(KEYINPUT50), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n642), .A2(new_n464), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT106), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n474), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n691), .B(new_n765), .C1(new_n722), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n691), .A2(new_n643), .ZN(new_n776));
  OR4_X1    g590(.A1(new_n551), .A2(new_n776), .A3(new_n628), .A4(new_n347), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(new_n555), .A3(new_n563), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n764), .A2(new_n643), .A3(new_n691), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n669), .A2(new_n675), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n762), .B1(new_n775), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n732), .A2(new_n754), .A3(new_n757), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n735), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n670), .B1(new_n662), .B2(new_n663), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n645), .B1(new_n788), .B2(new_n672), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n687), .A4(new_n733), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n790), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n785), .A2(new_n791), .B1(new_n758), .B2(new_n759), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n777), .A2(new_n564), .ZN(new_n795));
  NOR2_X1   g609(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT114), .Z(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n779), .A2(new_n339), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n779), .B2(new_n339), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n765), .A2(new_n655), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n795), .A2(new_n802), .A3(new_n344), .A4(new_n803), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT116), .Z(new_n805));
  NAND4_X1  g619(.A1(new_n761), .A2(new_n784), .A3(new_n794), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n808));
  AOI211_X1 g622(.A(new_n762), .B(new_n775), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n806), .A2(new_n809), .B1(G952), .B2(G953), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n772), .B(KEYINPUT49), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n473), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n343), .A3(new_n626), .A4(new_n627), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n813), .A2(new_n551), .A3(new_n630), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n810), .B1(new_n709), .B2(new_n814), .ZN(G75));
  NOR2_X1   g629(.A1(new_n321), .A2(G952), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(G210), .ZN(new_n818));
  INV_X1    g632(.A(new_n757), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n664), .A2(new_n727), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n664), .A2(KEYINPUT110), .A3(new_n727), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n756), .B1(new_n824), .B2(new_n755), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n791), .A3(new_n754), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n758), .A2(new_n759), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n818), .B(new_n266), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n397), .A2(new_n408), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(new_n403), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT55), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n817), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT56), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n829), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n827), .A2(new_n828), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n836), .A3(G210), .A4(G902), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n833), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT118), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(G210), .A3(G902), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT56), .B1(new_n842), .B2(KEYINPUT117), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n839), .A4(new_n833), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n834), .B1(new_n841), .B2(new_n845), .ZN(G51));
  NAND2_X1  g660(.A1(new_n469), .A2(KEYINPUT57), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n469), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g662(.A(new_n794), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n792), .A2(new_n793), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n640), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n792), .A2(new_n266), .A3(new_n701), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n816), .B1(new_n852), .B2(new_n853), .ZN(G54));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(KEYINPUT58), .B2(G475), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(KEYINPUT58), .A3(G475), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n838), .A2(G902), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(new_n507), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n507), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n860), .A2(new_n861), .A3(new_n816), .ZN(G60));
  XNOR2_X1  g676(.A(new_n562), .B(KEYINPUT59), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n557), .A2(new_n558), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT120), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n866), .C1(new_n849), .C2(new_n850), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n761), .B2(new_n794), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n867), .B(new_n817), .C1(new_n868), .C2(new_n866), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(G63));
  INV_X1    g684(.A(new_n330), .ZN(new_n871));
  NAND2_X1  g685(.A1(G217), .A2(G902), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT60), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n792), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n873), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n838), .A2(new_n586), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n876), .A3(new_n817), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT61), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n877), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(G66));
  INV_X1    g695(.A(G224), .ZN(new_n882));
  OAI21_X1  g696(.A(G953), .B1(new_n349), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n745), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n789), .A3(new_n733), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n886), .B2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n831), .B1(G898), .B2(new_n321), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(G69));
  AND2_X1   g703(.A1(new_n724), .A2(new_n716), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n755), .A2(new_n632), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n341), .A2(new_n438), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n480), .A2(new_n611), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n738), .A2(new_n564), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n691), .A4(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT123), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n890), .A2(new_n893), .A3(new_n900), .A4(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n504), .B(KEYINPUT122), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n271), .B(new_n903), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n321), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(G227), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n603), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n716), .A2(new_n755), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n716), .A2(KEYINPUT124), .A3(new_n755), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n910), .A2(new_n724), .A3(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n664), .A2(new_n340), .A3(new_n615), .A4(new_n706), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n692), .A2(new_n687), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT125), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n321), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(G227), .B2(new_n321), .ZN(new_n918));
  OAI221_X1 g732(.A(new_n905), .B1(new_n321), .B2(new_n907), .C1(new_n918), .C2(new_n904), .ZN(G72));
  INV_X1    g733(.A(new_n272), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(new_n920), .A3(new_n901), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n912), .A2(new_n915), .A3(new_n259), .A4(new_n913), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n273), .B(new_n885), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n265), .A2(new_n266), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n618), .A2(new_n273), .A3(KEYINPUT127), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n273), .A2(KEYINPUT127), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n760), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n618), .A2(new_n273), .A3(new_n926), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n923), .A2(new_n929), .A3(new_n816), .A4(new_n930), .ZN(G57));
endmodule


