

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707;

  NAND2_X1 U367 ( .A1(n627), .A2(n626), .ZN(n629) );
  INV_X1 U368 ( .A(G953), .ZN(n696) );
  NOR2_X2 U369 ( .A1(n498), .A2(n552), .ZN(n500) );
  XNOR2_X2 U370 ( .A(n466), .B(n467), .ZN(n491) );
  AND2_X2 U371 ( .A1(n508), .A2(n465), .ZN(n466) );
  XNOR2_X2 U372 ( .A(n529), .B(n352), .ZN(n630) );
  NAND2_X1 U373 ( .A1(n503), .A2(n494), .ZN(n495) );
  NOR2_X1 U374 ( .A1(n571), .A2(n570), .ZN(n572) );
  AND2_X1 U375 ( .A1(n358), .A2(n705), .ZN(n399) );
  XNOR2_X1 U376 ( .A(KEYINPUT32), .B(n490), .ZN(n705) );
  NOR2_X1 U377 ( .A1(n532), .A2(n538), .ZN(n533) );
  XNOR2_X1 U378 ( .A(n354), .B(n353), .ZN(n620) );
  NOR2_X1 U379 ( .A1(n616), .A2(n615), .ZN(n354) );
  XNOR2_X1 U380 ( .A(n462), .B(n461), .ZN(n473) );
  XNOR2_X1 U381 ( .A(n416), .B(G104), .ZN(n443) );
  XOR2_X1 U382 ( .A(G119), .B(KEYINPUT3), .Z(n406) );
  XNOR2_X1 U383 ( .A(G113), .B(G122), .ZN(n416) );
  XNOR2_X1 U384 ( .A(n456), .B(n443), .ZN(n349) );
  BUF_X1 U385 ( .A(n660), .Z(n672) );
  XNOR2_X2 U386 ( .A(n414), .B(n376), .ZN(n636) );
  XNOR2_X2 U387 ( .A(n488), .B(n487), .ZN(n529) );
  XNOR2_X1 U388 ( .A(n381), .B(n380), .ZN(n619) );
  INV_X1 U389 ( .A(KEYINPUT99), .ZN(n380) );
  OR2_X1 U390 ( .A1(n609), .A2(n604), .ZN(n381) );
  AND2_X1 U391 ( .A1(n386), .A2(n372), .ZN(n368) );
  XNOR2_X1 U392 ( .A(n539), .B(KEYINPUT38), .ZN(n616) );
  OR2_X1 U393 ( .A1(G237), .A2(G902), .ZN(n424) );
  XNOR2_X1 U394 ( .A(n410), .B(KEYINPUT5), .ZN(n379) );
  XNOR2_X1 U395 ( .A(G113), .B(G116), .ZN(n410) );
  XNOR2_X1 U396 ( .A(n345), .B(n405), .ZN(n481) );
  XNOR2_X1 U397 ( .A(G131), .B(G134), .ZN(n405) );
  XOR2_X1 U398 ( .A(KEYINPUT17), .B(KEYINPUT82), .Z(n418) );
  INV_X1 U399 ( .A(KEYINPUT101), .ZN(n396) );
  XNOR2_X1 U400 ( .A(n447), .B(n446), .ZN(n510) );
  NOR2_X1 U401 ( .A1(G902), .A2(n664), .ZN(n447) );
  NOR2_X1 U402 ( .A1(G902), .A2(n656), .ZN(n488) );
  INV_X1 U403 ( .A(KEYINPUT16), .ZN(n415) );
  XOR2_X1 U404 ( .A(G137), .B(G140), .Z(n480) );
  XOR2_X1 U405 ( .A(G119), .B(G110), .Z(n402) );
  XOR2_X1 U406 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n451) );
  XNOR2_X1 U407 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n450) );
  XNOR2_X1 U408 ( .A(n456), .B(KEYINPUT96), .ZN(n384) );
  XNOR2_X1 U409 ( .A(n442), .B(n355), .ZN(n691) );
  XNOR2_X1 U410 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n481), .B(n389), .ZN(n690) );
  INV_X1 U412 ( .A(n480), .ZN(n389) );
  NOR2_X2 U413 ( .A1(n651), .A2(n575), .ZN(n660) );
  XNOR2_X1 U414 ( .A(n523), .B(n524), .ZN(n532) );
  XNOR2_X1 U415 ( .A(n505), .B(n504), .ZN(n638) );
  XOR2_X1 U416 ( .A(KEYINPUT104), .B(n521), .Z(n346) );
  AND2_X1 U417 ( .A1(n522), .A2(n387), .ZN(n386) );
  INV_X1 U418 ( .A(n525), .ZN(n387) );
  XNOR2_X1 U419 ( .A(n375), .B(n516), .ZN(n522) );
  XNOR2_X1 U420 ( .A(n458), .B(n457), .ZN(n511) );
  XNOR2_X1 U421 ( .A(n690), .B(n388), .ZN(n656) );
  XNOR2_X1 U422 ( .A(n486), .B(n479), .ZN(n388) );
  XNOR2_X1 U423 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U424 ( .A(G146), .ZN(n484) );
  NOR2_X1 U425 ( .A1(G952), .A2(n696), .ZN(n676) );
  INV_X1 U426 ( .A(n619), .ZN(n536) );
  XOR2_X1 U427 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n460) );
  INV_X1 U428 ( .A(KEYINPUT107), .ZN(n353) );
  INV_X1 U429 ( .A(KEYINPUT39), .ZN(n372) );
  NOR2_X1 U430 ( .A1(n386), .A2(n372), .ZN(n371) );
  AND2_X1 U431 ( .A1(n346), .A2(n374), .ZN(n373) );
  INV_X1 U432 ( .A(n616), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n412) );
  XNOR2_X1 U434 ( .A(n409), .B(n411), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n417), .B(n379), .ZN(n378) );
  XNOR2_X1 U436 ( .A(G131), .B(G143), .ZN(n438) );
  XNOR2_X1 U437 ( .A(G101), .B(G110), .ZN(n390) );
  XNOR2_X1 U438 ( .A(n392), .B(KEYINPUT70), .ZN(n391) );
  INV_X1 U439 ( .A(KEYINPUT81), .ZN(n392) );
  XNOR2_X1 U440 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U441 ( .A(G107), .B(G104), .ZN(n482) );
  XNOR2_X1 U442 ( .A(n677), .B(n400), .ZN(n581) );
  XNOR2_X1 U443 ( .A(n421), .B(n420), .ZN(n400) );
  XNOR2_X1 U444 ( .A(n419), .B(KEYINPUT18), .ZN(n420) );
  INV_X1 U445 ( .A(n532), .ZN(n640) );
  XNOR2_X1 U446 ( .A(n393), .B(KEYINPUT73), .ZN(n357) );
  INV_X1 U447 ( .A(KEYINPUT45), .ZN(n393) );
  INV_X1 U448 ( .A(KEYINPUT1), .ZN(n352) );
  XNOR2_X1 U449 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n425) );
  INV_X1 U450 ( .A(G472), .ZN(n376) );
  NOR2_X1 U451 ( .A1(G902), .A2(n413), .ZN(n414) );
  INV_X1 U452 ( .A(n636), .ZN(n527) );
  XNOR2_X1 U453 ( .A(n691), .B(n472), .ZN(n356) );
  XNOR2_X1 U454 ( .A(n360), .B(n403), .ZN(n471) );
  XNOR2_X1 U455 ( .A(n480), .B(n402), .ZN(n472) );
  XNOR2_X1 U456 ( .A(n385), .B(n383), .ZN(n670) );
  XNOR2_X1 U457 ( .A(n452), .B(n384), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n453), .B(n455), .ZN(n385) );
  XNOR2_X1 U459 ( .A(n533), .B(n362), .ZN(n706) );
  INV_X1 U460 ( .A(KEYINPUT42), .ZN(n362) );
  XNOR2_X1 U461 ( .A(n535), .B(KEYINPUT40), .ZN(n707) );
  XNOR2_X1 U462 ( .A(KEYINPUT31), .B(n506), .ZN(n608) );
  NAND2_X1 U463 ( .A1(n386), .A2(n346), .ZN(n551) );
  XNOR2_X1 U464 ( .A(n513), .B(n382), .ZN(n609) );
  INV_X1 U465 ( .A(KEYINPUT98), .ZN(n382) );
  NOR2_X1 U466 ( .A1(n511), .A2(n512), .ZN(n604) );
  XNOR2_X1 U467 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U468 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U469 ( .A(KEYINPUT4), .B(n448), .Z(n345) );
  XNOR2_X1 U470 ( .A(n391), .B(n390), .ZN(n479) );
  XOR2_X1 U471 ( .A(n415), .B(n479), .Z(n347) );
  NAND2_X1 U472 ( .A1(G224), .A2(n696), .ZN(n348) );
  AND2_X1 U473 ( .A1(n559), .A2(n558), .ZN(n350) );
  AND2_X1 U474 ( .A1(G210), .A2(n424), .ZN(n351) );
  XNOR2_X1 U475 ( .A(n401), .B(n347), .ZN(n677) );
  XNOR2_X1 U476 ( .A(n397), .B(n396), .ZN(n395) );
  NOR2_X2 U477 ( .A1(n676), .A2(n667), .ZN(n668) );
  XNOR2_X1 U478 ( .A(n366), .B(n404), .ZN(n365) );
  NAND2_X1 U479 ( .A1(n365), .A2(n350), .ZN(n364) );
  NOR2_X1 U480 ( .A1(n586), .A2(n676), .ZN(n587) );
  NOR2_X1 U481 ( .A1(n578), .A2(n676), .ZN(n580) );
  XNOR2_X2 U482 ( .A(n423), .B(n351), .ZN(n539) );
  XNOR2_X1 U483 ( .A(n356), .B(n471), .ZN(n674) );
  NAND2_X1 U484 ( .A1(n369), .A2(n367), .ZN(n534) );
  NOR2_X1 U485 ( .A1(n373), .A2(n372), .ZN(n370) );
  XNOR2_X2 U486 ( .A(n394), .B(n357), .ZN(n681) );
  NAND2_X1 U487 ( .A1(n539), .A2(n540), .ZN(n426) );
  NOR2_X1 U488 ( .A1(n703), .A2(n359), .ZN(n358) );
  INV_X1 U489 ( .A(n597), .ZN(n359) );
  NAND2_X1 U490 ( .A1(n468), .A2(G221), .ZN(n360) );
  NOR2_X1 U491 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U492 ( .A1(n361), .A2(n681), .ZN(n573) );
  XNOR2_X1 U493 ( .A(n572), .B(KEYINPUT74), .ZN(n361) );
  NOR2_X2 U494 ( .A1(n571), .A2(n613), .ZN(n694) );
  NAND2_X1 U495 ( .A1(n565), .A2(n614), .ZN(n571) );
  XNOR2_X1 U496 ( .A(n349), .B(n417), .ZN(n401) );
  NAND2_X1 U497 ( .A1(n707), .A2(n706), .ZN(n366) );
  XNOR2_X1 U498 ( .A(n364), .B(n363), .ZN(n565) );
  INV_X1 U499 ( .A(KEYINPUT48), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n534), .A2(n604), .ZN(n535) );
  NAND2_X1 U501 ( .A1(n368), .A2(n373), .ZN(n367) );
  NAND2_X1 U502 ( .A1(n636), .A2(n540), .ZN(n375) );
  NAND2_X1 U503 ( .A1(n398), .A2(n395), .ZN(n394) );
  NOR2_X1 U504 ( .A1(n515), .A2(n588), .ZN(n397) );
  XNOR2_X1 U505 ( .A(n399), .B(KEYINPUT44), .ZN(n398) );
  XNOR2_X1 U506 ( .A(n345), .B(n348), .ZN(n421) );
  NAND2_X1 U507 ( .A1(n503), .A2(n636), .ZN(n505) );
  XNOR2_X2 U508 ( .A(n495), .B(KEYINPUT33), .ZN(n624) );
  XOR2_X1 U509 ( .A(n470), .B(n469), .Z(n403) );
  XOR2_X1 U510 ( .A(KEYINPUT46), .B(KEYINPUT76), .Z(n404) );
  XNOR2_X1 U511 ( .A(n426), .B(n425), .ZN(n537) );
  INV_X1 U512 ( .A(KEYINPUT72), .ZN(n555) );
  XNOR2_X1 U513 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT86), .ZN(n461) );
  INV_X1 U515 ( .A(KEYINPUT92), .ZN(n504) );
  XNOR2_X1 U516 ( .A(KEYINPUT13), .B(G475), .ZN(n446) );
  XNOR2_X1 U517 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X2 U518 ( .A(G143), .B(G128), .Z(n448) );
  XOR2_X1 U519 ( .A(KEYINPUT68), .B(n406), .Z(n417) );
  XOR2_X1 U520 ( .A(KEYINPUT91), .B(G137), .Z(n408) );
  XNOR2_X1 U521 ( .A(G101), .B(G146), .ZN(n407) );
  XNOR2_X1 U522 ( .A(n408), .B(n407), .ZN(n409) );
  NOR2_X1 U523 ( .A1(G953), .A2(G237), .ZN(n435) );
  NAND2_X1 U524 ( .A1(n435), .A2(G210), .ZN(n411) );
  XNOR2_X1 U525 ( .A(n481), .B(n412), .ZN(n413) );
  XNOR2_X1 U526 ( .A(n413), .B(KEYINPUT62), .ZN(n577) );
  XOR2_X1 U527 ( .A(n527), .B(KEYINPUT6), .Z(n542) );
  INV_X1 U528 ( .A(n542), .ZN(n494) );
  INV_X1 U529 ( .A(KEYINPUT22), .ZN(n467) );
  XOR2_X1 U530 ( .A(G116), .B(G107), .Z(n456) );
  XOR2_X1 U531 ( .A(G146), .B(G125), .Z(n442) );
  XNOR2_X1 U532 ( .A(n442), .B(n418), .ZN(n419) );
  XNOR2_X2 U533 ( .A(G902), .B(KEYINPUT15), .ZN(n422) );
  XNOR2_X2 U534 ( .A(n422), .B(KEYINPUT80), .ZN(n575) );
  NAND2_X1 U535 ( .A1(n581), .A2(n575), .ZN(n423) );
  NAND2_X1 U536 ( .A1(G214), .A2(n424), .ZN(n540) );
  XOR2_X1 U537 ( .A(KEYINPUT14), .B(KEYINPUT83), .Z(n428) );
  NAND2_X1 U538 ( .A1(G234), .A2(G237), .ZN(n427) );
  XNOR2_X1 U539 ( .A(n428), .B(n427), .ZN(n430) );
  AND2_X1 U540 ( .A1(G953), .A2(n430), .ZN(n429) );
  NAND2_X1 U541 ( .A1(G902), .A2(n429), .ZN(n517) );
  NOR2_X1 U542 ( .A1(G898), .A2(n517), .ZN(n432) );
  NAND2_X1 U543 ( .A1(G952), .A2(n430), .ZN(n646) );
  NOR2_X1 U544 ( .A1(G953), .A2(n646), .ZN(n431) );
  XNOR2_X1 U545 ( .A(KEYINPUT84), .B(n431), .ZN(n520) );
  NOR2_X1 U546 ( .A1(n432), .A2(n520), .ZN(n433) );
  NOR2_X2 U547 ( .A1(n537), .A2(n433), .ZN(n434) );
  XNOR2_X2 U548 ( .A(n434), .B(KEYINPUT0), .ZN(n508) );
  XOR2_X1 U549 ( .A(KEYINPUT12), .B(KEYINPUT93), .Z(n437) );
  NAND2_X1 U550 ( .A1(G214), .A2(n435), .ZN(n436) );
  XNOR2_X1 U551 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U552 ( .A(KEYINPUT11), .B(G140), .Z(n439) );
  XNOR2_X1 U553 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U554 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U555 ( .A(n691), .B(n443), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n445), .B(n444), .ZN(n664) );
  XNOR2_X1 U557 ( .A(n448), .B(G134), .ZN(n449) );
  XNOR2_X1 U558 ( .A(n449), .B(G122), .ZN(n453) );
  XNOR2_X1 U559 ( .A(n451), .B(n450), .ZN(n452) );
  NAND2_X1 U560 ( .A1(G234), .A2(n696), .ZN(n454) );
  XOR2_X1 U561 ( .A(KEYINPUT8), .B(n454), .Z(n468) );
  NAND2_X1 U562 ( .A1(G217), .A2(n468), .ZN(n455) );
  NOR2_X1 U563 ( .A1(G902), .A2(n670), .ZN(n458) );
  XNOR2_X1 U564 ( .A(KEYINPUT97), .B(G478), .ZN(n457) );
  NOR2_X1 U565 ( .A1(n510), .A2(n511), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n459), .B(KEYINPUT100), .ZN(n617) );
  NAND2_X1 U567 ( .A1(G234), .A2(n575), .ZN(n462) );
  NAND2_X1 U568 ( .A1(n473), .A2(G221), .ZN(n463) );
  XNOR2_X1 U569 ( .A(n463), .B(KEYINPUT90), .ZN(n464) );
  XOR2_X1 U570 ( .A(KEYINPUT21), .B(n464), .Z(n626) );
  AND2_X1 U571 ( .A1(n617), .A2(n626), .ZN(n465) );
  NOR2_X2 U572 ( .A1(n494), .A2(n491), .ZN(n501) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n470) );
  XNOR2_X1 U574 ( .A(G128), .B(KEYINPUT85), .ZN(n469) );
  NOR2_X1 U575 ( .A1(G902), .A2(n674), .ZN(n478) );
  XOR2_X1 U576 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n475) );
  NAND2_X1 U577 ( .A1(G217), .A2(n473), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U579 ( .A(n476), .B(KEYINPUT25), .ZN(n477) );
  XNOR2_X2 U580 ( .A(n478), .B(n477), .ZN(n627) );
  NAND2_X1 U581 ( .A1(G227), .A2(n696), .ZN(n483) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(G469), .ZN(n487) );
  NOR2_X1 U583 ( .A1(n627), .A2(n630), .ZN(n489) );
  NAND2_X1 U584 ( .A1(n501), .A2(n489), .ZN(n490) );
  INV_X1 U585 ( .A(n630), .ZN(n548) );
  NOR2_X1 U586 ( .A1(n491), .A2(n548), .ZN(n493) );
  NOR2_X1 U587 ( .A1(n627), .A2(n636), .ZN(n492) );
  NAND2_X1 U588 ( .A1(n493), .A2(n492), .ZN(n597) );
  NOR2_X1 U589 ( .A1(n630), .A2(n629), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n624), .A2(n508), .ZN(n497) );
  XOR2_X1 U591 ( .A(KEYINPUT69), .B(KEYINPUT34), .Z(n496) );
  XNOR2_X1 U592 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U593 ( .A1(n511), .A2(n510), .ZN(n552) );
  XNOR2_X1 U594 ( .A(KEYINPUT75), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U595 ( .A(n500), .B(n499), .ZN(n703) );
  NAND2_X1 U596 ( .A1(n627), .A2(n501), .ZN(n502) );
  NOR2_X1 U597 ( .A1(n548), .A2(n502), .ZN(n588) );
  NAND2_X1 U598 ( .A1(n508), .A2(n638), .ZN(n506) );
  INV_X1 U599 ( .A(n629), .ZN(n507) );
  NAND2_X1 U600 ( .A1(n529), .A2(n507), .ZN(n521) );
  NAND2_X1 U601 ( .A1(n527), .A2(n508), .ZN(n509) );
  NOR2_X1 U602 ( .A1(n521), .A2(n509), .ZN(n594) );
  NOR2_X1 U603 ( .A1(n608), .A2(n594), .ZN(n514) );
  INV_X1 U604 ( .A(n510), .ZN(n512) );
  NAND2_X1 U605 ( .A1(n512), .A2(n511), .ZN(n513) );
  NOR2_X1 U606 ( .A1(n514), .A2(n536), .ZN(n515) );
  XNOR2_X1 U607 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n516) );
  NOR2_X1 U608 ( .A1(G900), .A2(n517), .ZN(n518) );
  XNOR2_X1 U609 ( .A(n518), .B(KEYINPUT102), .ZN(n519) );
  NOR2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n525) );
  NAND2_X1 U611 ( .A1(n609), .A2(n534), .ZN(n568) );
  INV_X1 U612 ( .A(n568), .ZN(n613) );
  XOR2_X1 U613 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n524) );
  INV_X1 U614 ( .A(n540), .ZN(n615) );
  NAND2_X1 U615 ( .A1(n620), .A2(n617), .ZN(n523) );
  NOR2_X1 U616 ( .A1(n627), .A2(n525), .ZN(n526) );
  NAND2_X1 U617 ( .A1(n626), .A2(n526), .ZN(n541) );
  NOR2_X1 U618 ( .A1(n527), .A2(n541), .ZN(n528) );
  XNOR2_X1 U619 ( .A(KEYINPUT28), .B(n528), .ZN(n531) );
  XNOR2_X1 U620 ( .A(n529), .B(KEYINPUT106), .ZN(n530) );
  NAND2_X1 U621 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U622 ( .A1(n537), .A2(n538), .ZN(n601) );
  NAND2_X1 U623 ( .A1(n619), .A2(n601), .ZN(n550) );
  OR2_X1 U624 ( .A1(n550), .A2(KEYINPUT47), .ZN(n559) );
  BUF_X1 U625 ( .A(n539), .Z(n562) );
  NAND2_X1 U626 ( .A1(n604), .A2(n540), .ZN(n545) );
  NOR2_X1 U627 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n543), .B(KEYINPUT103), .ZN(n544) );
  NOR2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n562), .A2(n560), .ZN(n547) );
  XNOR2_X1 U631 ( .A(KEYINPUT77), .B(KEYINPUT36), .ZN(n546) );
  XNOR2_X1 U632 ( .A(n547), .B(n546), .ZN(n549) );
  NAND2_X1 U633 ( .A1(n549), .A2(n548), .ZN(n612) );
  NAND2_X1 U634 ( .A1(n550), .A2(KEYINPUT47), .ZN(n554) );
  NOR2_X1 U635 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U636 ( .A1(n562), .A2(n553), .ZN(n600) );
  NAND2_X1 U637 ( .A1(n554), .A2(n600), .ZN(n556) );
  AND2_X1 U638 ( .A1(n612), .A2(n557), .ZN(n558) );
  NAND2_X1 U639 ( .A1(n630), .A2(n560), .ZN(n561) );
  XNOR2_X1 U640 ( .A(n561), .B(KEYINPUT43), .ZN(n564) );
  INV_X1 U641 ( .A(n562), .ZN(n563) );
  NAND2_X1 U642 ( .A1(n564), .A2(n563), .ZN(n614) );
  NAND2_X1 U643 ( .A1(n681), .A2(n694), .ZN(n567) );
  INV_X1 U644 ( .A(KEYINPUT2), .ZN(n566) );
  NAND2_X1 U645 ( .A1(n567), .A2(n566), .ZN(n574) );
  NAND2_X1 U646 ( .A1(KEYINPUT2), .A2(n568), .ZN(n569) );
  XOR2_X1 U647 ( .A(KEYINPUT71), .B(n569), .Z(n570) );
  NAND2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n651) );
  NAND2_X1 U649 ( .A1(n660), .A2(G472), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U651 ( .A(KEYINPUT63), .B(KEYINPUT79), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n580), .B(n579), .ZN(G57) );
  XOR2_X1 U653 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n583) );
  XNOR2_X1 U654 ( .A(n581), .B(KEYINPUT55), .ZN(n582) );
  XNOR2_X1 U655 ( .A(n583), .B(n582), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n660), .A2(G210), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U659 ( .A(G101), .B(n588), .Z(G3) );
  XOR2_X1 U660 ( .A(G104), .B(KEYINPUT109), .Z(n590) );
  NAND2_X1 U661 ( .A1(n594), .A2(n604), .ZN(n589) );
  XNOR2_X1 U662 ( .A(n590), .B(n589), .ZN(G6) );
  XOR2_X1 U663 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n592) );
  XNOR2_X1 U664 ( .A(G107), .B(KEYINPUT26), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT110), .B(n593), .Z(n596) );
  NAND2_X1 U667 ( .A1(n594), .A2(n609), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n596), .B(n595), .ZN(G9) );
  XNOR2_X1 U669 ( .A(G110), .B(n597), .ZN(G12) );
  XOR2_X1 U670 ( .A(G128), .B(KEYINPUT29), .Z(n599) );
  NAND2_X1 U671 ( .A1(n601), .A2(n609), .ZN(n598) );
  XNOR2_X1 U672 ( .A(n599), .B(n598), .ZN(G30) );
  XNOR2_X1 U673 ( .A(G143), .B(n600), .ZN(G45) );
  NAND2_X1 U674 ( .A1(n601), .A2(n604), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT112), .ZN(n603) );
  XNOR2_X1 U676 ( .A(G146), .B(n603), .ZN(G48) );
  XOR2_X1 U677 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n606) );
  NAND2_X1 U678 ( .A1(n608), .A2(n604), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U680 ( .A(G113), .B(n607), .ZN(G15) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(G116), .ZN(G18) );
  XOR2_X1 U683 ( .A(G125), .B(KEYINPUT37), .Z(n611) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(G27) );
  XOR2_X1 U685 ( .A(G134), .B(n613), .Z(G36) );
  XNOR2_X1 U686 ( .A(G140), .B(n614), .ZN(G42) );
  AND2_X1 U687 ( .A1(n640), .A2(n624), .ZN(n649) );
  XNOR2_X1 U688 ( .A(KEYINPUT117), .B(KEYINPUT52), .ZN(n645) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(KEYINPUT116), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n643) );
  NOR2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT49), .B(n628), .ZN(n634) );
  XOR2_X1 U697 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n632) );
  NAND2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U700 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U702 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U703 ( .A(n639), .B(KEYINPUT51), .ZN(n641) );
  NAND2_X1 U704 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U705 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U706 ( .A(n645), .B(n644), .ZN(n647) );
  NOR2_X1 U707 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U708 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U709 ( .A(n650), .B(KEYINPUT118), .ZN(n652) );
  NAND2_X1 U710 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U711 ( .A1(n653), .A2(G953), .ZN(n654) );
  XNOR2_X1 U712 ( .A(n654), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U713 ( .A1(n672), .A2(G469), .ZN(n658) );
  XOR2_X1 U714 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n655) );
  NOR2_X1 U715 ( .A1(n676), .A2(n659), .ZN(G54) );
  NAND2_X1 U716 ( .A1(n660), .A2(G475), .ZN(n666) );
  XOR2_X1 U717 ( .A(KEYINPUT78), .B(KEYINPUT64), .Z(n662) );
  XNOR2_X1 U718 ( .A(KEYINPUT59), .B(KEYINPUT120), .ZN(n661) );
  XNOR2_X1 U719 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U720 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n668), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U722 ( .A1(G478), .A2(n672), .ZN(n669) );
  XNOR2_X1 U723 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U724 ( .A1(n676), .A2(n671), .ZN(G63) );
  NAND2_X1 U725 ( .A1(G217), .A2(n672), .ZN(n673) );
  XNOR2_X1 U726 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U727 ( .A1(n676), .A2(n675), .ZN(G66) );
  OR2_X1 U728 ( .A1(G898), .A2(n696), .ZN(n678) );
  NAND2_X1 U729 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U730 ( .A(n679), .B(KEYINPUT124), .ZN(n680) );
  XNOR2_X1 U731 ( .A(KEYINPUT123), .B(n680), .ZN(n689) );
  NAND2_X1 U732 ( .A1(n681), .A2(n696), .ZN(n682) );
  XNOR2_X1 U733 ( .A(n682), .B(KEYINPUT122), .ZN(n687) );
  XOR2_X1 U734 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n684) );
  NAND2_X1 U735 ( .A1(G224), .A2(G953), .ZN(n683) );
  XNOR2_X1 U736 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U737 ( .A1(n685), .A2(G898), .ZN(n686) );
  NAND2_X1 U738 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U739 ( .A(n689), .B(n688), .ZN(G69) );
  XOR2_X1 U740 ( .A(n690), .B(n691), .Z(n692) );
  XOR2_X1 U741 ( .A(KEYINPUT125), .B(n692), .Z(n698) );
  INV_X1 U742 ( .A(n698), .ZN(n693) );
  XOR2_X1 U743 ( .A(n693), .B(KEYINPUT126), .Z(n695) );
  XNOR2_X1 U744 ( .A(n695), .B(n694), .ZN(n697) );
  NAND2_X1 U745 ( .A1(n697), .A2(n696), .ZN(n702) );
  XOR2_X1 U746 ( .A(G227), .B(n698), .Z(n699) );
  NAND2_X1 U747 ( .A1(n699), .A2(G900), .ZN(n700) );
  NAND2_X1 U748 ( .A1(n700), .A2(G953), .ZN(n701) );
  NAND2_X1 U749 ( .A1(n702), .A2(n701), .ZN(G72) );
  XNOR2_X1 U750 ( .A(n703), .B(G122), .ZN(n704) );
  XNOR2_X1 U751 ( .A(n704), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U752 ( .A(G119), .B(n705), .ZN(G21) );
  XNOR2_X1 U753 ( .A(n706), .B(G137), .ZN(G39) );
  XNOR2_X1 U754 ( .A(n707), .B(G131), .ZN(G33) );
endmodule

