//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT64), .B(G77), .Z(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT67), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT66), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n211), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n209), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n224), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT68), .Z(G361));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT70), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G250), .ZN(new_n239));
  INV_X1    g0039(.A(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G226), .B(G232), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT71), .ZN(new_n251));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G20), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT72), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n262), .A2(new_n263), .B1(G1), .B2(G13), .ZN(new_n264));
  NAND4_X1  g0064(.A1(KEYINPUT72), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n266), .B1(new_n208), .B2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n261), .B1(new_n267), .B2(new_n257), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT7), .B1(new_n272), .B2(new_n209), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(G68), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT81), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n209), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G159), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT81), .A3(G159), .ZN(new_n285));
  XNOR2_X1  g0085(.A(G58), .B(G68), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n285), .B1(G20), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n278), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT16), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT82), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n274), .A2(new_n209), .A3(new_n275), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n294), .B2(new_n276), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n283), .A2(new_n285), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n286), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT82), .B(new_n289), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n290), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n266), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT80), .ZN(new_n303));
  OAI21_X1  g0103(.A(G68), .B1(new_n276), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n294), .A2(new_n303), .A3(new_n276), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n302), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n269), .B1(new_n301), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  INV_X1    g0110(.A(G223), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n270), .B2(new_n271), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT83), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G87), .ZN(new_n316));
  OAI211_X1 g0116(.A(G226), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n312), .B(KEYINPUT83), .C1(new_n271), .C2(new_n270), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n315), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G41), .ZN(new_n322));
  INV_X1    g0122(.A(G45), .ZN(new_n323));
  AOI21_X1  g0123(.A(G1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G41), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G1), .A3(G13), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n326), .A3(G274), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(G232), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n310), .B1(new_n321), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT73), .B(G179), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n330), .B(new_n333), .C1(new_n319), .C2(new_n320), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT84), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n333), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n321), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT84), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n330), .B1(new_n319), .B2(new_n320), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n338), .C1(new_n310), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT18), .B1(new_n309), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n289), .B1(new_n295), .B2(new_n298), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT82), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n294), .A2(new_n303), .A3(new_n276), .ZN(new_n346));
  OAI211_X1 g0146(.A(KEYINPUT16), .B(new_n287), .C1(new_n346), .C2(new_n304), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n345), .A2(new_n266), .A3(new_n347), .A4(new_n299), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n268), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT18), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n340), .A4(new_n335), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT85), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n339), .A2(G190), .ZN(new_n354));
  INV_X1    g0154(.A(G200), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n339), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n348), .A2(new_n354), .A3(new_n268), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT17), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT85), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n342), .A2(new_n361), .A3(new_n351), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n353), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n327), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n326), .A2(new_n328), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(G226), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n274), .A2(new_n275), .ZN(new_n368));
  INV_X1    g0168(.A(G1698), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G222), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n370), .C1(new_n311), .C2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(new_n212), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n320), .C1(new_n372), .C2(new_n368), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G190), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n355), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n267), .A2(G50), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n284), .A2(G150), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n209), .A2(G33), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n378), .B1(new_n201), .B2(new_n209), .C1(new_n256), .C2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G50), .ZN(new_n381));
  INV_X1    g0181(.A(new_n260), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n380), .A2(new_n266), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n376), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT10), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n387), .B(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(new_n374), .A2(G169), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n374), .A2(new_n333), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n394));
  INV_X1    g0194(.A(G232), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G1698), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n368), .B(new_n396), .C1(G226), .C2(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G97), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n320), .ZN(new_n400));
  INV_X1    g0200(.A(G238), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n327), .B1(new_n401), .B2(new_n365), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n394), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n326), .B1(new_n397), .B2(new_n398), .ZN(new_n405));
  INV_X1    g0205(.A(new_n394), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n405), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(G169), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n409));
  NAND2_X1  g0209(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n410));
  OAI211_X1 g0210(.A(G169), .B(new_n410), .C1(new_n404), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT13), .B1(new_n405), .B2(new_n402), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT78), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n407), .ZN(new_n415));
  OAI211_X1 g0215(.A(KEYINPUT78), .B(KEYINPUT13), .C1(new_n405), .C2(new_n402), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(G179), .A4(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n409), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n291), .A2(G20), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(new_n379), .B2(new_n202), .C1(new_n381), .C2(new_n281), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n259), .A2(KEYINPUT12), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n421), .B1(KEYINPUT12), .B2(new_n382), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT11), .B1(new_n420), .B2(new_n266), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n267), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n291), .B1(new_n426), .B2(KEYINPUT12), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n414), .A2(new_n415), .A3(G190), .A4(new_n416), .ZN(new_n431));
  OAI21_X1  g0231(.A(G200), .B1(new_n404), .B2(new_n407), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n428), .A4(new_n425), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n327), .B1(new_n213), .B2(new_n365), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G238), .A2(G1698), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n368), .B(new_n436), .C1(new_n395), .C2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n272), .A2(new_n205), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n320), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT74), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n435), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n333), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT15), .B(G87), .Z(new_n448));
  INV_X1    g0248(.A(new_n379), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(KEYINPUT75), .A3(new_n449), .ZN(new_n450));
  OAI221_X1 g0250(.A(new_n450), .B1(new_n209), .B2(new_n212), .C1(new_n256), .C2(new_n281), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT75), .B1(new_n448), .B2(new_n449), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n266), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n267), .A2(G77), .B1(new_n212), .B2(new_n382), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n441), .A2(new_n310), .A3(new_n443), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n443), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n442), .B1(new_n435), .B2(new_n439), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT76), .B(new_n333), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n447), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n444), .A2(G190), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n441), .A2(G200), .A3(new_n443), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n430), .A2(new_n433), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n363), .A2(new_n393), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n468), .A2(new_n209), .A3(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT23), .B1(new_n205), .B2(G20), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G116), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n469), .A2(new_n470), .B1(G20), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n209), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n368), .A2(new_n475), .A3(new_n209), .A4(G87), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n266), .B1(new_n477), .B2(KEYINPUT24), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n479), .B(new_n472), .C1(new_n474), .C2(new_n476), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n259), .A2(G20), .B1(new_n208), .B2(G33), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(G107), .A3(new_n265), .A4(new_n264), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n208), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT25), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n483), .B(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT96), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n482), .B2(new_n485), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n478), .A2(new_n480), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT97), .ZN(new_n491));
  INV_X1    g0291(.A(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n487), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT97), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n493), .B(new_n494), .C1(new_n480), .C2(new_n478), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n323), .A2(G1), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n322), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G41), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n326), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G264), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n369), .C1(new_n270), .C2(new_n271), .ZN(new_n504));
  OAI211_X1 g0304(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G294), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n320), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n326), .A2(G274), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(new_n500), .A3(KEYINPUT90), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n512));
  INV_X1    g0312(.A(G274), .ZN(new_n513));
  INV_X1    g0313(.A(new_n230), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n325), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n503), .B(new_n508), .C1(new_n510), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G169), .ZN(new_n518));
  INV_X1    g0318(.A(G179), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n517), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n491), .A2(new_n495), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G190), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  OR2_X1    g0323(.A1(new_n478), .A2(new_n480), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(G200), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n493), .A4(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT94), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n209), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT91), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT91), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n368), .A2(new_n531), .A3(new_n209), .A4(G68), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  XNOR2_X1  g0334(.A(KEYINPUT87), .B(G97), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(new_n379), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT92), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT92), .B(new_n534), .C1(new_n535), .C2(new_n379), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n540), .A3(new_n205), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n209), .B1(new_n398), .B2(new_n534), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n533), .A2(new_n538), .A3(new_n539), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n266), .ZN(new_n545));
  INV_X1    g0345(.A(new_n448), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n382), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n481), .A2(new_n265), .A3(new_n264), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G87), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT93), .ZN(new_n551));
  INV_X1    g0351(.A(G250), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n323), .B2(G1), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n208), .A2(new_n513), .A3(G45), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n326), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(G238), .A2(G1698), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n213), .B2(G1698), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n368), .B1(G33), .B2(G116), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n555), .B1(new_n558), .B2(new_n326), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n551), .B1(new_n559), .B2(new_n522), .ZN(new_n560));
  INV_X1    g0360(.A(new_n555), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n213), .A2(G1698), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G238), .B2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n471), .B1(new_n563), .B2(new_n272), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(new_n320), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(KEYINPUT93), .A3(G190), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n559), .A2(G200), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n550), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n559), .A2(new_n310), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n333), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n544), .A2(new_n266), .B1(new_n382), .B2(new_n546), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n548), .A2(new_n448), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n528), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  INV_X1    g0377(.A(new_n572), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n565), .A2(G190), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n551), .B1(new_n559), .B2(G200), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n581), .A2(new_n573), .A3(new_n549), .A4(new_n566), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(KEYINPUT94), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n552), .B1(new_n274), .B2(new_n275), .ZN(new_n585));
  NOR2_X1   g0385(.A1(KEYINPUT88), .A2(KEYINPUT4), .ZN(new_n586));
  OAI21_X1  g0386(.A(G1698), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(G244), .B1(new_n270), .B2(new_n271), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(new_n586), .B1(G33), .B2(G283), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n368), .A2(G244), .A3(new_n369), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT88), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n320), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n512), .A2(new_n515), .A3(new_n511), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT90), .B1(new_n509), .B2(new_n500), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(new_n597), .B1(new_n502), .B2(G257), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n535), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT6), .B1(new_n206), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(G20), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n284), .A2(G77), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT86), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n205), .B1(new_n294), .B2(new_n276), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n266), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n260), .A2(G97), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n548), .B2(G97), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n599), .A2(new_n310), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n595), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT89), .B(new_n320), .C1(new_n590), .C2(new_n594), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n333), .A3(new_n615), .A4(new_n598), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n516), .A2(new_n510), .B1(new_n240), .B2(new_n501), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n595), .B2(new_n613), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n355), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n609), .B(new_n611), .C1(new_n599), .C2(new_n522), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G20), .B1(G33), .B2(G283), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n535), .B2(G33), .ZN(new_n624));
  INV_X1    g0424(.A(G116), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G20), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n266), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT20), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n624), .A2(new_n266), .A3(KEYINPUT20), .A4(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n302), .A2(G116), .A3(new_n481), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n382), .A2(new_n625), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n596), .A2(new_n597), .B1(new_n502), .B2(G270), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n369), .A2(G257), .ZN(new_n637));
  NAND2_X1  g0437(.A1(G264), .A2(G1698), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n637), .B(new_n638), .C1(new_n270), .C2(new_n271), .ZN(new_n639));
  INV_X1    g0439(.A(G303), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n274), .A2(new_n640), .A3(new_n275), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n320), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT95), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT95), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n639), .A2(new_n641), .A3(new_n644), .A4(new_n320), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n635), .B(new_n310), .C1(new_n636), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n636), .A2(G179), .A3(new_n646), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n634), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n636), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G200), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n632), .A2(new_n633), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n629), .B2(new_n630), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n652), .B(new_n654), .C1(new_n522), .C2(new_n651), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(G169), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n635), .B1(new_n656), .B2(new_n654), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n650), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n622), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n467), .A2(new_n527), .A3(new_n584), .A4(new_n659), .ZN(G372));
  INV_X1    g0460(.A(new_n392), .ZN(new_n661));
  INV_X1    g0461(.A(new_n352), .ZN(new_n662));
  INV_X1    g0462(.A(new_n461), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n433), .B1(new_n418), .B2(new_n429), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n662), .B1(new_n664), .B2(new_n359), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n661), .B1(new_n665), .B2(new_n389), .ZN(new_n666));
  INV_X1    g0466(.A(new_n467), .ZN(new_n667));
  INV_X1    g0467(.A(new_n617), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n569), .A2(new_n575), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n617), .B1(new_n576), .B2(new_n583), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n579), .B(new_n671), .C1(new_n672), .C2(new_n670), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n651), .A2(KEYINPUT21), .A3(G169), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n654), .B1(new_n674), .B2(new_n648), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n310), .B1(new_n636), .B2(new_n646), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT21), .B1(new_n634), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(KEYINPUT98), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT98), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n650), .A2(new_n679), .A3(new_n657), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n520), .A2(new_n490), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n678), .A2(new_n680), .A3(KEYINPUT99), .A4(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n621), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n619), .A2(new_n615), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G200), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n686), .A2(new_n669), .A3(new_n526), .A4(new_n617), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT99), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n673), .B1(new_n682), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n666), .B1(new_n667), .B2(new_n691), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n259), .A2(new_n209), .ZN(new_n693));
  OAI21_X1  g0493(.A(G213), .B1(new_n693), .B2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n697), .A3(KEYINPUT27), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G343), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n658), .B1(new_n634), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n634), .A2(new_n701), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n678), .B2(new_n680), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n491), .A2(new_n495), .A3(new_n701), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n527), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n521), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n701), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n700), .B(KEYINPUT101), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n681), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n701), .B1(new_n650), .B2(new_n657), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n527), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n227), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n541), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n232), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n565), .A2(new_n503), .A3(new_n508), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(G179), .A3(new_n646), .A4(new_n636), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT30), .B1(new_n728), .B2(new_n599), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n565), .A2(new_n503), .A3(new_n508), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n648), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  INV_X1    g0532(.A(new_n599), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n565), .A2(new_n336), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n684), .A2(new_n517), .A3(new_n651), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n726), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n599), .A2(new_n648), .A3(KEYINPUT30), .A4(new_n730), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n701), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n714), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n659), .A2(new_n527), .A3(new_n584), .A4(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n706), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT29), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n691), .B2(new_n714), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n672), .A2(new_n670), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n579), .A2(new_n582), .A3(new_n616), .A4(new_n612), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n575), .B1(new_n751), .B2(KEYINPUT26), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT102), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n650), .A2(new_n657), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n710), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n521), .A2(KEYINPUT102), .A3(new_n657), .A4(new_n650), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n687), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(KEYINPUT29), .B(new_n700), .C1(new_n753), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n747), .B1(new_n749), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n725), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n258), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n208), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n720), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n707), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n705), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(G330), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n227), .A2(new_n368), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n227), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n227), .A2(new_n272), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT103), .Z(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n323), .B2(new_n233), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n254), .A2(G45), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n230), .B1(G20), .B2(new_n310), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n765), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n333), .A2(new_n209), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G200), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n522), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n785), .A2(G190), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT33), .B(G317), .Z(new_n790));
  OAI21_X1  g0590(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n522), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G311), .A2(new_n794), .B1(new_n797), .B2(G322), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n209), .A2(G179), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n792), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n368), .B1(new_n802), .B2(G329), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(G190), .A3(G200), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n640), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n209), .B1(new_n795), .B2(new_n519), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n800), .A2(new_n522), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n806), .A2(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n791), .A2(new_n799), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT104), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n804), .A2(new_n540), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n802), .A2(G159), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n815), .A2(KEYINPUT32), .B1(new_n205), .B2(new_n808), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(KEYINPUT32), .C2(new_n815), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n368), .B1(new_n204), .B2(new_n806), .C1(new_n793), .C2(new_n212), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G58), .B2(new_n797), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n788), .A2(G68), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n786), .A2(G50), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n812), .A2(KEYINPUT104), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n813), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n783), .B1(new_n824), .B2(new_n780), .ZN(new_n825));
  INV_X1    g0625(.A(new_n779), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n767), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n768), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n688), .A2(new_n689), .ZN(new_n830));
  INV_X1    g0630(.A(new_n687), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n682), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n579), .B1(new_n751), .B2(KEYINPUT26), .ZN(new_n833));
  INV_X1    g0633(.A(new_n672), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(KEYINPUT26), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT107), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n460), .A2(new_n456), .A3(new_n455), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT76), .B1(new_n444), .B2(new_n333), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n465), .B(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n462), .A2(new_n700), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n461), .B(new_n841), .C1(new_n837), .C2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n843), .A2(new_n845), .A3(new_n745), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n714), .B1(new_n832), .B2(new_n835), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n843), .A2(new_n845), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n747), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n765), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  INV_X1    g0654(.A(new_n765), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n780), .A2(new_n777), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n202), .B2(new_n856), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n625), .A2(new_n793), .B1(new_n796), .B2(new_n807), .ZN(new_n858));
  INV_X1    g0658(.A(G311), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n272), .B1(new_n801), .B2(new_n859), .C1(new_n806), .C2(new_n204), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n540), .A2(new_n808), .B1(new_n804), .B2(new_n205), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n786), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n862), .B1(new_n809), .B2(new_n789), .C1(new_n640), .C2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n786), .B1(new_n788), .B2(G150), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT105), .Z(new_n866));
  INV_X1    g0666(.A(G143), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n867), .B2(new_n796), .C1(new_n282), .C2(new_n793), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT34), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G132), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n368), .B1(new_n801), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G58), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n806), .A2(new_n873), .B1(new_n808), .B2(new_n291), .ZN(new_n874));
  INV_X1    g0674(.A(new_n804), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n872), .B(new_n874), .C1(G50), .C2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n868), .B2(new_n869), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n864), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT106), .ZN(new_n879));
  INV_X1    g0679(.A(new_n780), .ZN(new_n880));
  OAI221_X1 g0680(.A(new_n857), .B1(new_n778), .B2(new_n850), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n854), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(G384));
  NOR2_X1   g0683(.A1(new_n601), .A2(new_n603), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(G116), .B(new_n231), .C1(new_n885), .C2(KEYINPUT35), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n886), .A2(KEYINPUT108), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(KEYINPUT108), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n372), .B(new_n233), .C1(new_n873), .C2(new_n291), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n381), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n208), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n347), .A2(new_n266), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n307), .A2(KEYINPUT16), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n268), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n340), .A3(new_n335), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n699), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(new_n357), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n349), .A2(new_n340), .A3(new_n335), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n349), .A2(new_n699), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n357), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n900), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n907), .B1(new_n363), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n909), .A2(KEYINPUT38), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n911), .B(new_n907), .C1(new_n363), .C2(new_n908), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT39), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n349), .B(new_n699), .C1(new_n359), .C2(new_n352), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n357), .A3(new_n904), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n906), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n918), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n430), .A2(new_n701), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n662), .A2(new_n699), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n430), .A2(new_n433), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n429), .A3(new_n701), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n429), .A2(new_n701), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n430), .A2(new_n433), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n461), .A2(new_n701), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n848), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n352), .A2(KEYINPUT85), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n900), .B1(new_n936), .B2(new_n362), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n911), .B1(new_n937), .B2(new_n907), .ZN(new_n938));
  INV_X1    g0738(.A(new_n907), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n342), .A2(new_n361), .A3(new_n351), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n361), .B1(new_n342), .B2(new_n351), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n940), .A2(new_n941), .A3(new_n359), .ZN(new_n942));
  OAI211_X1 g0742(.A(KEYINPUT38), .B(new_n939), .C1(new_n942), .C2(new_n900), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n924), .B1(new_n933), .B2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n922), .A2(new_n923), .B1(new_n945), .B2(KEYINPUT109), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n467), .B(new_n759), .C1(new_n849), .C2(KEYINPUT29), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n666), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n742), .A2(new_n743), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n701), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n746), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n929), .A3(new_n850), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT40), .B1(new_n944), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n914), .A2(new_n917), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n911), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n943), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n955), .A2(new_n929), .A3(KEYINPUT40), .A4(new_n850), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n958), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n955), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n667), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n706), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n964), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n952), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n208), .B2(new_n762), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n952), .A2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n895), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT110), .Z(G367));
  INV_X1    g0773(.A(new_n241), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n781), .B1(new_n227), .B2(new_n546), .C1(new_n974), .C2(new_n773), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n975), .A2(new_n765), .ZN(new_n976));
  INV_X1    g0776(.A(new_n550), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n669), .B1(new_n977), .B2(new_n700), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n575), .A2(new_n550), .A3(new_n701), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n272), .B1(new_n801), .B2(new_n981), .C1(new_n806), .C2(new_n205), .ZN(new_n982));
  INV_X1    g0782(.A(new_n535), .ZN(new_n983));
  INV_X1    g0783(.A(new_n808), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n863), .B2(new_n859), .C1(new_n807), .C2(new_n789), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n875), .A2(G116), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n809), .B2(new_n793), .C1(new_n640), .C2(new_n796), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n212), .A2(new_n808), .B1(new_n804), .B2(new_n873), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n806), .A2(new_n291), .ZN(new_n991));
  INV_X1    g0791(.A(G137), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n368), .B1(new_n801), .B2(new_n992), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(G150), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(new_n381), .B2(new_n793), .C1(new_n995), .C2(new_n796), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n867), .A2(new_n863), .B1(new_n789), .B2(new_n282), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n986), .A2(new_n989), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT47), .Z(new_n999));
  OAI221_X1 g0799(.A(new_n976), .B1(new_n826), .B2(new_n980), .C1(new_n880), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n713), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n609), .A2(new_n611), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n714), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n617), .B(new_n1003), .C1(new_n620), .C2(new_n621), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n612), .A2(new_n714), .A3(new_n616), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT111), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT111), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT45), .B1(new_n1010), .B2(new_n717), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1004), .A2(new_n1008), .A3(new_n1005), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1008), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1013));
  OAI211_X1 g0813(.A(KEYINPUT45), .B(new_n717), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n716), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n521), .A2(new_n526), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1017), .A2(new_n1018), .B1(new_n681), .B2(new_n714), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT44), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT44), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1001), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1022), .B2(new_n1019), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n1014), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1029), .A2(new_n713), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n749), .A2(new_n759), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n527), .A2(new_n716), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n712), .B2(new_n716), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(new_n707), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n852), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n760), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n720), .B(KEYINPUT41), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n763), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT112), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1012), .A2(new_n1013), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT112), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n710), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1045), .A2(KEYINPUT113), .A3(new_n617), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT113), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1042), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1007), .A2(KEYINPUT112), .A3(new_n1009), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n521), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1047), .B1(new_n1050), .B2(new_n668), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1051), .A3(new_n745), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1022), .A2(new_n1033), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT42), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n980), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT43), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1055), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n713), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1052), .A2(new_n1059), .A3(new_n1058), .A4(new_n1054), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1064), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1041), .B(new_n1066), .C1(new_n1067), .C2(KEYINPUT114), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1064), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1056), .B(new_n1060), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1065), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT114), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1000), .B1(new_n1068), .B2(new_n1074), .ZN(G387));
  NAND3_X1  g0875(.A1(new_n709), .A2(new_n711), .A3(new_n779), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n246), .A2(G45), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1077), .A2(new_n773), .B1(new_n722), .B2(new_n769), .ZN(new_n1078));
  AOI21_X1  g0878(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n257), .A2(KEYINPUT50), .A3(new_n381), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT50), .B1(new_n257), .B2(new_n381), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n722), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1078), .A2(new_n1082), .B1(new_n205), .B2(new_n719), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n765), .B1(new_n1083), .B2(new_n782), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G159), .A2(new_n786), .B1(new_n788), .B2(new_n257), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n212), .A2(new_n804), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n272), .B(new_n1086), .C1(G150), .C2(new_n802), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n546), .A2(new_n806), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G97), .B2(new_n984), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G50), .A2(new_n797), .B1(new_n794), .B2(G68), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n368), .B1(new_n802), .B2(G326), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n806), .A2(new_n809), .B1(new_n804), .B2(new_n807), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G303), .A2(new_n794), .B1(new_n797), .B2(G317), .ZN(new_n1094));
  INV_X1    g0894(.A(G322), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1094), .B1(new_n863), .B2(new_n1095), .C1(new_n859), .C2(new_n789), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT48), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1093), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n1097), .B2(new_n1096), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT49), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1092), .B1(new_n625), .B2(new_n808), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1091), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1084), .B1(new_n1103), .B2(new_n780), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1035), .A2(new_n764), .B1(new_n1076), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1036), .A2(new_n720), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n760), .A2(new_n1035), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(G393));
  NAND2_X1  g0908(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n760), .A2(new_n1026), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n720), .A3(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n368), .B1(new_n801), .B2(new_n867), .C1(new_n540), .C2(new_n808), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n806), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(G77), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n291), .B2(new_n804), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(new_n257), .C2(new_n794), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n381), .B2(new_n789), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n786), .A2(G150), .B1(new_n797), .B2(G159), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n786), .A2(G317), .B1(new_n797), .B2(G311), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT52), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n806), .A2(new_n625), .B1(new_n804), .B2(new_n809), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n272), .B1(new_n801), .B2(new_n1095), .C1(new_n205), .C2(new_n808), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(G294), .C2(new_n794), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n640), .B2(new_n789), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1117), .A2(new_n1119), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n780), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n250), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n781), .B1(new_n227), .B2(new_n535), .C1(new_n773), .C2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n765), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1063), .B2(new_n779), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n764), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1111), .A2(KEYINPUT115), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT115), .B1(new_n1111), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G390));
  AOI21_X1  g0937(.A(new_n855), .B1(new_n256), .B2(new_n856), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n786), .A2(G283), .B1(new_n794), .B2(new_n983), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n205), .B2(new_n789), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT118), .Z(new_n1141));
  OAI221_X1 g0941(.A(new_n1114), .B1(new_n291), .B2(new_n808), .C1(new_n807), .C2(new_n801), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n814), .A2(new_n368), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G116), .C2(new_n797), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n786), .A2(G128), .B1(new_n797), .B2(G132), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT117), .Z(new_n1147));
  OR3_X1    g0947(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n995), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n804), .B2(new_n995), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n1149), .C1(new_n793), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n272), .B1(new_n802), .B2(G125), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n381), .B2(new_n808), .C1(new_n282), .C2(new_n806), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(G137), .C2(new_n788), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1141), .A2(new_n1145), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1138), .B1(new_n880), .B2(new_n1155), .C1(new_n922), .C2(new_n778), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n846), .B1(new_n832), .B2(new_n835), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n929), .B1(new_n1157), .B2(new_n931), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n923), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n913), .A2(new_n1160), .A3(new_n921), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n850), .B(new_n700), .C1(new_n753), .C2(new_n758), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(new_n932), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n961), .B(new_n1159), .C1(new_n1163), .C2(new_n930), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n747), .A2(new_n850), .A3(new_n929), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n930), .B1(new_n1162), .B2(new_n932), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n919), .A2(new_n1167), .A3(new_n923), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n920), .B1(new_n938), .B2(new_n943), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n943), .A2(new_n920), .A3(new_n960), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1168), .B1(new_n1171), .B2(new_n1160), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n955), .A2(new_n929), .A3(G330), .A4(new_n850), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1166), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1156), .B1(new_n1174), .B2(new_n763), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n965), .A2(new_n706), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n467), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n950), .A3(new_n666), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n848), .A2(new_n932), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n929), .B1(new_n747), .B2(new_n850), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT116), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1173), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(KEYINPUT116), .B(new_n929), .C1(new_n747), .C2(new_n850), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n955), .A2(G330), .A3(new_n850), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1163), .B(new_n1165), .C1(new_n1185), .C2(new_n929), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1178), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1187), .B(new_n1166), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1187), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n721), .B1(new_n1174), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1175), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(G378));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n393), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n384), .A2(new_n699), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1193), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n389), .A2(new_n392), .A3(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1194), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1196), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(G330), .B1(new_n919), .B2(new_n962), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n958), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n706), .B1(new_n961), .B2(new_n963), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n956), .B1(new_n938), .B2(new_n943), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1205), .B(new_n1201), .C1(KEYINPUT40), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n948), .A3(new_n946), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n924), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n910), .A2(new_n912), .ZN(new_n1211));
  OAI211_X1 g1011(.A(KEYINPUT109), .B(new_n1210), .C1(new_n1211), .C2(new_n1158), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n923), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1207), .B(new_n1204), .C1(new_n1214), .C2(new_n947), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(new_n1215), .A3(KEYINPUT121), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1178), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1188), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n949), .A2(new_n1219), .A3(new_n1207), .A4(new_n1204), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1209), .A2(new_n1215), .A3(KEYINPUT122), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT122), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n949), .A2(new_n1225), .A3(new_n1207), .A4(new_n1204), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n1226), .A3(new_n1218), .A4(KEYINPUT57), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n720), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1216), .A2(new_n764), .A3(new_n1220), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n856), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n765), .B1(G50), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n381), .B1(G33), .B2(G41), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n272), .B2(new_n322), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G97), .A2(new_n788), .B1(new_n786), .B2(G116), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n322), .B(new_n272), .C1(new_n801), .C2(new_n809), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n808), .A2(new_n873), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n991), .A2(new_n1236), .A3(new_n1086), .A4(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G107), .A2(new_n797), .B1(new_n794), .B2(new_n448), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1234), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n797), .A2(G128), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1113), .A2(G150), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n804), .A2(new_n1150), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n786), .A2(G125), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n789), .B2(new_n871), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G137), .C2(new_n794), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n984), .A2(G159), .ZN(new_n1252));
  AOI211_X1 g1052(.A(G33), .B(G41), .C1(new_n802), .C2(G124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1242), .B1(new_n1241), .B2(new_n1240), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1232), .B1(new_n1256), .B2(new_n780), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1202), .B2(new_n778), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT120), .Z(new_n1259));
  AND2_X1   g1059(.A1(new_n1230), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1229), .A2(new_n1260), .ZN(G375));
  AND2_X1   g1061(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1178), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1039), .A3(new_n1189), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n763), .B(KEYINPUT123), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n930), .A2(new_n777), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n765), .B1(G68), .B2(new_n1231), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n368), .B(new_n1088), .C1(G303), .C2(new_n802), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G107), .A2(new_n794), .B1(new_n797), .B2(G283), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n875), .A2(G97), .B1(new_n984), .B2(G77), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n625), .A2(new_n789), .B1(new_n863), .B2(new_n807), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G137), .A2(new_n797), .B1(new_n794), .B2(G150), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n272), .B(new_n1237), .C1(G128), .C2(new_n802), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1113), .A2(G50), .B1(new_n875), .B2(G159), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n871), .A2(new_n863), .B1(new_n789), .B2(new_n1150), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1272), .A2(new_n1273), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1268), .B1(new_n1279), .B2(new_n780), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1265), .A2(new_n1266), .B1(new_n1267), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1264), .A2(new_n1281), .ZN(G381));
  NAND3_X1  g1082(.A1(new_n1229), .A2(new_n1191), .A3(new_n1260), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1136), .B(new_n1000), .C1(new_n1068), .C2(new_n1074), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1281), .A3(new_n1264), .A4(new_n1286), .ZN(new_n1287));
  OR2_X1    g1087(.A1(new_n1283), .A2(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(new_n1287), .ZN(new_n1289));
  INV_X1    g1089(.A(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(G343), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1291), .B(KEYINPUT124), .Z(new_n1292));
  NOR2_X1   g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(G213), .B1(new_n1293), .B2(new_n1283), .ZN(G409));
  AOI21_X1  g1094(.A(new_n1038), .B1(new_n1188), .B2(new_n1217), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT125), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1295), .A2(new_n1216), .A3(new_n1298), .A4(new_n1220), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1224), .A2(new_n1226), .A3(new_n1266), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1297), .A2(new_n1258), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1191), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1260), .C1(new_n1223), .C2(new_n1228), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1291), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1262), .A2(KEYINPUT60), .A3(new_n1178), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n720), .A3(new_n1189), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT60), .B1(new_n1262), .B2(new_n1178), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1281), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n882), .ZN(new_n1311));
  OAI211_X1 g1111(.A(G384), .B(new_n1281), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(G2897), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1313), .A2(new_n1314), .A3(new_n1305), .ZN(new_n1315));
  AOI22_X1  g1115(.A1(new_n1311), .A2(new_n1312), .B1(G2897), .B2(new_n1292), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1292), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1313), .A2(new_n1320), .ZN(new_n1321));
  AOI22_X1  g1121(.A1(new_n1306), .A2(new_n1318), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(G393), .B(new_n828), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1041), .A4(new_n1066), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1136), .B1(new_n1326), .B2(new_n1000), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1323), .B1(new_n1285), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT61), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G387), .A2(G390), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1323), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1284), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1328), .A2(new_n1329), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1333), .B(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1313), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1304), .A2(new_n1305), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(new_n1320), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1322), .A2(new_n1335), .A3(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1329), .B1(new_n1319), .B2(new_n1317), .ZN(new_n1340));
  XOR2_X1   g1140(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1341));
  NAND2_X1  g1141(.A1(new_n1337), .A2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1319), .A2(KEYINPUT62), .A3(new_n1336), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1328), .A2(new_n1332), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1339), .B1(new_n1344), .B2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1191), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(new_n1313), .A3(new_n1303), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1313), .B1(new_n1348), .B2(new_n1303), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1345), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1348), .A2(new_n1303), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1336), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1354), .A2(new_n1346), .A3(new_n1349), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1352), .A2(new_n1355), .ZN(G402));
endmodule


