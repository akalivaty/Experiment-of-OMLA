//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n205), .B1(new_n209), .B2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G50), .ZN(new_n222));
  INV_X1    g0022(.A(G226), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT65), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT66), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n229), .B(new_n230), .C1(new_n226), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n220), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XOR2_X1   g0047(.A(G58), .B(G77), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  OAI211_X1 g0057(.A(G250), .B(new_n257), .C1(new_n254), .C2(new_n255), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G294), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT5), .B(G41), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G264), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  AND2_X1   g0068(.A1(G1), .A2(G13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(new_n264), .A3(new_n265), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n262), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G200), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n262), .A2(new_n267), .A3(G190), .A4(new_n272), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n216), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT90), .B1(new_n207), .B2(G107), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT23), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT23), .ZN(new_n282));
  OAI211_X1 g0082(.A(KEYINPUT90), .B(new_n282), .C1(new_n207), .C2(G107), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n207), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n281), .A2(new_n283), .B1(G116), .B2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n207), .B(G87), .C1(new_n254), .C2(new_n255), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT89), .A2(KEYINPUT22), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n288), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n292), .A2(new_n294), .A3(new_n207), .A4(G87), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT24), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT24), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n286), .A2(new_n289), .A3(new_n295), .A4(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n279), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(new_n216), .A3(new_n277), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT81), .B1(new_n304), .B2(G1), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT81), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(new_n206), .A3(G33), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT82), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n303), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT82), .B1(new_n311), .B2(new_n302), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(G107), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n301), .ZN(new_n314));
  INV_X1    g0114(.A(G107), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT25), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT25), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n301), .A2(new_n317), .A3(G107), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n276), .A2(new_n300), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n254), .A2(new_n255), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT7), .B1(new_n321), .B2(new_n207), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  NOR4_X1   g0123(.A1(new_n254), .A2(new_n255), .A3(new_n323), .A4(G20), .ZN(new_n324));
  OAI21_X1  g0124(.A(G107), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT6), .ZN(new_n326));
  AND2_X1   g0126(.A1(G97), .A2(G107), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(new_n202), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n315), .A2(KEYINPUT6), .A3(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G20), .A2(G33), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(G20), .B1(G77), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n279), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n310), .A2(G97), .A3(new_n312), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n301), .A2(G97), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT5), .A2(G41), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT5), .A2(G41), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n264), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n269), .A2(new_n270), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G257), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n272), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(G244), .B(new_n257), .C1(new_n254), .C2(new_n255), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G283), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT83), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  AOI211_X1 g0151(.A(G179), .B(new_n343), .C1(new_n261), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n261), .ZN(new_n353));
  INV_X1    g0153(.A(new_n343), .ZN(new_n354));
  AOI21_X1  g0154(.A(G169), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n336), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT84), .ZN(new_n357));
  AOI211_X1 g0157(.A(G190), .B(new_n343), .C1(new_n261), .C2(new_n351), .ZN(new_n358));
  AOI21_X1  g0158(.A(G200), .B1(new_n353), .B2(new_n354), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OR3_X1    g0160(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G190), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n353), .A2(new_n363), .A3(new_n354), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n343), .B1(new_n351), .B2(new_n261), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(G200), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT84), .A3(new_n336), .ZN(new_n367));
  AOI211_X1 g0167(.A(new_n320), .B(new_n356), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n331), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n222), .B1(new_n207), .B2(G68), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n284), .A2(new_n225), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n278), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT11), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT11), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n373), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT70), .B1(new_n207), .B2(G1), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(new_n206), .A3(G20), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G68), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n302), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT12), .B1(new_n301), .B2(G68), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n376), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G41), .ZN(new_n390));
  AOI21_X1  g0190(.A(G1), .B1(new_n390), .B2(new_n263), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n261), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G238), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  INV_X1    g0194(.A(G232), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(G1698), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n292), .B1(G33), .B2(G97), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(new_n340), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n391), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT69), .B1(new_n271), .B2(new_n391), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT13), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n395), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G226), .B2(G1698), .ZN(new_n404));
  INV_X1    g0204(.A(G97), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n321), .B1(new_n304), .B2(new_n405), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(new_n261), .B1(G238), .B2(new_n392), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n271), .A2(new_n391), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT69), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n391), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n363), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n389), .B1(new_n402), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n402), .A2(new_n418), .A3(new_n414), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n407), .A2(new_n412), .A3(KEYINPUT75), .A4(new_n413), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(G200), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n419), .A2(new_n424), .A3(G169), .A4(new_n420), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT77), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n419), .A2(G169), .A3(new_n420), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n415), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n429), .A2(KEYINPUT14), .B1(new_n402), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n423), .B1(new_n433), .B2(new_n389), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n392), .A2(G226), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n412), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n292), .A2(G222), .A3(new_n257), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n292), .A2(G223), .A3(G1698), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n225), .C2(new_n292), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n261), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(KEYINPUT71), .A3(new_n430), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT8), .B(G58), .ZN(new_n442));
  INV_X1    g0242(.A(G150), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n442), .A2(new_n284), .B1(new_n443), .B2(new_n369), .ZN(new_n444));
  NOR2_X1   g0244(.A1(G58), .A2(G68), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n207), .B1(new_n445), .B2(new_n222), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n278), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n222), .B1(new_n380), .B2(new_n382), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n303), .A2(new_n448), .B1(new_n222), .B2(new_n314), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n441), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(new_n412), .A3(new_n435), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT71), .B1(new_n453), .B2(G169), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n430), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n383), .A2(new_n225), .ZN(new_n457));
  OAI22_X1  g0257(.A1(new_n457), .A2(new_n302), .B1(G77), .B2(new_n301), .ZN(new_n458));
  INV_X1    g0258(.A(new_n442), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(new_n331), .B1(G20), .B2(G77), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT15), .B(G87), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n285), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n279), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n292), .A2(G232), .A3(new_n257), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n467), .C1(new_n315), .C2(new_n292), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n261), .ZN(new_n469));
  INV_X1    g0269(.A(new_n224), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n392), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n412), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G169), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(G179), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(G200), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n476), .B(new_n465), .C1(new_n363), .C2(new_n472), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT74), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n479), .B1(new_n452), .B2(new_n363), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n436), .A2(KEYINPUT74), .A3(G190), .A4(new_n440), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT9), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n450), .A2(KEYINPUT72), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT72), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n447), .A2(new_n486), .A3(new_n449), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(KEYINPUT9), .A3(new_n487), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT73), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n452), .B2(G200), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n482), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT10), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n492), .A2(new_n490), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT10), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n482), .A4(new_n489), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n456), .B(new_n478), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT16), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n290), .A2(new_n207), .A3(new_n291), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n323), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n291), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n384), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G58), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n384), .ZN(new_n505));
  OAI21_X1  g0305(.A(G20), .B1(new_n505), .B2(new_n445), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n331), .A2(G159), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n499), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G68), .B1(new_n322), .B2(new_n324), .ZN(new_n510));
  INV_X1    g0310(.A(new_n508), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(KEYINPUT16), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n512), .A3(new_n278), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n383), .A2(new_n302), .A3(new_n442), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n314), .B2(new_n442), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n223), .A2(G1698), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G223), .B2(G1698), .ZN(new_n518));
  INV_X1    g0318(.A(G87), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n518), .A2(new_n321), .B1(new_n304), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n261), .B1(G232), .B2(new_n392), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n521), .A2(new_n430), .A3(new_n412), .ZN(new_n522));
  AOI21_X1  g0322(.A(G169), .B1(new_n521), .B2(new_n412), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n526), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n516), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n521), .A2(new_n412), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  AND2_X1   g0333(.A1(KEYINPUT79), .A2(G190), .ZN(new_n534));
  NOR2_X1   g0334(.A1(KEYINPUT79), .A2(G190), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n521), .A2(new_n412), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n513), .A2(new_n533), .A3(new_n515), .A4(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT17), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n531), .A2(new_n540), .A3(KEYINPUT80), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n516), .A2(new_n524), .A3(new_n528), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n528), .B1(new_n516), .B2(new_n524), .ZN(new_n544));
  INV_X1    g0344(.A(new_n530), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT17), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n539), .B(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n542), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AND4_X1   g0349(.A1(new_n434), .A2(new_n498), .A3(new_n541), .A4(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT85), .ZN(new_n551));
  OR2_X1    g0351(.A1(G238), .A2(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G1698), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n552), .B(new_n554), .C1(new_n254), .C2(new_n255), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n340), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n340), .A2(G274), .A3(new_n264), .ZN(new_n558));
  INV_X1    g0358(.A(G250), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n206), .B2(G45), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n340), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n551), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n271), .A2(new_n264), .B1(new_n340), .B2(new_n560), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G238), .A2(G1698), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n553), .B2(G1698), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n566), .A2(new_n292), .B1(G33), .B2(G116), .ZN(new_n567));
  OAI211_X1 g0367(.A(KEYINPUT85), .B(new_n564), .C1(new_n567), .C2(new_n340), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n568), .A3(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT86), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n563), .A2(new_n568), .A3(new_n571), .A4(G190), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(G200), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n563), .B2(new_n568), .ZN(new_n575));
  NAND3_X1  g0375(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n207), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n203), .B2(G87), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n207), .B(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n284), .B2(new_n405), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n278), .B1(new_n314), .B2(new_n461), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n310), .A2(G87), .A3(new_n312), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n573), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n563), .A2(new_n568), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n473), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n563), .A2(new_n568), .A3(new_n430), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n310), .A2(new_n312), .A3(new_n462), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n587), .A2(new_n593), .A3(KEYINPUT87), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT87), .B1(new_n587), .B2(new_n593), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n292), .A2(G264), .A3(G1698), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n292), .A2(G257), .A3(new_n257), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT88), .B(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n292), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n261), .ZN(new_n601));
  INV_X1    g0401(.A(G270), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n272), .B1(new_n341), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n303), .A2(new_n308), .A3(G116), .ZN(new_n607));
  INV_X1    g0407(.A(G116), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n314), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT20), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT83), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n348), .B(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n207), .B1(new_n405), .B2(G33), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(G20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n278), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n611), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n617), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(KEYINPUT20), .C1(new_n613), .C2(new_n614), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n610), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n606), .B(new_n621), .C1(new_n605), .C2(new_n536), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n342), .B1(new_n290), .B2(new_n291), .ZN(new_n624));
  XOR2_X1   g0424(.A(KEYINPUT88), .B(G303), .Z(new_n625));
  AOI22_X1  g0425(.A1(new_n257), .A2(new_n624), .B1(new_n625), .B2(new_n321), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n340), .B1(new_n626), .B2(new_n597), .ZN(new_n627));
  OAI21_X1  g0427(.A(G169), .B1(new_n627), .B2(new_n603), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n618), .A2(new_n620), .ZN(new_n630));
  INV_X1    g0430(.A(new_n610), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n601), .A2(new_n604), .A3(G179), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n632), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n622), .A2(new_n629), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n262), .A2(new_n267), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n430), .A3(new_n272), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n273), .A2(new_n473), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n639), .B(new_n640), .C1(new_n300), .C2(new_n319), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n368), .A2(new_n550), .A3(new_n596), .A4(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n429), .A2(KEYINPUT14), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n431), .A2(new_n402), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n428), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n425), .A2(new_n426), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n389), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n423), .A2(new_n475), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n540), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT92), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n516), .A2(new_n524), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(new_n516), .B2(new_n524), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n525), .A2(KEYINPUT92), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n516), .A2(new_n524), .A3(new_n655), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n653), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n494), .A2(new_n497), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n456), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n641), .A2(new_n629), .A3(new_n636), .A4(new_n633), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n564), .B1(new_n567), .B2(new_n340), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n473), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n590), .A2(new_n592), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n585), .B1(G200), .B2(new_n667), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n669), .B1(new_n573), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n356), .B1(new_n362), .B2(new_n367), .ZN(new_n674));
  INV_X1    g0474(.A(new_n320), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n356), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n366), .A2(KEYINPUT84), .A3(new_n336), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT84), .B1(new_n366), .B2(new_n336), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n677), .B(new_n675), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n666), .A2(new_n671), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT91), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n671), .A2(new_n684), .A3(new_n356), .ZN(new_n685));
  INV_X1    g0485(.A(new_n669), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  AOI211_X1 g0488(.A(new_n575), .B(new_n585), .C1(new_n570), .C2(new_n572), .ZN(new_n689));
  INV_X1    g0489(.A(new_n593), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n587), .A2(new_n593), .A3(KEYINPUT87), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n356), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n687), .B1(new_n693), .B2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n683), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n550), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n665), .A2(new_n696), .ZN(G369));
  AND2_X1   g0497(.A1(new_n633), .A2(new_n636), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n629), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n621), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n637), .B2(new_n707), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n709), .B(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n705), .B1(new_n300), .B2(new_n319), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n642), .B1(new_n675), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n641), .A2(new_n705), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(G330), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n699), .A2(new_n706), .ZN(new_n717));
  OAI22_X1  g0517(.A1(new_n717), .A2(new_n713), .B1(new_n641), .B2(new_n705), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n716), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n213), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n202), .A2(new_n519), .A3(new_n608), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT95), .Z(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n218), .B2(new_n723), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT96), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n674), .A2(new_n675), .A3(new_n671), .A4(new_n666), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n691), .A2(new_n684), .A3(new_n356), .A4(new_n692), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n671), .A2(new_n356), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n669), .B1(new_n733), .B2(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .A3(new_n706), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n705), .B1(new_n683), .B2(new_n694), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n737), .B2(KEYINPUT29), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n365), .A2(new_n638), .A3(new_n563), .A4(new_n568), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n634), .ZN(new_n742));
  AND4_X1   g0542(.A1(new_n267), .A2(new_n563), .A3(new_n568), .A4(new_n262), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n635), .A2(new_n743), .A3(KEYINPUT30), .A4(new_n365), .ZN(new_n744));
  INV_X1    g0544(.A(new_n365), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n667), .A2(new_n430), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n746), .A3(new_n605), .A4(new_n273), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n742), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n705), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT31), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n596), .A2(new_n368), .A3(new_n643), .A4(new_n706), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n739), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n738), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n730), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n211), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n206), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n722), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n473), .A2(KEYINPUT98), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n207), .B1(KEYINPUT98), .B2(new_n473), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n216), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n213), .A2(new_n321), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT97), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n219), .A2(new_n263), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n773), .B(new_n774), .C1(new_n249), .C2(new_n263), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n721), .A2(new_n321), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G355), .B1(new_n608), .B2(new_n721), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n771), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n574), .A2(G179), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n780), .A2(new_n207), .A3(new_n363), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n292), .B1(new_n782), .B2(new_n519), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n207), .A2(new_n430), .A3(new_n574), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G190), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(G68), .B2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n207), .A2(new_n430), .A3(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n537), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n785), .A2(new_n536), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(G58), .B1(new_n791), .B2(G50), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n363), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n207), .B1(new_n795), .B2(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(G77), .B1(G97), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n363), .A2(G20), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT99), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n780), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G107), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n787), .A2(new_n792), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n801), .A2(G179), .A3(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G159), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n794), .A2(G311), .B1(G294), .B2(new_n797), .ZN(new_n808));
  INV_X1    g0608(.A(G322), .ZN(new_n809));
  INV_X1    g0609(.A(G326), .ZN(new_n810));
  INV_X1    g0610(.A(new_n791), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(new_n809), .B2(new_n789), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n805), .A2(G329), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n802), .A2(G283), .ZN(new_n814));
  INV_X1    g0614(.A(G317), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n786), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n292), .B1(new_n781), .B2(G303), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n813), .A2(new_n814), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n804), .A2(new_n807), .B1(new_n812), .B2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n761), .B(new_n778), .C1(new_n765), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT100), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n709), .B2(new_n770), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n711), .A2(G330), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n761), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n711), .A2(G330), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G396));
  OR2_X1    g0628(.A1(new_n475), .A2(new_n705), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n477), .B1(new_n465), .B2(new_n706), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n475), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n737), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n760), .B1(new_n834), .B2(new_n753), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n753), .B2(new_n834), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n766), .A2(new_n768), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n760), .B1(G77), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n791), .A2(G137), .B1(new_n794), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  INV_X1    g0640(.A(new_n786), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n789), .C1(new_n443), .C2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT101), .Z(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(KEYINPUT34), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n292), .B1(new_n504), .B2(new_n796), .C1(new_n782), .C2(new_n222), .ZN(new_n846));
  INV_X1    g0646(.A(new_n802), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n384), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n846), .B(new_n848), .C1(G132), .C2(new_n805), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n844), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n321), .B1(new_n405), .B2(new_n796), .C1(new_n782), .C2(new_n315), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G87), .B2(new_n802), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n790), .A2(G294), .B1(new_n791), .B2(G303), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n786), .A2(G283), .B1(new_n794), .B2(G116), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n805), .A2(G311), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n838), .B1(new_n857), .B2(new_n765), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n768), .B2(new_n833), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n836), .A2(KEYINPUT102), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT102), .B1(new_n836), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  NAND2_X1  g0663(.A1(new_n217), .A2(G116), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n330), .B2(KEYINPUT35), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n330), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OAI21_X1  g0667(.A(G77), .B1(new_n504), .B2(new_n384), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n868), .A2(new_n218), .B1(G50), .B2(new_n384), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n211), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT103), .Z(new_n872));
  NAND2_X1  g0672(.A1(new_n389), .A2(new_n705), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n649), .A2(new_n422), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n389), .B(new_n705), .C1(new_n433), .C2(new_n423), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n737), .A2(new_n833), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n877), .B1(new_n878), .B2(new_n829), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n703), .B1(new_n513), .B2(new_n515), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n546), .B2(new_n548), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n525), .A2(new_n882), .A3(new_n539), .ZN(new_n883));
  INV_X1    g0683(.A(new_n703), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT104), .B1(new_n516), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n886), .B(new_n703), .C1(new_n513), .C2(new_n515), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n516), .A2(new_n884), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n525), .A2(new_n890), .A3(new_n539), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n881), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n531), .B2(new_n540), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n883), .A2(new_n888), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n879), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n539), .B1(new_n656), .B2(new_n657), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n880), .B(KEYINPUT104), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n658), .A2(new_n661), .A3(new_n540), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n889), .A2(new_n904), .B1(new_n905), .B2(new_n903), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n901), .B(new_n894), .C1(new_n906), .C2(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n896), .A2(new_n897), .A3(new_n895), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n881), .B2(new_n893), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT39), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n910), .A3(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n889), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n905), .A2(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n914), .B2(new_n895), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n916), .A3(new_n901), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n649), .A2(new_n705), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n662), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n703), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n900), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n550), .B(new_n736), .C1(new_n737), .C2(KEYINPUT29), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(new_n665), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  INV_X1    g0725(.A(KEYINPUT31), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT106), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n749), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n926), .A4(new_n705), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n832), .B1(new_n751), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n876), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT40), .B1(new_n932), .B2(new_n915), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT40), .B1(new_n894), .B2(new_n898), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n876), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n751), .A2(new_n930), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n550), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n739), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n925), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n206), .B2(new_n757), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n925), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n872), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n674), .B1(new_n336), .B2(new_n706), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n356), .A2(new_n705), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n717), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n715), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n677), .B1(new_n945), .B2(new_n641), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(KEYINPUT42), .B1(new_n706), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT42), .B2(new_n949), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n585), .A2(new_n705), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n686), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n671), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n953), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g0759(.A(new_n947), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n716), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n722), .B(KEYINPUT41), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n948), .B(new_n715), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n825), .B(new_n964), .Z(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n755), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT107), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n825), .B(new_n964), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n754), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n716), .A2(KEYINPUT108), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n960), .A2(new_n972), .A3(new_n718), .ZN(new_n973));
  AOI21_X1  g0773(.A(KEYINPUT45), .B1(new_n719), .B2(new_n947), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n716), .A2(KEYINPUT108), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT44), .B1(new_n960), .B2(new_n718), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n719), .A2(new_n947), .A3(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n971), .A2(new_n975), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n975), .A2(new_n980), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(KEYINPUT108), .A3(new_n716), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT109), .B1(new_n970), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n981), .A2(new_n983), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT109), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n986), .A2(new_n966), .A3(new_n987), .A4(new_n969), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n963), .B1(new_n989), .B2(new_n755), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n962), .B1(new_n990), .B2(new_n759), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n773), .A2(new_n244), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n771), .B1(new_n721), .B2(new_n462), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n761), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n782), .B2(new_n608), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(G294), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n997), .C1(new_n998), .C2(new_n841), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT110), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n791), .A2(G311), .B1(new_n794), .B2(G283), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n315), .B2(new_n796), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n292), .B1(new_n790), .B2(new_n625), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n805), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n847), .B2(new_n405), .C1(new_n1004), .C2(new_n815), .ZN(new_n1005));
  NOR3_X1   g0805(.A1(new_n1000), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT111), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n796), .A2(new_n384), .ZN(new_n1008));
  INV_X1    g0808(.A(G159), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n840), .A2(new_n811), .B1(new_n841), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G50), .C2(new_n794), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n802), .A2(G77), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n805), .A2(G137), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n292), .B1(new_n782), .B2(new_n504), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n790), .B2(G150), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n994), .B1(new_n1018), .B2(new_n766), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n769), .B2(new_n956), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n991), .A2(new_n1021), .ZN(G387));
  OAI211_X1 g0822(.A(new_n970), .B(new_n722), .C1(new_n755), .C2(new_n965), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n773), .B1(new_n241), .B2(new_n263), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n776), .A2(new_n725), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n442), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT50), .B1(new_n442), .B2(G50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n726), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(new_n315), .B2(new_n721), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n760), .B1(new_n1031), .B2(new_n771), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT113), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n292), .B1(new_n384), .B2(new_n793), .C1(new_n782), .C2(new_n225), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G97), .B2(new_n802), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n791), .A2(G159), .B1(new_n797), .B2(new_n462), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n790), .A2(G50), .B1(new_n786), .B2(new_n459), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n805), .A2(G150), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n292), .B1(new_n805), .B2(G326), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G322), .A2(new_n791), .B1(new_n786), .B2(G311), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(KEYINPUT114), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n790), .A2(G317), .B1(new_n625), .B2(new_n794), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n781), .A2(G294), .B1(G283), .B2(new_n797), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT115), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1040), .B1(new_n608), .B2(new_n847), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1051), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1039), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1033), .B1(new_n1056), .B2(new_n765), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT116), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n715), .B2(new_n770), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1023), .B1(new_n758), .B2(new_n968), .C1(new_n1059), .C2(new_n1061), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n773), .A2(new_n252), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n771), .B1(new_n721), .B2(G97), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n761), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n790), .A2(G311), .B1(new_n791), .B2(G317), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT52), .Z(new_n1067));
  OAI21_X1  g0867(.A(new_n803), .B1(new_n1004), .B2(new_n809), .ZN(new_n1068));
  INV_X1    g0868(.A(G283), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n321), .B1(new_n608), .B2(new_n796), .C1(new_n782), .C2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n841), .A2(new_n599), .B1(new_n998), .B2(new_n793), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1004), .A2(new_n840), .B1(new_n847), .B2(new_n519), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n292), .B1(new_n782), .B2(new_n384), .C1(new_n841), .C2(new_n222), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n793), .A2(new_n442), .B1(new_n225), .B2(new_n796), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n811), .A2(new_n443), .B1(new_n1009), .B2(new_n789), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1067), .A2(new_n1072), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1065), .B1(new_n766), .B2(new_n1079), .C1(new_n947), .C2(new_n770), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n984), .B2(new_n758), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n723), .B1(new_n970), .B2(new_n984), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1081), .B1(new_n989), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(new_n918), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n829), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n737), .B2(new_n833), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1087), .B2(new_n877), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n911), .A2(new_n917), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n735), .A2(new_n706), .A3(new_n831), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n829), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n876), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n905), .A2(new_n903), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n659), .A2(new_n660), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n888), .A3(new_n539), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1096), .A2(KEYINPUT37), .B1(new_n888), .B2(new_n883), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n895), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n918), .B1(new_n1098), .B2(new_n894), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1093), .A2(KEYINPUT117), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT117), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1091), .A2(new_n829), .B1(new_n874), .B2(new_n875), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT38), .B1(new_n912), .B2(new_n913), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1085), .B1(new_n1103), .B2(new_n908), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n752), .A2(new_n833), .A3(new_n876), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1090), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1089), .A2(new_n1088), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n931), .A2(G330), .A3(new_n876), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n550), .A2(G330), .A3(new_n937), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n923), .A2(new_n665), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n750), .A2(new_n751), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(G330), .A3(new_n833), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n877), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1110), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1087), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n931), .A2(G330), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n877), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1092), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n1107), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1113), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1111), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1108), .B(new_n1124), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n722), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1108), .B(new_n759), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1089), .A2(new_n767), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n760), .B1(new_n459), .B2(new_n837), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n781), .A2(G150), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT53), .Z(new_n1133));
  AOI22_X1  g0933(.A1(new_n790), .A2(G132), .B1(G159), .B2(new_n797), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n321), .B1(new_n794), .B2(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(G128), .A2(new_n791), .B1(new_n786), .B2(G137), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n805), .A2(G125), .B1(new_n802), .B2(G50), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1135), .A2(new_n1138), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n848), .B1(G294), .B2(new_n805), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT118), .Z(new_n1143));
  OAI221_X1 g0943(.A(new_n321), .B1(new_n225), .B2(new_n796), .C1(new_n782), .C2(new_n519), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n841), .A2(new_n315), .B1(new_n793), .B2(new_n405), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n811), .A2(new_n1069), .B1(new_n608), .B2(new_n789), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1141), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1131), .B1(new_n1148), .B2(new_n765), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1130), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1129), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1128), .A2(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(new_n456), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n664), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n703), .B1(new_n484), .B2(new_n487), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n664), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1158), .B1(new_n664), .B2(new_n1154), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n456), .B(new_n1156), .C1(new_n494), .C2(new_n497), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1162), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n936), .B2(G330), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n739), .B(new_n1166), .C1(new_n933), .C2(new_n935), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n922), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n931), .B(new_n876), .C1(new_n1103), .C2(new_n908), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n876), .A2(new_n937), .A3(new_n833), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(KEYINPUT40), .A2(new_n1171), .B1(new_n1172), .B2(new_n934), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1166), .B1(new_n1173), .B2(new_n739), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT40), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1098), .A2(new_n894), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n935), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n1167), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n879), .A2(new_n899), .B1(new_n920), .B2(new_n703), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1174), .A2(new_n919), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1166), .A2(new_n767), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n760), .B1(G50), .B2(new_n837), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n791), .A2(G116), .B1(new_n794), .B2(new_n462), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n405), .B2(new_n841), .C1(new_n315), .C2(new_n789), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n847), .A2(new_n504), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n782), .A2(new_n225), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n321), .A2(new_n390), .ZN(new_n1189));
  OR4_X1    g0989(.A1(new_n1008), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1186), .B(new_n1190), .C1(G283), .C2(new_n805), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1193));
  AOI21_X1  g0993(.A(G50), .B1(new_n304), .B2(new_n390), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1192), .A2(new_n1193), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n790), .A2(G128), .B1(G137), .B2(new_n794), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G125), .A2(new_n791), .B1(new_n786), .B2(G132), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n781), .A2(new_n1137), .B1(G150), .B2(new_n797), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT59), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT120), .B(G124), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n805), .C2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(new_n1009), .C2(new_n847), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1195), .B1(new_n1200), .B2(new_n1204), .C1(new_n1193), .C2(new_n1192), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1184), .B1(new_n1205), .B2(new_n765), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1182), .A2(new_n759), .B1(new_n1183), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1113), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1127), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n1170), .B2(new_n1181), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n722), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1182), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(G375));
  INV_X1    g1015(.A(new_n963), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1119), .A2(new_n1113), .A3(new_n1123), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1125), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1122), .A2(new_n1107), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1219), .A2(new_n1121), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n877), .A2(new_n767), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n760), .B1(G68), .B2(new_n837), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n321), .B1(new_n461), .B2(new_n796), .C1(new_n782), .C2(new_n405), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G77), .B2(new_n802), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n791), .A2(G294), .B1(new_n794), .B2(G107), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n790), .A2(G283), .B1(new_n786), .B2(G116), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n805), .A2(G303), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1187), .A2(new_n321), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT122), .Z(new_n1232));
  AOI22_X1  g1032(.A1(new_n790), .A2(G137), .B1(G159), .B2(new_n781), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n805), .A2(G128), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n786), .A2(new_n1137), .B1(new_n794), .B2(G150), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n791), .A2(G132), .B1(new_n797), .B2(G50), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1230), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1224), .B1(new_n1238), .B2(new_n765), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1221), .A2(new_n759), .B1(new_n1222), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1218), .A2(new_n1240), .ZN(G381));
  OR4_X1    g1041(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1242), .A2(G387), .A3(G390), .A4(G378), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n1207), .C1(new_n1214), .C2(new_n1213), .ZN(G407));
  AOI21_X1  g1044(.A(new_n723), .B1(new_n1111), .B2(new_n1125), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1151), .B1(new_n1245), .B2(new_n1127), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n704), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  XNOR2_X1  g1048(.A(G393), .B(G396), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n991), .A2(G390), .A3(new_n1021), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G390), .B1(new_n991), .B2(new_n1021), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1083), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1249), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1255), .A3(new_n1250), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1253), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1207), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1209), .A2(new_n1216), .A3(new_n1182), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1207), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1246), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n704), .A2(G213), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT60), .B1(new_n1220), .B2(new_n1113), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n723), .B1(new_n1267), .B2(new_n1217), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1220), .A2(KEYINPUT60), .A3(new_n1113), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1266), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1217), .B1(new_n1124), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(new_n722), .A3(new_n1269), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1273), .A2(KEYINPUT124), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1240), .B1(new_n1270), .B2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n862), .A2(KEYINPUT125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n862), .A2(KEYINPUT125), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1273), .B(KEYINPUT124), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1279), .A2(new_n862), .A3(KEYINPUT125), .A4(new_n1240), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1281), .A2(KEYINPUT63), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1258), .B1(new_n1265), .B2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n704), .A2(G213), .A3(G2897), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1281), .B(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT123), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1259), .A2(new_n1286), .A3(new_n1262), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1264), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1286), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1288), .A2(new_n1292), .A3(new_n1289), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1293), .A2(KEYINPUT63), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1283), .A2(new_n1291), .A3(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1285), .B2(new_n1265), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1293), .B2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1289), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1300), .A2(new_n1264), .A3(new_n1281), .A4(new_n1287), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(KEYINPUT127), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1265), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1297), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1295), .B1(new_n1306), .B2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(G375), .A2(new_n1246), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1259), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1292), .B(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1307), .B(new_n1311), .ZN(G402));
endmodule


