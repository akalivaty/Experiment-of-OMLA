//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT0), .A2(G128), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G137), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n195), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n189), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n187), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(G128), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n197), .A2(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n199), .A2(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(G131), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND4_X1   g029(.A1(new_n203), .A2(new_n210), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT2), .A2(G113), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(KEYINPUT2), .B2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT2), .A2(G113), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(KEYINPUT2), .A3(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n217), .A3(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n206), .A2(new_n216), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n231), .B2(KEYINPUT28), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n228), .A2(new_n217), .A3(new_n223), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n223), .B1(new_n228), .B2(new_n217), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n205), .A2(new_n203), .ZN(new_n236));
  INV_X1    g050(.A(new_n195), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n210), .A2(new_n203), .A3(new_n215), .A4(new_n212), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT28), .B1(new_n231), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n235), .A3(new_n239), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT65), .A2(G953), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(G210), .A3(new_n249), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT27), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT65), .A2(G953), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT65), .A2(G953), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n255), .A2(new_n256), .A3(G210), .A4(new_n249), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n252), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n252), .B2(new_n257), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n232), .A2(new_n241), .A3(new_n245), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n259), .A2(new_n260), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT30), .B1(new_n206), .B2(new_n216), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n238), .A2(new_n266), .A3(new_n239), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n235), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n268), .B2(new_n231), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n262), .A2(new_n263), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n264), .A2(new_n263), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n232), .A2(new_n241), .A3(new_n245), .A4(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n230), .B1(new_n206), .B2(new_n216), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n244), .B1(new_n276), .B2(new_n242), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n278), .A2(KEYINPUT69), .A3(new_n232), .A4(new_n271), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n270), .A2(new_n274), .A3(new_n279), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G472), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(KEYINPUT70), .A3(G472), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NOR2_X1   g101(.A1(G472), .A2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n232), .A2(new_n241), .A3(new_n245), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n264), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n206), .A2(new_n216), .A3(KEYINPUT30), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n266), .B1(new_n238), .B2(new_n239), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n230), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n242), .A2(new_n261), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n298), .B1(new_n268), .B2(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n289), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT67), .B(KEYINPUT32), .Z(new_n302));
  OAI21_X1  g116(.A(new_n287), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n302), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n290), .A2(new_n264), .B1(new_n297), .B2(new_n299), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT68), .B(new_n304), .C1(new_n305), .C2(new_n289), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT71), .B1(new_n301), .B2(KEYINPUT32), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n286), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n314));
  NOR2_X1   g128(.A1(G475), .A2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(G113), .B(G122), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT85), .B(G104), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT72), .B(G125), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G125), .A2(G140), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n319), .B2(G140), .ZN(new_n324));
  OAI211_X1 g138(.A(G146), .B(new_n322), .C1(new_n324), .C2(new_n320), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT72), .A2(G125), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT72), .A2(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(G140), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT19), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G125), .B(G140), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT19), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n187), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n325), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n248), .A2(G214), .A3(new_n249), .A4(new_n250), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n189), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n255), .A2(G143), .A3(G214), .A4(new_n249), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n201), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT18), .A2(G131), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(KEYINPUT82), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n338), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n328), .A2(G146), .A3(new_n329), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n331), .A2(new_n187), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND4_X1   g165(.A1(KEYINPUT83), .A2(new_n346), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n339), .A2(new_n345), .B1(new_n350), .B2(new_n349), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT83), .B1(new_n353), .B2(new_n348), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n343), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT84), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n336), .B(G143), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n348), .B(new_n351), .C1(new_n358), .C2(new_n344), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n353), .A2(KEYINPUT83), .A3(new_n348), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT84), .A3(new_n343), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n318), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n340), .A2(new_n366), .A3(new_n341), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT86), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n340), .A2(new_n369), .A3(new_n366), .A4(new_n341), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n320), .B1(new_n328), .B2(new_n329), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n326), .A2(new_n327), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n372), .A2(KEYINPUT16), .A3(G140), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n187), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n325), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n366), .B(new_n201), .C1(new_n337), .C2(new_n338), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n370), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n318), .A3(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n314), .B(new_n315), .C1(new_n365), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n315), .ZN(new_n382));
  INV_X1    g196(.A(new_n318), .ZN(new_n383));
  AOI221_X4 g197(.A(new_n356), .B1(new_n335), .B2(new_n342), .C1(new_n361), .C2(new_n362), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT84), .B1(new_n363), .B2(new_n343), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n386), .B2(new_n379), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n388));
  OAI21_X1  g202(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n318), .A2(KEYINPUT87), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(new_n363), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n280), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n378), .B2(new_n363), .ZN(new_n393));
  OAI21_X1  g207(.A(G475), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(new_n396), .A3(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n189), .B2(G128), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n211), .A2(KEYINPUT88), .A3(G143), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n189), .A2(G128), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n197), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n399), .A2(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT13), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n404), .A2(new_n405), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n211), .A2(G143), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(KEYINPUT89), .B1(KEYINPUT13), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n211), .B2(G143), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n406), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n410), .B1(new_n419), .B2(G134), .ZN(new_n420));
  INV_X1    g234(.A(G116), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(G122), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(G107), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n399), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n424), .A2(new_n399), .ZN(new_n426));
  INV_X1    g240(.A(new_n408), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n197), .B1(new_n406), .B2(new_n407), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n398), .B1(new_n420), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n197), .B1(new_n414), .B2(new_n418), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n429), .B(new_n397), .C1(new_n432), .C2(new_n410), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n280), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n437), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n434), .B2(new_n280), .ZN(new_n440));
  INV_X1    g254(.A(G952), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  INV_X1    g256(.A(G234), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n249), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n280), .B(new_n255), .C1(G234), .C2(G237), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(G898), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n438), .A2(new_n440), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n389), .A2(new_n394), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n395), .B2(G902), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(G110), .B(G140), .Z(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT74), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n255), .A2(G227), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n236), .ZN(new_n458));
  INV_X1    g272(.A(G104), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT3), .B1(new_n459), .B2(G107), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n401), .A3(G104), .ZN(new_n462));
  INV_X1    g276(.A(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(G107), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n459), .A2(G107), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n401), .A2(G104), .ZN(new_n467));
  OAI21_X1  g281(.A(G101), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n210), .A2(new_n465), .A3(new_n468), .A4(new_n212), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT75), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT10), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT10), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT4), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(G101), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n476), .A2(G101), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n237), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n458), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT10), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT10), .B1(new_n469), .B2(new_n470), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n458), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n457), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(KEYINPUT76), .A3(new_n456), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n210), .A2(new_n212), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n465), .A2(new_n468), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n469), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT12), .B1(new_n492), .B2(new_n236), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(KEYINPUT12), .A3(new_n236), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n488), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT76), .B1(new_n485), .B2(new_n456), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n487), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n280), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n280), .ZN(new_n502));
  INV_X1    g316(.A(new_n482), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n485), .A2(new_n456), .ZN(new_n504));
  INV_X1    g318(.A(new_n495), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n485), .B1(new_n505), .B2(new_n493), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n503), .A2(new_n504), .B1(new_n506), .B2(new_n457), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(G469), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n452), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  INV_X1    g324(.A(G119), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G116), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n421), .A2(G119), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT5), .ZN(new_n514));
  OR3_X1    g328(.A1(new_n421), .A2(KEYINPUT5), .A3(G119), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(G113), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n229), .A3(new_n465), .A4(new_n468), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n478), .B1(new_n233), .B2(new_n234), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n479), .A2(new_n480), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n510), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n210), .A2(new_n212), .A3(new_n372), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n192), .B(new_n319), .C1(new_n193), .C2(new_n194), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n247), .A2(G224), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT79), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n521), .A2(KEYINPUT7), .A3(new_n526), .A4(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n510), .B(KEYINPUT8), .ZN(new_n531));
  AND4_X1   g345(.A1(new_n229), .A2(new_n516), .A3(new_n465), .A4(new_n468), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n516), .A2(new_n229), .B1(new_n465), .B2(new_n468), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n520), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n280), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT80), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n538));
  INV_X1    g352(.A(new_n510), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT78), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n520), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n538), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n523), .B(new_n526), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT80), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n535), .A2(new_n548), .A3(new_n280), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n537), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G210), .B1(G237), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n537), .A2(new_n547), .A3(new_n551), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n556), .B(KEYINPUT77), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n509), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n450), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n511), .A2(G128), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n511), .A2(G128), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(KEYINPUT23), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(G110), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n325), .B(new_n350), .C1(new_n565), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(G110), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT73), .B1(new_n375), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT73), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n575), .B(new_n572), .C1(new_n374), .C2(new_n325), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n569), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n255), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n569), .B(new_n580), .C1(new_n574), .C2(new_n576), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n280), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n582), .A2(KEYINPUT25), .A3(new_n280), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n396), .B1(G234), .B2(new_n280), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n583), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(G902), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n313), .A2(new_n560), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT90), .B(G101), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT91), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n555), .B2(new_n556), .ZN(new_n600));
  INV_X1    g414(.A(new_n556), .ZN(new_n601));
  AOI211_X1 g415(.A(KEYINPUT91), .B(new_n601), .C1(new_n553), .C2(new_n554), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n448), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n436), .A2(G902), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT33), .B1(new_n434), .B2(KEYINPUT92), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n607), .B(new_n608), .C1(new_n431), .C2(new_n433), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n605), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n435), .A2(new_n436), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n605), .ZN(new_n614));
  INV_X1    g428(.A(new_n433), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n211), .A2(KEYINPUT88), .A3(G143), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT88), .B1(new_n211), .B2(G143), .ZN(new_n617));
  OAI211_X1 g431(.A(KEYINPUT89), .B(new_n415), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n621));
  OAI21_X1  g435(.A(G134), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n410), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n397), .B1(new_n624), .B2(new_n429), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT92), .B1(new_n615), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n608), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n434), .A2(KEYINPUT92), .A3(KEYINPUT33), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n614), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n612), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT93), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n389), .A2(new_n394), .B1(new_n613), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n603), .A2(new_n604), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n297), .A2(new_n299), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n261), .B1(new_n278), .B2(new_n232), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n280), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n301), .B1(new_n636), .B2(G472), .ZN(new_n637));
  AND4_X1   g451(.A1(new_n590), .A2(new_n509), .A3(new_n637), .A4(new_n594), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NAND3_X1  g455(.A1(new_n555), .A2(new_n599), .A3(new_n556), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n438), .A2(new_n440), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n387), .A2(new_n388), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n315), .B1(new_n365), .B2(new_n380), .ZN(new_n645));
  INV_X1    g459(.A(new_n388), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n535), .A2(new_n548), .A3(new_n280), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n548), .B1(new_n535), .B2(new_n280), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n551), .B1(new_n651), .B2(new_n547), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n551), .A2(new_n537), .A3(new_n547), .A4(new_n549), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n556), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT91), .ZN(new_n655));
  INV_X1    g469(.A(new_n394), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n448), .B(KEYINPUT94), .Z(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n642), .A2(new_n648), .A3(new_n655), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n638), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  OR2_X1    g477(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n577), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n577), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n665), .A2(new_n593), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n590), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n560), .A2(new_n637), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI21_X1  g486(.A(new_n667), .B1(new_n588), .B2(new_n589), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n600), .A2(new_n602), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n445), .B1(new_n446), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n394), .A2(new_n677), .ZN(new_n678));
  AOI211_X1 g492(.A(new_n643), .B(new_n678), .C1(new_n644), .C2(new_n647), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n313), .A2(new_n674), .A3(new_n509), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  AOI21_X1  g495(.A(new_n643), .B1(new_n389), .B2(new_n394), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n556), .A3(new_n673), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT96), .Z(new_n684));
  INV_X1    g498(.A(KEYINPUT95), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n303), .B(new_n306), .C1(new_n686), .C2(new_n309), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n261), .B1(new_n268), .B2(new_n231), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n264), .A2(new_n276), .A3(new_n242), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n280), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n685), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n308), .A2(new_n312), .A3(KEYINPUT95), .A4(new_n692), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n555), .B(KEYINPUT38), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n676), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n509), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT40), .Z(new_n700));
  AND4_X1   g514(.A1(new_n684), .A2(new_n696), .A3(new_n697), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT97), .B(G143), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G45));
  AOI221_X4 g517(.A(new_n676), .B1(new_n631), .B2(new_n613), .C1(new_n389), .C2(new_n394), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n313), .A2(new_n704), .A3(new_n674), .A4(new_n509), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n595), .ZN(new_n707));
  INV_X1    g521(.A(new_n687), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(new_n286), .ZN(new_n709));
  INV_X1    g523(.A(new_n501), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n500), .B1(new_n499), .B2(new_n280), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n452), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(new_n633), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND3_X1  g529(.A1(new_n709), .A2(new_n660), .A3(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AND3_X1   g531(.A1(new_n389), .A2(new_n394), .A3(new_n449), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n281), .A2(KEYINPUT70), .A3(G472), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT70), .B1(new_n281), .B2(G472), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n718), .B1(new_n721), .B2(new_n687), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n655), .A2(new_n669), .A3(new_n712), .A4(new_n642), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT98), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n642), .A2(new_n655), .A3(new_n669), .A4(new_n712), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT98), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n726), .A3(new_n313), .A4(new_n718), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  INV_X1    g543(.A(KEYINPUT99), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n278), .A2(new_n730), .A3(new_n232), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n261), .B1(new_n290), .B2(KEYINPUT99), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n634), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(G472), .ZN(new_n734));
  AOI21_X1  g548(.A(G902), .B1(new_n291), .B2(new_n300), .ZN(new_n735));
  OAI22_X1  g549(.A1(new_n733), .A2(new_n289), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n595), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT100), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n595), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n603), .A2(new_n682), .ZN(new_n743));
  INV_X1    g557(.A(new_n712), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n658), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NOR2_X1   g561(.A1(new_n673), .A2(new_n736), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n704), .A2(new_n603), .A3(new_n712), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT32), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n305), .B2(new_n289), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n305), .A2(KEYINPUT103), .A3(new_n751), .A4(new_n289), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n301), .B2(KEYINPUT32), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n595), .B1(new_n721), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n758));
  OAI221_X1 g572(.A(new_n752), .B1(new_n753), .B2(new_n755), .C1(new_n719), .C2(new_n720), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n760), .A3(new_n595), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n677), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT102), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n553), .A2(KEYINPUT102), .A3(new_n554), .A4(new_n556), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n503), .A2(new_n504), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n506), .A2(new_n457), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT101), .B1(new_n770), .B2(new_n500), .ZN(new_n771));
  INV_X1    g585(.A(new_n502), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT101), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n507), .A2(new_n773), .A3(G469), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n771), .A2(new_n501), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n766), .A2(new_n451), .A3(new_n767), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n763), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n776), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n704), .A2(new_n778), .A3(new_n313), .A4(new_n595), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n762), .A2(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n201), .ZN(G33));
  NAND3_X1  g596(.A1(new_n709), .A2(new_n679), .A3(new_n778), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n766), .A2(new_n767), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n507), .A2(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n507), .A2(KEYINPUT45), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(G469), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT46), .B1(new_n788), .B2(new_n772), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(KEYINPUT46), .A3(new_n772), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n501), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n789), .B1(new_n791), .B2(KEYINPUT105), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT105), .B2(new_n791), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n451), .A3(new_n698), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n631), .A2(new_n613), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n389), .A3(new_n394), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT106), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT107), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT107), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n673), .A2(new_n637), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n785), .B(new_n794), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n793), .A2(new_n809), .A3(new_n451), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n793), .B2(new_n451), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT109), .B(KEYINPUT47), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n812), .ZN(new_n814));
  NAND2_X1  g628(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n815));
  OR2_X1    g629(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n313), .A2(new_n595), .A3(new_n785), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n704), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND3_X1  g635(.A1(new_n595), .A2(new_n558), .A3(new_n451), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n697), .A3(new_n796), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n710), .A2(new_n711), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT49), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n823), .A2(new_n694), .A3(new_n695), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n800), .B2(new_n444), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n798), .B(KEYINPUT43), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n445), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n829), .A2(new_n831), .B1(new_n741), .B2(new_n739), .ZN(new_n832));
  INV_X1    g646(.A(new_n785), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n710), .A2(new_n711), .A3(new_n451), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n813), .A2(new_n817), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n832), .A2(KEYINPUT115), .A3(new_n833), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n833), .A2(new_n712), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n829), .B2(new_n831), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n696), .A2(new_n707), .A3(new_n842), .A4(new_n444), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n656), .B(new_n795), .C1(new_n647), .C2(new_n381), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n843), .A2(new_n748), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n697), .A2(new_n744), .A3(new_n556), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n832), .A2(KEYINPUT50), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT50), .B1(new_n832), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n827), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n853));
  INV_X1    g667(.A(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n855), .A3(KEYINPUT51), .A4(new_n846), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n832), .A2(new_n603), .A3(new_n712), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n844), .A2(new_n632), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n442), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n843), .ZN(new_n860));
  INV_X1    g674(.A(new_n762), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n860), .A2(KEYINPUT48), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT48), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n856), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n709), .B(new_n712), .C1(new_n633), .C2(new_n660), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n728), .A2(new_n746), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n632), .A2(new_n748), .A3(new_n677), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT111), .B1(new_n869), .B2(new_n776), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT111), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n778), .A2(new_n704), .A3(new_n871), .A4(new_n748), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n509), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n708), .B2(new_n286), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n644), .A2(new_n647), .ZN(new_n876));
  INV_X1    g690(.A(new_n438), .ZN(new_n877));
  INV_X1    g691(.A(new_n440), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(KEYINPUT110), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n438), .B2(new_n440), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n876), .A2(new_n673), .A3(new_n678), .A4(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n833), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n873), .A2(new_n783), .A3(new_n884), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n557), .B(new_n658), .C1(new_n553), .C2(new_n554), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n389), .A2(new_n882), .A3(new_n394), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n638), .B(new_n886), .C1(new_n887), .C2(new_n632), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n596), .A2(new_n670), .A3(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n760), .B1(new_n759), .B2(new_n595), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n777), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n779), .A2(new_n780), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n868), .A2(new_n885), .A3(new_n889), .A4(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n705), .A2(new_n680), .A3(new_n749), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n775), .A2(new_n451), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n676), .B(new_n667), .C1(new_n588), .C2(new_n589), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n603), .A2(new_n900), .A3(new_n682), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n694), .B2(new_n695), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n897), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n875), .B(new_n674), .C1(new_n679), .C2(new_n704), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n899), .A2(new_n669), .A3(new_n676), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n696), .A2(new_n743), .A3(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n907), .A3(KEYINPUT52), .A4(new_n749), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n866), .B1(new_n896), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n908), .ZN(new_n911));
  AND4_X1   g725(.A1(new_n728), .A2(new_n889), .A3(new_n746), .A4(new_n867), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n873), .A2(new_n783), .A3(new_n884), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n781), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n890), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n913), .A2(new_n781), .A3(new_n890), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(KEYINPUT112), .A3(new_n911), .A4(new_n912), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n910), .A2(new_n916), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n915), .B(KEYINPUT53), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n920), .B(KEYINPUT113), .C1(new_n921), .C2(new_n917), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n916), .A2(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT113), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n923), .A2(new_n924), .A3(new_n917), .A4(new_n910), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n865), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n826), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NAND2_X1  g742(.A1(new_n544), .A2(new_n545), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT116), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT55), .Z(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n546), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n910), .A2(new_n916), .A3(new_n919), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(G210), .A3(G902), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT56), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n255), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n441), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT118), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n935), .A3(new_n932), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n934), .A2(KEYINPUT117), .A3(new_n935), .A4(new_n932), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n936), .B(new_n941), .C1(new_n944), .C2(new_n945), .ZN(G51));
  NAND2_X1  g760(.A1(new_n933), .A2(KEYINPUT54), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n920), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n933), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n502), .B(KEYINPUT57), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n499), .ZN(new_n953));
  INV_X1    g767(.A(new_n788), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n933), .A2(G902), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n939), .B1(new_n953), .B2(new_n956), .ZN(G54));
  AND4_X1   g771(.A1(KEYINPUT58), .A2(new_n933), .A3(G475), .A4(G902), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n386), .A2(new_n379), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n960), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n939), .B1(new_n961), .B2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n922), .A2(new_n925), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n606), .A2(new_n609), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n949), .A2(new_n969), .A3(new_n950), .A4(new_n965), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n968), .A2(new_n940), .A3(new_n970), .ZN(G63));
  AND2_X1   g785(.A1(new_n665), .A2(new_n666), .ZN(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  NAND3_X1  g788(.A1(new_n933), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n933), .A2(new_n977), .A3(new_n972), .A4(new_n974), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n592), .B1(new_n933), .B2(new_n974), .ZN(new_n980));
  NOR2_X1   g794(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n941), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n933), .A2(new_n974), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n941), .B1(new_n984), .B2(new_n591), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n986));
  INV_X1    g800(.A(new_n981), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n975), .A3(new_n987), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT61), .B2(new_n988), .ZN(G66));
  INV_X1    g803(.A(new_n447), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n247), .B1(new_n990), .B2(G224), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n912), .B(KEYINPUT124), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n255), .ZN(new_n993));
  INV_X1    g807(.A(G898), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n930), .B1(new_n994), .B2(new_n937), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  AOI21_X1  g810(.A(new_n255), .B1(G227), .B2(G900), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n762), .A2(new_n743), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n794), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n783), .ZN(new_n1001));
  NOR4_X1   g815(.A1(new_n1000), .A2(new_n781), .A3(new_n1001), .A4(new_n898), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n807), .A2(new_n1002), .A3(new_n255), .A4(new_n820), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n292), .A2(new_n293), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n330), .A2(new_n333), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT125), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(G900), .B2(new_n937), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n701), .A2(new_n898), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT62), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n887), .A2(new_n632), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1012), .A2(new_n699), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n709), .A3(new_n833), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1011), .A2(new_n807), .A3(new_n820), .A4(new_n1014), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(new_n255), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1007), .B(KEYINPUT126), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n998), .B(new_n1009), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1009), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1015), .B2(new_n255), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n997), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(G72));
  XNOR2_X1  g836(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n734), .A2(new_n280), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1023), .B(new_n1024), .Z(new_n1025));
  NAND3_X1  g839(.A1(new_n807), .A2(new_n1002), .A3(new_n820), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n992), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1027), .A2(new_n242), .A3(new_n264), .A4(new_n294), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1025), .B1(new_n1015), .B2(new_n992), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(new_n689), .ZN(new_n1030));
  INV_X1    g844(.A(new_n921), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1025), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n294), .A2(new_n296), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1032), .B1(new_n269), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n939), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g849(.A1(new_n1028), .A2(new_n1030), .A3(new_n1035), .ZN(G57));
endmodule


