//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT67), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  OAI211_X1 g039(.A(new_n464), .B(G125), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT66), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n473), .A3(G137), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n460), .A2(new_n461), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT66), .B(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT69), .A4(G137), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n478), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n475), .A2(new_n486), .ZN(G160));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n483), .C2(G112), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n474), .A2(new_n484), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n481), .B2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n484), .A2(KEYINPUT70), .A3(new_n470), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(G136), .B2(new_n496), .ZN(G162));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n460), .B2(new_n461), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n471), .A2(new_n473), .A3(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n504), .B2(new_n481), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n483), .A2(new_n484), .A3(new_n506), .A4(G138), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(G75), .A2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n515), .B2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n515), .A2(G651), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n520), .A2(G50), .A3(G543), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(new_n511), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n514), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AOI22_X1  g102(.A1(new_n516), .A2(new_n519), .B1(new_n515), .B2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G51), .A3(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n524), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n520), .A2(new_n521), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(G52), .A2(new_n542), .B1(new_n536), .B2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n510), .A2(new_n511), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(KEYINPUT72), .A3(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n518), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n543), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n536), .A2(G81), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n528), .A2(G43), .A3(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n545), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND4_X1  g142(.A1(new_n520), .A2(G53), .A3(G543), .A4(new_n521), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n545), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n536), .A2(G91), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  NAND4_X1  g149(.A1(new_n520), .A2(G87), .A3(new_n521), .A4(new_n523), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n528), .A2(KEYINPUT73), .A3(G87), .A4(new_n523), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n520), .A2(G49), .A3(G543), .A4(new_n521), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(G288));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n510), .B2(new_n511), .ZN(new_n585));
  AND2_X1   g160(.A1(G73), .A2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n520), .A2(G86), .A3(new_n521), .A4(new_n523), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n545), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n518), .B1(new_n593), .B2(KEYINPUT74), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(KEYINPUT74), .B2(new_n593), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT75), .B(G47), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n542), .A2(new_n596), .B1(new_n536), .B2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(G290));
  NAND4_X1  g173(.A1(new_n520), .A2(G92), .A3(new_n521), .A4(new_n523), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n545), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n542), .A2(G54), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(KEYINPUT76), .B1(G299), .B2(new_n607), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(KEYINPUT76), .B2(new_n611), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(KEYINPUT76), .B2(new_n611), .ZN(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT77), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n620), .A2(KEYINPUT78), .B1(G868), .B2(new_n562), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(KEYINPUT78), .B2(new_n620), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n484), .A2(new_n477), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n496), .A2(G135), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT80), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n483), .C2(G111), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n490), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n628), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n629), .B2(new_n635), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  OAI21_X1  g227(.A(G14), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(new_n655), .ZN(new_n662));
  INV_X1    g237(.A(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n658), .A3(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(new_n657), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n660), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n671), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n677), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  NAND3_X1  g261(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT25), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n496), .A2(G139), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n688), .B(new_n689), .C1(new_n483), .C2(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(G33), .B(new_n691), .S(G29), .Z(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(G2072), .Z(new_n693));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G34), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(G34), .ZN(new_n697));
  AOI21_X1  g272(.A(G29), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(G160), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G2084), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(G2084), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G5), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G301), .B2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n693), .A2(new_n702), .A3(new_n703), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G32), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n496), .A2(G141), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT26), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n715), .A2(new_n716), .B1(G105), .B2(new_n477), .ZN(new_n717));
  INV_X1    g292(.A(G129), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n490), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n711), .B1(new_n720), .B2(new_n700), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT27), .B(G1996), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n700), .A2(G27), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G164), .B2(new_n700), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G2078), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n700), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n700), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2090), .ZN(new_n734));
  INV_X1    g309(.A(G2090), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n721), .A2(new_n723), .B1(G2078), .B2(new_n726), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n728), .A2(new_n734), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n710), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n700), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n474), .A2(new_n484), .A3(G128), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT86), .Z(new_n743));
  OAI221_X1 g318(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n483), .C2(G116), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n496), .A2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2067), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n704), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n615), .B2(new_n704), .ZN(new_n751));
  INV_X1    g326(.A(G1348), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n704), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n562), .B2(new_n704), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(G1341), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n749), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n704), .A2(G21), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G168), .B2(new_n704), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n761), .A2(G1966), .B1(new_n707), .B2(new_n708), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G11), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT30), .B(G28), .Z(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n635), .B2(G29), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n761), .A2(G1966), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n704), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT90), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT89), .B(G1956), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n757), .B2(new_n758), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n739), .A2(new_n759), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n704), .A2(G23), .ZN(new_n780));
  INV_X1    g355(.A(G288), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(new_n704), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT33), .B(G1976), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n704), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n704), .ZN(new_n786));
  INV_X1    g361(.A(G1971), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G6), .B(G305), .S(G16), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT85), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT35), .B(G1991), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT83), .B1(G95), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(KEYINPUT83), .A2(G95), .A3(G2105), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n800), .A2(new_n801), .A3(new_n476), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G107), .B2(new_n483), .ZN(new_n803));
  INV_X1    g378(.A(G119), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n490), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G131), .B2(new_n496), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT84), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n700), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n700), .A2(G25), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n798), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n809), .A2(new_n810), .A3(new_n798), .ZN(new_n812));
  MUX2_X1   g387(.A(G24), .B(G290), .S(G16), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1986), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n796), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT36), .B1(new_n795), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n793), .B(KEYINPUT85), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n779), .B1(new_n817), .B2(new_n821), .ZN(G311));
  XNOR2_X1  g397(.A(G311), .B(KEYINPUT91), .ZN(G150));
  NAND3_X1  g398(.A1(new_n528), .A2(G93), .A3(new_n523), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT93), .B(G55), .Z(new_n825));
  NAND3_X1  g400(.A1(new_n528), .A2(G543), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n510), .B2(new_n511), .ZN(new_n828));
  AND2_X1   g403(.A1(G80), .A2(G543), .ZN(new_n829));
  OAI21_X1  g404(.A(G651), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n824), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT94), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT94), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n824), .A2(new_n826), .A3(new_n830), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND3_X1  g412(.A1(new_n832), .A2(new_n561), .A3(new_n834), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n831), .A2(new_n555), .A3(new_n556), .A4(new_n560), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT95), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n615), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT96), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n837), .B1(new_n851), .B2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n691), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n720), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n720), .ZN(new_n858));
  OAI221_X1 g433(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n483), .C2(G118), .ZN(new_n859));
  INV_X1    g434(.A(G130), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n859), .B1(new_n860), .B2(new_n490), .C1(new_n495), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n626), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n857), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n505), .A2(new_n507), .ZN(new_n868));
  INV_X1    g443(.A(new_n503), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n747), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n806), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n806), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n866), .B2(new_n865), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(G160), .B(KEYINPUT97), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n879), .B(new_n635), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n881), .B2(new_n877), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g459(.A(new_n619), .B(new_n844), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n569), .A2(new_n601), .A3(new_n573), .A4(new_n605), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n569), .A2(new_n573), .B1(new_n601), .B2(new_n605), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT99), .Z(new_n890));
  AND2_X1   g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT41), .B1(new_n887), .B2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(G299), .A2(new_n606), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n885), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n891), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n891), .B2(new_n897), .ZN(new_n900));
  XOR2_X1   g475(.A(G303), .B(G305), .Z(new_n901));
  XNOR2_X1  g476(.A(G290), .B(new_n781), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(KEYINPUT100), .ZN(new_n903));
  XNOR2_X1  g478(.A(G290), .B(G288), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n901), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n909), .A2(KEYINPUT101), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(KEYINPUT101), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT42), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT42), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n914), .A3(new_n911), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n899), .A2(new_n900), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(new_n900), .A3(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(G868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n835), .A2(new_n607), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(G295));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n919), .ZN(G331));
  INV_X1    g496(.A(new_n909), .ZN(new_n922));
  XNOR2_X1  g497(.A(G301), .B(G286), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n838), .A2(new_n842), .A3(new_n839), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(G301), .A2(G286), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n543), .A2(new_n552), .B1(new_n537), .B2(new_n535), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n841), .A2(new_n929), .A3(new_n843), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n892), .A2(new_n933), .A3(new_n895), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n889), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n934), .A2(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT105), .B1(new_n939), .B2(new_n931), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT103), .B1(new_n844), .B2(new_n923), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT103), .B1(new_n926), .B2(new_n930), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n943), .A2(new_n890), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n922), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n896), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n932), .A2(new_n889), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n922), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G37), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT106), .B1(new_n946), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n937), .B1(new_n932), .B2(new_n936), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n931), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n931), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n942), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n953), .B(new_n954), .C1(new_n957), .C2(new_n890), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n909), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n950), .A4(new_n949), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n922), .B1(new_n947), .B2(new_n948), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n951), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n959), .A2(new_n966), .A3(new_n950), .A4(new_n949), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n966), .B2(new_n965), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n963), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n968), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NOR3_X1   g548(.A1(G164), .A2(new_n973), .A3(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n475), .A2(G40), .A3(new_n486), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(G164), .B2(G1384), .ZN(new_n977));
  AOI21_X1  g552(.A(G1971), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n475), .A2(G40), .A3(new_n486), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n870), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n735), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT108), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n988));
  NAND2_X1  g563(.A1(G303), .A2(G8), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT109), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT110), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n993), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT110), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G164), .A2(G1384), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(G40), .A3(new_n475), .A4(new_n486), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n579), .A2(G1976), .A3(new_n582), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1000), .A2(G8), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G305), .A2(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1007), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1010), .A2(G8), .A3(new_n1002), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n870), .A2(new_n981), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1003), .B(G8), .C1(new_n1013), .C2(new_n975), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n995), .A2(new_n998), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n999), .A3(new_n781), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n1007), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(G8), .A3(new_n1002), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1016), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1004), .A2(new_n1012), .A3(new_n1015), .A4(KEYINPUT114), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n995), .A2(new_n998), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n983), .A2(G40), .A3(new_n475), .A4(new_n486), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n982), .A2(new_n1030), .ZN(new_n1031));
  NOR4_X1   g606(.A1(G164), .A2(new_n1030), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1029), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n978), .B1(new_n1034), .B2(new_n735), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  OAI211_X1 g611(.A(KEYINPUT113), .B(new_n997), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n980), .B1(new_n870), .B2(new_n981), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n975), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT112), .B1(new_n1001), .B2(new_n980), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1040), .B(new_n735), .C1(new_n1041), .C2(new_n1032), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n979), .A2(new_n977), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n787), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1038), .B1(new_n1046), .B2(new_n996), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n979), .A2(new_n1049), .A3(new_n1043), .A4(new_n977), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(KEYINPUT124), .A3(KEYINPUT53), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT124), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n979), .A2(new_n982), .A3(new_n983), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1052), .A2(new_n1055), .B1(new_n708), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1050), .A2(KEYINPUT123), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT123), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G301), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1051), .A2(KEYINPUT53), .B1(new_n708), .B2(new_n1056), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(G301), .C1(new_n1060), .C2(new_n1059), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT54), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1028), .B(new_n1048), .C1(new_n1062), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1056), .A2(G2084), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1966), .B1(new_n976), .B2(new_n977), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1966), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1044), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1072), .B(KEYINPUT121), .C1(G2084), .C2(new_n1056), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1073), .A3(G168), .ZN(new_n1074));
  AND2_X1   g649(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G168), .A2(new_n1036), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1074), .A2(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1036), .B(G168), .C1(new_n1070), .C2(new_n1073), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1057), .A2(new_n1061), .A3(G301), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1063), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1084));
  OAI21_X1  g659(.A(G171), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT54), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1066), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(G299), .B(KEYINPUT57), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n976), .A2(new_n977), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1089), .B(new_n1091), .C1(G1956), .C2(new_n1034), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1034), .B2(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1088), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n975), .A2(new_n1013), .ZN(new_n1096));
  INV_X1    g671(.A(G2067), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1056), .A2(new_n752), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n606), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(KEYINPUT117), .B(new_n1092), .C1(new_n1095), .C2(new_n1099), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1093), .A2(KEYINPUT120), .A3(new_n1088), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1092), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1094), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1098), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT118), .B(G1996), .Z(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1044), .A2(new_n1111), .B1(new_n1096), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n562), .ZN(new_n1114));
  NAND2_X1  g689(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1110), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1094), .A2(new_n1092), .A3(KEYINPUT61), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1098), .A2(KEYINPUT60), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1098), .A2(KEYINPUT60), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n615), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1102), .B(new_n1103), .C1(new_n1109), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1024), .B1(new_n1087), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1076), .A2(G286), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1028), .A2(new_n1048), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT63), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1028), .A2(new_n1048), .A3(KEYINPUT115), .A4(new_n1126), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n985), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n997), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n995), .A2(new_n998), .ZN(new_n1137));
  NOR4_X1   g712(.A1(new_n1076), .A2(new_n1016), .A3(new_n1130), .A4(G286), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1079), .A2(new_n1080), .A3(KEYINPUT62), .ZN(new_n1141));
  AOI21_X1  g716(.A(G301), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1028), .A2(new_n1048), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT125), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1028), .A2(new_n1048), .A3(new_n1142), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1077), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1146), .B(new_n1148), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1145), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT62), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1144), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1125), .A2(new_n1140), .A3(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n806), .B(new_n798), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n975), .A2(new_n977), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n747), .A2(G2067), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n745), .A2(new_n1097), .A3(new_n746), .ZN(new_n1162));
  INV_X1    g737(.A(G1996), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1161), .B(new_n1162), .C1(new_n1163), .C2(new_n720), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1158), .ZN(new_n1165));
  INV_X1    g740(.A(new_n720), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT107), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(G290), .B(G1986), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1160), .B(new_n1169), .C1(new_n1158), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1156), .A2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1168), .B(KEYINPUT46), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1161), .A2(new_n720), .A3(new_n1162), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1158), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1176), .A2(KEYINPUT47), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(KEYINPUT47), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(KEYINPUT126), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n808), .A2(new_n797), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1162), .B1(new_n1169), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1169), .A2(new_n1160), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1159), .A2(G1986), .A3(G290), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1181), .A2(new_n1158), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1179), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(KEYINPUT126), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1172), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g765(.A(G319), .ZN(new_n1192));
  NOR4_X1   g766(.A1(G401), .A2(G229), .A3(new_n1192), .A4(G227), .ZN(new_n1193));
  NAND3_X1  g767(.A1(new_n970), .A2(new_n883), .A3(new_n1193), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


