//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G58), .C2(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  INV_X1    g0023(.A(new_n201), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n225), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G13), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT0), .Z(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n227), .A3(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  INV_X1    g0036(.A(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n210), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n209), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND3_X1  g0050(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT68), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G77), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT66), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n255), .A2(new_n256), .B1(new_n220), .B2(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n220), .A2(G33), .ZN(new_n261));
  XOR2_X1   g0061(.A(KEYINPUT15), .B(G87), .Z(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n226), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n253), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n266), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n219), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(KEYINPUT68), .A3(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n257), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G232), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G107), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(G1698), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n279), .B1(new_n280), .B2(new_n277), .C1(new_n281), .C2(new_n214), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n283), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n274), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G244), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n267), .A2(new_n272), .B1(new_n273), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n289), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G200), .B2(new_n289), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n253), .B(new_n271), .C1(new_n264), .C2(new_n266), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n290), .A2(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n203), .A2(G20), .ZN(new_n299));
  INV_X1    g0099(.A(G150), .ZN(new_n300));
  INV_X1    g0100(.A(new_n254), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT8), .A2(G58), .ZN(new_n302));
  OR2_X1    g0102(.A1(KEYINPUT65), .A2(G58), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT65), .A2(G58), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT8), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n299), .B1(new_n300), .B2(new_n301), .C1(new_n307), .C2(new_n261), .ZN(new_n308));
  INV_X1    g0108(.A(new_n251), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n308), .A2(new_n266), .B1(new_n202), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n268), .A2(G50), .A3(new_n269), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT9), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n277), .A2(G222), .A3(new_n278), .ZN(new_n317));
  INV_X1    g0117(.A(G223), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n257), .B2(new_n277), .C1(new_n281), .C2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n283), .B1(G226), .B2(new_n287), .ZN(new_n320));
  INV_X1    g0120(.A(new_n276), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n294), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT10), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n329), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n316), .A2(new_n326), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n322), .A2(new_n273), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(new_n312), .C1(G179), .C2(new_n322), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n298), .A2(new_n330), .A3(new_n333), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT70), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n277), .A2(G226), .A3(new_n278), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n277), .A2(G232), .A3(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n283), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n287), .A2(G238), .ZN(new_n346));
  AND4_X1   g0146(.A1(new_n340), .A2(new_n345), .A3(new_n346), .A4(new_n321), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n276), .B1(new_n344), .B2(new_n283), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n340), .B1(new_n348), .B2(new_n346), .ZN(new_n349));
  OAI21_X1  g0149(.A(G169), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(new_n340), .A3(new_n346), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n349), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n340), .A4(new_n346), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(G179), .A4(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(G169), .C1(new_n347), .C2(new_n349), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n351), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n213), .A2(G20), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n361), .B1(new_n261), .B2(new_n257), .C1(new_n301), .C2(new_n202), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n266), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT72), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n365), .A3(new_n266), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT11), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n270), .A2(KEYINPUT12), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G68), .ZN(new_n370));
  INV_X1    g0170(.A(new_n252), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n370), .B(new_n372), .C1(KEYINPUT12), .C2(new_n309), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT73), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n368), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n360), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n368), .A2(new_n375), .A3(new_n376), .ZN(new_n379));
  OAI21_X1  g0179(.A(G200), .B1(new_n347), .B2(new_n349), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n354), .A2(new_n355), .A3(G190), .A4(new_n356), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NOR2_X1   g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  OAI211_X1 g0185(.A(G226), .B(G1698), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(G223), .B(new_n278), .C1(new_n384), .C2(new_n385), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n283), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n285), .A2(G232), .A3(new_n274), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n321), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(G190), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n276), .B1(new_n389), .B2(new_n283), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n394), .A2(KEYINPUT75), .A3(new_n391), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT75), .B1(new_n394), .B2(new_n391), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n397), .B2(new_n324), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n303), .A2(G68), .A3(new_n304), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n220), .B1(new_n400), .B2(new_n224), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n301), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n399), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n403), .ZN(new_n405));
  AND2_X1   g0205(.A1(KEYINPUT65), .A2(G58), .ZN(new_n406));
  NOR2_X1   g0206(.A1(KEYINPUT65), .A2(G58), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n201), .B1(new_n408), .B2(G68), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT74), .B(new_n405), .C1(new_n409), .C2(new_n220), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n277), .B2(G20), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n384), .A2(new_n385), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n213), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(KEYINPUT16), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n405), .B1(new_n409), .B2(new_n220), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n416), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n266), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n307), .A2(new_n309), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n268), .A2(new_n269), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n307), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(KEYINPUT17), .B1(new_n398), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n416), .B1(new_n404), .B2(new_n410), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n268), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n425), .B1(new_n430), .B2(new_n421), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n392), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n394), .A2(KEYINPUT75), .A3(new_n391), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n324), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G190), .B2(new_n392), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT18), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n433), .A2(new_n273), .A3(new_n434), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G179), .B2(new_n392), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n431), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n392), .A2(G179), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n397), .B2(new_n273), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n427), .A3(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n338), .A2(new_n339), .A3(new_n383), .A4(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n220), .B(G87), .C1(new_n384), .C2(new_n385), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT83), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n277), .A2(new_n453), .A3(new_n220), .A4(G87), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT22), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n220), .A2(G107), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT23), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT22), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(KEYINPUT83), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n220), .A2(G33), .A3(G116), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n455), .A2(new_n457), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT24), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n459), .A2(new_n460), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n457), .A4(new_n455), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n266), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n251), .A2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT25), .ZN(new_n470));
  INV_X1    g0270(.A(G33), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n268), .A2(new_n251), .A3(new_n473), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n474), .A2(new_n280), .B1(new_n469), .B2(KEYINPUT25), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n467), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n277), .A2(G250), .A3(new_n278), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n277), .A2(G257), .A3(G1698), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n277), .A2(new_n481), .A3(G250), .A4(new_n278), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G294), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n479), .A2(new_n480), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n285), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n484), .A2(new_n283), .B1(G264), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n489), .A2(new_n275), .ZN(new_n492));
  AOI21_X1  g0292(.A(G169), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n491), .A2(new_n292), .A3(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n477), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n475), .B1(new_n466), .B2(new_n266), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(new_n492), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(G190), .A3(new_n492), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n470), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n498), .B1(new_n497), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n474), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n262), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n205), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT78), .A2(KEYINPUT19), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n511), .A2(new_n512), .A3(new_n343), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(G20), .ZN(new_n514));
  INV_X1    g0314(.A(new_n385), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT3), .A2(G33), .ZN(new_n516));
  AOI21_X1  g0316(.A(G20), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G68), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n220), .A2(G33), .A3(G97), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT78), .B(KEYINPUT19), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n514), .A2(new_n518), .A3(new_n521), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n266), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n252), .A2(new_n262), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT80), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n530), .B(new_n527), .C1(new_n525), .C2(new_n266), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n508), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n277), .A2(G238), .A3(new_n278), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n277), .A2(G244), .A3(G1698), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G116), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n283), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n486), .A2(G274), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n285), .B(G250), .C1(G1), .C2(new_n485), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n292), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n273), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n521), .A2(new_n524), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n220), .B1(new_n522), .B2(new_n343), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n510), .B1(G68), .B2(new_n517), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n268), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n530), .B1(new_n548), .B2(new_n527), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n528), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n541), .A2(G190), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n474), .A2(new_n509), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n540), .A2(G200), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n551), .A2(new_n552), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n544), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT81), .ZN(new_n558));
  OAI211_X1 g0358(.A(G244), .B(new_n278), .C1(new_n384), .C2(new_n385), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT4), .B1(new_n560), .B2(KEYINPUT77), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n277), .A2(G250), .A3(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G283), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n561), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n283), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n490), .A2(G257), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n492), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT6), .B1(new_n206), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(KEYINPUT6), .A2(G97), .ZN(new_n574));
  OAI21_X1  g0374(.A(KEYINPUT76), .B1(new_n574), .B2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n280), .A3(KEYINPUT6), .A4(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n579), .A2(new_n220), .B1(new_n257), .B2(new_n301), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n280), .B1(new_n413), .B2(new_n415), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n266), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n251), .A2(G97), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n507), .A2(G97), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n571), .B(new_n587), .C1(new_n294), .C2(new_n570), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n570), .A2(new_n273), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n568), .A2(new_n292), .A3(new_n492), .A4(new_n569), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n371), .A2(new_n209), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n252), .A2(G116), .A3(new_n268), .A4(new_n473), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n209), .A2(G20), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT82), .B1(new_n266), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n595), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n566), .B(new_n220), .C1(G33), .C2(new_n215), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT20), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n266), .A2(KEYINPUT82), .A3(new_n595), .ZN(new_n602));
  OAI211_X1 g0402(.A(KEYINPUT20), .B(new_n600), .C1(new_n602), .C2(new_n596), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n593), .B(new_n594), .C1(new_n601), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n277), .A2(G257), .A3(new_n278), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  INV_X1    g0408(.A(G264), .ZN(new_n609));
  OAI221_X1 g0409(.A(new_n607), .B1(new_n608), .B2(new_n277), .C1(new_n281), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n283), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n490), .A2(G270), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n492), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G200), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n606), .B(new_n614), .C1(new_n294), .C2(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n605), .A2(G169), .A3(new_n613), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n613), .A2(new_n292), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n605), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n605), .A2(new_n613), .A3(KEYINPUT21), .A4(G169), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n615), .A2(new_n618), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT81), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n544), .A2(new_n624), .A3(new_n556), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n558), .A2(new_n592), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n450), .A2(new_n506), .A3(new_n626), .ZN(G372));
  INV_X1    g0427(.A(new_n447), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n267), .A2(new_n272), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n289), .A2(new_n273), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n629), .A2(new_n630), .A3(new_n293), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n382), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n378), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT87), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n633), .A2(KEYINPUT87), .B1(new_n428), .B2(new_n438), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n330), .A2(new_n333), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n335), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n591), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT86), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n543), .A2(new_n642), .B1(new_n541), .B2(new_n292), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n273), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n532), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n641), .A2(new_n645), .A3(new_n646), .A4(new_n556), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n503), .A2(new_n588), .A3(new_n591), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n497), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n556), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n544), .A2(new_n624), .A3(new_n556), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n624), .B1(new_n544), .B2(new_n556), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n655), .A2(new_n656), .A3(new_n591), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n648), .B(new_n654), .C1(new_n657), .C2(new_n646), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n640), .B1(new_n450), .B2(new_n659), .ZN(G369));
  AOI211_X1 g0460(.A(new_n493), .B(new_n495), .C1(new_n499), .C2(new_n470), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n470), .A2(new_n499), .A3(new_n501), .A4(new_n502), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT85), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n497), .A2(new_n498), .A3(new_n503), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n228), .A2(G20), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n219), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT88), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n477), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n665), .A2(new_n675), .B1(new_n661), .B2(new_n674), .ZN(new_n676));
  INV_X1    g0476(.A(new_n650), .ZN(new_n677));
  INV_X1    g0477(.A(new_n674), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n606), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n622), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g0481(.A(KEYINPUT89), .B(G330), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n497), .A2(new_n674), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n677), .A2(new_n678), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n665), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n685), .A2(new_n689), .ZN(G399));
  NAND3_X1  g0490(.A1(new_n205), .A2(new_n509), .A3(new_n209), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT90), .Z(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n229), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n225), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n558), .A2(new_n646), .A3(new_n641), .A4(new_n625), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT26), .B1(new_n652), .B2(new_n591), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n654), .A2(new_n699), .A3(new_n645), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n678), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n658), .A2(new_n704), .A3(new_n678), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n682), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n655), .A2(new_n656), .A3(new_n622), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n665), .A2(new_n592), .A3(new_n709), .A4(new_n678), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n613), .A2(new_n292), .A3(new_n540), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n568), .A2(new_n492), .A3(new_n569), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n712), .A3(new_n491), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n613), .A2(new_n292), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n500), .A3(new_n570), .A4(new_n540), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n674), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(new_n674), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n708), .B1(new_n710), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n707), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n698), .B1(new_n728), .B2(G1), .ZN(G364));
  AOI21_X1  g0529(.A(new_n219), .B1(new_n666), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n694), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT91), .Z(new_n733));
  OR2_X1    g0533(.A1(new_n681), .A2(new_n682), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n683), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n226), .B1(G20), .B2(new_n273), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n294), .A2(new_n324), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n220), .A2(G179), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n509), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n414), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n324), .A2(G190), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G107), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n294), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n292), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n741), .B(new_n745), .C1(new_n215), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(G20), .A2(G179), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n737), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n742), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n202), .A2(new_n754), .B1(new_n755), .B2(new_n213), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n746), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n750), .B(new_n756), .C1(new_n408), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G190), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n738), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n402), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n763));
  XNOR2_X1  g0563(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n753), .A2(new_n760), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n759), .B(new_n764), .C1(new_n257), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT95), .Z(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  INV_X1    g0568(.A(G326), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n757), .B1(new_n754), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n755), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n739), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G303), .ZN(new_n775));
  INV_X1    g0575(.A(new_n761), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n414), .B(new_n777), .C1(new_n749), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G283), .B2(new_n744), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n765), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G311), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n736), .B1(new_n767), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n246), .A2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n229), .A2(new_n277), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(G45), .C2(new_n225), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n230), .A2(G355), .A3(new_n277), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(G116), .C2(new_n230), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT92), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n736), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n792), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n784), .B(new_n794), .C1(new_n681), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n735), .B1(new_n796), .B2(new_n733), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT96), .Z(G396));
  INV_X1    g0598(.A(new_n733), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n800), .A2(new_n754), .B1(new_n755), .B2(new_n300), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g0602(.A1(new_n758), .A2(G143), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n402), .C2(new_n765), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT34), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n743), .A2(new_n213), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n277), .B1(new_n749), .B2(new_n305), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G50), .C2(new_n774), .ZN(new_n808));
  INV_X1    g0608(.A(G132), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n805), .B(new_n808), .C1(new_n809), .C2(new_n761), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n744), .A2(G87), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n280), .B2(new_n739), .C1(new_n749), .C2(new_n215), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n277), .B(new_n812), .C1(G311), .C2(new_n776), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT98), .B(G283), .Z(new_n814));
  OAI22_X1  g0614(.A1(new_n778), .A2(new_n757), .B1(new_n755), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n754), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G303), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n813), .B(new_n817), .C1(new_n209), .C2(new_n765), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n810), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n799), .B1(new_n819), .B2(new_n736), .ZN(new_n820));
  INV_X1    g0620(.A(new_n791), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n736), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT97), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n257), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n631), .A2(KEYINPUT100), .A3(new_n674), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n290), .A2(new_n293), .A3(new_n674), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n629), .A2(new_n674), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n825), .A2(new_n828), .B1(new_n298), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n820), .B(new_n824), .C1(new_n791), .C2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n558), .A2(new_n641), .A3(new_n625), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n652), .B1(new_n650), .B2(new_n497), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(KEYINPUT26), .B1(new_n834), .B2(new_n649), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n674), .B1(new_n835), .B2(new_n648), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(new_n830), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(new_n725), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n832), .B1(new_n838), .B2(new_n733), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n445), .A2(new_n427), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n431), .A2(new_n436), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n427), .A2(new_n671), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n411), .A2(new_n417), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n419), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n425), .B1(new_n430), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT102), .B1(new_n847), .B2(new_n672), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n418), .A2(new_n266), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n429), .A2(KEYINPUT16), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n426), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(new_n671), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n445), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n848), .A2(new_n853), .A3(new_n842), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n844), .B1(KEYINPUT37), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n439), .A2(new_n447), .B1(new_n853), .B2(new_n848), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n840), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n848), .A2(new_n853), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n448), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT39), .B1(new_n859), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT103), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n439), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n428), .A2(KEYINPUT104), .A3(new_n438), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(new_n447), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n843), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n874), .A2(new_n875), .B1(new_n861), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n869), .B(new_n870), .C1(new_n878), .C2(KEYINPUT38), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n870), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(KEYINPUT103), .A3(KEYINPUT39), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n868), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n378), .A2(new_n674), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n377), .A2(new_n674), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n378), .A2(new_n382), .A3(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT101), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT101), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n360), .A2(new_n377), .A3(new_n674), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n658), .A2(new_n831), .A3(new_n678), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n631), .A2(new_n678), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n896), .A2(new_n881), .B1(new_n628), .B2(new_n672), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  AOI211_X1 g0698(.A(KEYINPUT105), .B(new_n450), .C1(new_n703), .C2(new_n705), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  INV_X1    g0700(.A(new_n339), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n383), .B1(new_n336), .B2(new_n337), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n901), .A2(new_n902), .A3(new_n448), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n900), .B1(new_n706), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n640), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n898), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n830), .B1(new_n891), .B2(new_n892), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n710), .A2(new_n724), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n881), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n870), .B1(new_n878), .B2(KEYINPUT38), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n912), .A2(KEYINPUT40), .A3(new_n908), .A4(new_n907), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n903), .A2(new_n908), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n708), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n906), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n219), .B2(new_n666), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT35), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n220), .B(new_n226), .C1(new_n579), .C2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(G116), .C1(new_n920), .C2(new_n579), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n400), .A2(G50), .A3(G77), .A4(new_n224), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(G50), .B2(new_n213), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n228), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n923), .A3(new_n926), .ZN(G367));
  NOR2_X1   g0727(.A1(new_n743), .A2(new_n257), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n816), .A2(G143), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n928), .B(new_n929), .C1(G150), .C2(new_n758), .ZN(new_n930));
  AOI22_X1  g0730(.A1(G50), .A2(new_n782), .B1(new_n771), .B2(G159), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(KEYINPUT109), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n749), .A2(new_n213), .B1(new_n739), .B2(new_n305), .ZN(new_n934));
  AOI211_X1 g0734(.A(new_n414), .B(new_n934), .C1(G137), .C2(new_n776), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n930), .A2(new_n932), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT46), .B1(new_n774), .B2(G116), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n816), .A2(G311), .B1(G107), .B2(new_n748), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n778), .B2(new_n755), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n414), .B1(new_n761), .B2(new_n940), .C1(new_n215), .C2(new_n743), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT108), .Z(new_n942));
  NAND3_X1  g0742(.A1(new_n774), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(new_n765), .B2(new_n814), .C1(new_n608), .C2(new_n757), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n936), .B1(new_n937), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT110), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n736), .ZN(new_n949));
  INV_X1    g0749(.A(new_n786), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n793), .B1(new_n230), .B2(new_n263), .C1(new_n242), .C2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n949), .A2(new_n733), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT111), .Z(new_n953));
  INV_X1    g0753(.A(new_n551), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n674), .B1(new_n954), .B2(new_n553), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n653), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n645), .B2(new_n955), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n957), .A2(new_n795), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n674), .A2(new_n586), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n592), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n641), .A2(new_n674), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n689), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(KEYINPUT107), .A3(new_n966), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n964), .A2(KEYINPUT107), .A3(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n689), .A2(new_n963), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n684), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n676), .A2(new_n687), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n665), .A2(new_n688), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n683), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n727), .ZN(new_n977));
  INV_X1    g0777(.A(new_n971), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n967), .A2(new_n978), .A3(new_n685), .A4(new_n968), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n972), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n728), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n982));
  XOR2_X1   g0782(.A(new_n694), .B(new_n982), .Z(new_n983));
  AOI21_X1  g0783(.A(new_n731), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n974), .A2(new_n961), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n986), .A2(new_n987), .B1(new_n591), .B2(new_n674), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n686), .A2(new_n987), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n689), .A2(new_n961), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n985), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n684), .A2(new_n963), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n959), .B1(new_n984), .B2(new_n995), .ZN(G387));
  AOI22_X1  g0796(.A1(G303), .A2(new_n782), .B1(new_n816), .B2(G322), .ZN(new_n997));
  INV_X1    g0797(.A(G311), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n998), .B2(new_n755), .C1(new_n940), .C2(new_n757), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n778), .B2(new_n739), .C1(new_n749), .C2(new_n814), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT49), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n277), .B1(new_n744), .B2(G116), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n769), .C2(new_n761), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n749), .A2(new_n263), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G77), .B2(new_n774), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n414), .B1(new_n744), .B2(G97), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(new_n300), .C2(new_n761), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n758), .A2(G50), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n213), .B2(new_n765), .C1(new_n307), .C2(new_n755), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n816), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT113), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n799), .B1(new_n1013), .B2(new_n736), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n256), .A2(G50), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1016));
  AND2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n485), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n213), .A2(new_n257), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n692), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n786), .B1(new_n238), .B2(new_n485), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n692), .A2(new_n230), .A3(new_n277), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n230), .A2(G107), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n793), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n676), .A2(new_n792), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1014), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n976), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n694), .B1(new_n1028), .B2(new_n728), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1027), .B1(new_n730), .B2(new_n976), .C1(new_n1029), .C2(new_n977), .ZN(G393));
  INV_X1    g0830(.A(KEYINPUT115), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT114), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n972), .A2(new_n1032), .A3(new_n979), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n979), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n694), .B(new_n980), .C1(new_n1034), .C2(new_n977), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n961), .A2(new_n792), .A3(new_n962), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n793), .B1(new_n215), .B2(new_n230), .C1(new_n249), .C2(new_n950), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n414), .B1(new_n761), .B2(new_n768), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n745), .B1(new_n739), .B2(new_n814), .C1(new_n749), .C2(new_n209), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G303), .C2(new_n771), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n998), .A2(new_n757), .B1(new_n754), .B2(new_n940), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n778), .C2(new_n765), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n816), .B1(new_n758), .B2(G159), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT51), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n749), .A2(new_n257), .B1(new_n739), .B2(new_n213), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n414), .B(new_n1046), .C1(G143), .C2(new_n776), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n811), .B1(new_n765), .B2(new_n256), .C1(new_n202), .C2(new_n755), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1044), .A2(KEYINPUT51), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n799), .B1(new_n1052), .B2(new_n736), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1036), .A2(new_n1037), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1034), .B2(new_n731), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1031), .B1(new_n1035), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1035), .A2(new_n1031), .A3(new_n1055), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(G390));
  INV_X1    g0859(.A(new_n884), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n895), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n701), .A2(new_n678), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n831), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1060), .B(new_n912), .C1(new_n1063), .C2(new_n893), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n896), .A2(new_n884), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n883), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n891), .A2(new_n892), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n908), .A2(G330), .A3(new_n831), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n708), .B(new_n830), .C1(new_n710), .C2(new_n724), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1067), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1064), .B(new_n1072), .C1(new_n883), .C2(new_n1065), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n731), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G107), .A2(new_n771), .B1(new_n816), .B2(G283), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n215), .B2(new_n765), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT118), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n414), .B1(new_n778), .B2(new_n761), .C1(new_n757), .C2(new_n209), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n749), .A2(new_n257), .B1(new_n213), .B2(new_n743), .ZN(new_n1080));
  NOR4_X1   g0880(.A1(new_n1078), .A2(new_n740), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n739), .A2(new_n300), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n414), .B1(new_n744), .B2(G50), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n402), .C2(new_n749), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G128), .A2(new_n816), .B1(new_n758), .B2(G132), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  NAND2_X1  g0888(.A1(new_n782), .A2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(new_n800), .C2(new_n755), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1086), .B(new_n1090), .C1(G125), .C2(new_n776), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1081), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT119), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n799), .B1(new_n1093), .B2(new_n736), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n823), .A2(new_n307), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n791), .C2(new_n883), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1075), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n908), .A2(G330), .A3(new_n831), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1071), .B(new_n1063), .C1(new_n1067), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT116), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1061), .B1(new_n836), .B2(new_n831), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n506), .A2(new_n626), .A3(new_n674), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n721), .A2(new_n723), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n682), .B(new_n831), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n893), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1103), .B(new_n1104), .C1(new_n1108), .C2(new_n1068), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1068), .B1(new_n1070), .B2(new_n1067), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n894), .A2(new_n895), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT116), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1102), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n903), .A2(G330), .A3(new_n908), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n658), .A2(new_n704), .A3(new_n678), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n704), .B1(new_n701), .B2(new_n678), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n903), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(KEYINPUT105), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n706), .A2(new_n900), .A3(new_n903), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n639), .B(new_n1115), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1074), .A2(new_n1121), .A3(new_n1113), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n694), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1075), .A2(KEYINPUT120), .A3(new_n1096), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1099), .A2(new_n1125), .A3(new_n1126), .ZN(G378));
  INV_X1    g0927(.A(KEYINPUT122), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n911), .A2(G330), .A3(new_n913), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n885), .A2(new_n897), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n885), .B2(new_n897), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n330), .A2(new_n333), .A3(new_n335), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n312), .A2(new_n671), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1132), .B(new_n1133), .Z(new_n1134));
  AND2_X1   g0934(.A1(new_n1134), .A2(KEYINPUT55), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(KEYINPUT55), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT56), .ZN(new_n1137));
  OR3_X1    g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1130), .A2(new_n1131), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1140), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1129), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT103), .B1(new_n881), .B2(KEYINPUT39), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n867), .B(new_n869), .C1(new_n880), .C2(new_n870), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1060), .B1(new_n1146), .B2(new_n879), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n897), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n885), .A2(new_n897), .A3(new_n1129), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1142), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1128), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1142), .A3(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(KEYINPUT122), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1121), .B1(new_n1100), .B2(new_n1122), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1124), .A2(new_n1121), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n695), .B1(new_n1160), .B2(KEYINPUT57), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1142), .A2(new_n821), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n822), .A2(new_n202), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n277), .A2(G41), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n776), .A2(G283), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n257), .B2(new_n739), .C1(new_n305), .C2(new_n743), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G68), .C2(new_n748), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n209), .A2(new_n754), .B1(new_n765), .B2(new_n263), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G97), .B2(new_n771), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(new_n280), .C2(new_n757), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G128), .A2(new_n758), .B1(new_n771), .B2(G132), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n782), .A2(G137), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n774), .A2(new_n1088), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n816), .A2(G125), .B1(G150), .B2(new_n748), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n776), .A2(G124), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(G33), .A2(G41), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT121), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G159), .B2(new_n744), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1165), .A2(new_n202), .A3(new_n1182), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1172), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n799), .B1(new_n1186), .B2(new_n736), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1163), .A2(new_n1164), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1155), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT122), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1189), .B1(new_n1192), .B2(new_n731), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1162), .A2(new_n1193), .ZN(G375));
  OAI21_X1  g0994(.A(new_n277), .B1(new_n743), .B2(new_n305), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n749), .A2(new_n202), .B1(new_n739), .B2(new_n402), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G128), .C2(new_n776), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1088), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n300), .A2(new_n765), .B1(new_n755), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G132), .B2(new_n816), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(new_n800), .C2(new_n757), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n280), .A2(new_n765), .B1(new_n754), .B2(new_n778), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G116), .B2(new_n771), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n928), .B(new_n1005), .C1(G97), .C2(new_n774), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n758), .A2(G283), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n277), .B1(new_n776), .B2(G303), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n799), .B1(new_n1208), .B2(new_n736), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1067), .B2(new_n791), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n213), .B2(new_n823), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1113), .B2(new_n731), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1122), .A2(new_n983), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(G381));
  XOR2_X1   g1015(.A(G375), .B(KEYINPUT123), .Z(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  INV_X1    g1017(.A(G387), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1057), .A2(new_n1218), .A3(new_n1058), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(G381), .A3(G384), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1216), .A2(new_n1217), .A3(new_n1220), .A4(new_n1221), .ZN(G407));
  NAND3_X1  g1022(.A1(new_n1216), .A2(new_n673), .A3(new_n1217), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(new_n1058), .ZN(new_n1225));
  OAI21_X1  g1025(.A(G387), .B1(new_n1225), .B2(new_n1056), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1219), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G393), .B(G396), .Z(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1228), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1219), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n673), .A2(G213), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1162), .A2(G378), .A3(new_n1193), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n731), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n983), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1157), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1217), .B1(new_n1237), .B2(new_n1189), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1233), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1241));
  AND4_X1   g1041(.A1(G330), .A2(new_n908), .A3(new_n831), .A4(new_n1067), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1067), .B1(new_n725), .B2(new_n831), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1111), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1103), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1110), .A2(KEYINPUT116), .A3(new_n1111), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n640), .B(new_n1114), .C1(new_n899), .C2(new_n904), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT60), .A4(new_n1102), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1241), .A2(new_n694), .A3(new_n1122), .A4(new_n1249), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1250), .A2(G384), .A3(new_n1212), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1250), .B2(new_n1212), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1239), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1232), .B1(new_n1255), .B2(KEYINPUT63), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT124), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1233), .A2(G2897), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(new_n1251), .A2(new_n1252), .A3(KEYINPUT124), .A4(new_n1258), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1257), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT63), .B1(new_n1239), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1254), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1239), .B2(new_n1263), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT125), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1239), .A2(new_n1253), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1254), .A2(new_n1270), .ZN(new_n1274));
  OAI211_X1 g1074(.A(KEYINPUT125), .B(new_n1266), .C1(new_n1239), .C2(new_n1263), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1269), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI221_X4 g1076(.A(KEYINPUT127), .B1(new_n1256), .B2(new_n1265), .C1(new_n1276), .C2(new_n1232), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1232), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1256), .A2(new_n1265), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1277), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1217), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1234), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1253), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1232), .ZN(G402));
endmodule


