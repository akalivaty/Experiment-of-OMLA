//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n211), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n214), .B(new_n219), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n217), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n208), .A2(G20), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G50), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G50), .B2(new_n247), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n209), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n250), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G223), .A3(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  OAI221_X1 g0074(.A(new_n270), .B1(new_n271), .B2(new_n269), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT65), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  OAI211_X1 g0084(.A(G1), .B(G13), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n285), .A2(new_n278), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G226), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n277), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G200), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n268), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT68), .B(G179), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n267), .B(new_n295), .C1(new_n297), .C2(new_n288), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT74), .ZN(new_n300));
  OR2_X1    g0100(.A1(G226), .A2(G1698), .ZN(new_n301));
  INV_X1    g0101(.A(G232), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G1698), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n269), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT72), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n276), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n279), .A2(new_n281), .B1(new_n286), .B2(G238), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT13), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n313), .A2(G179), .A3(new_n315), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n310), .A2(new_n311), .A3(new_n314), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n310), .B2(new_n311), .ZN(new_n318));
  OAI21_X1  g0118(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(KEYINPUT14), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(new_n315), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n321), .B1(new_n322), .B2(G169), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n300), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(KEYINPUT14), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n321), .A3(G169), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT74), .A4(new_n316), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n248), .A2(new_n202), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n251), .A2(G68), .A3(new_n252), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(G50), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n260), .A2(new_n333), .B1(new_n209), .B2(G68), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n262), .A2(new_n271), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n250), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n330), .B(new_n331), .C1(new_n332), .C2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n332), .B2(new_n336), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT73), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n322), .A2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n313), .A2(G190), .A3(new_n315), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n269), .A2(G238), .A3(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G33), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n283), .A2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(G107), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n346), .B(new_n351), .C1(new_n273), .C2(new_n302), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n276), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n279), .A2(new_n281), .B1(new_n286), .B2(G244), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n289), .B2(new_n355), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n247), .A2(KEYINPUT71), .A3(G77), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT71), .B1(new_n247), .B2(G77), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n271), .B1(new_n208), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n358), .A2(new_n359), .B1(new_n251), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT8), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G58), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT69), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT69), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n261), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n260), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n370), .A2(new_n262), .B1(new_n209), .B2(new_n271), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n250), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n372), .A2(new_n373), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n361), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n357), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n355), .A2(new_n294), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n353), .A2(new_n296), .A3(new_n354), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n299), .A2(new_n345), .A3(new_n377), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT82), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n286), .A2(G232), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n282), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n348), .A2(new_n349), .A3(G223), .A4(new_n272), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT79), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n269), .A2(KEYINPUT79), .A3(G223), .A4(new_n272), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n348), .A2(new_n349), .A3(G226), .A4(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n285), .B1(new_n395), .B2(KEYINPUT80), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n388), .B2(new_n389), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n385), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(KEYINPUT81), .A3(new_n289), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT81), .ZN(new_n402));
  INV_X1    g0202(.A(new_n385), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n276), .B1(new_n397), .B2(new_n398), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n390), .A2(new_n398), .A3(new_n394), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n402), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n289), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n401), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n251), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n365), .A2(new_n252), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n412), .A2(new_n413), .B1(new_n247), .B2(new_n365), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT7), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(G20), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n350), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT7), .B1(new_n350), .B2(new_n209), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(G58), .B(G68), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n250), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g0224(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n283), .B2(KEYINPUT3), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n347), .A2(KEYINPUT76), .A3(G33), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n349), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n416), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n415), .B1(new_n269), .B2(G20), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n202), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n421), .B1(new_n432), .B2(KEYINPUT77), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n434), .B(new_n202), .C1(new_n430), .C2(new_n431), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n425), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT78), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n424), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(KEYINPUT78), .B(new_n425), .C1(new_n433), .C2(new_n435), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n414), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT17), .B1(new_n411), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n383), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n436), .A2(new_n437), .ZN(new_n444));
  INV_X1    g0244(.A(new_n424), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n414), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n406), .A2(G169), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n296), .B2(new_n406), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n448), .B2(new_n451), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n409), .A2(new_n402), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT81), .B1(new_n400), .B2(G200), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n409), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(new_n448), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n411), .A2(new_n440), .A3(KEYINPUT17), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(KEYINPUT82), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n443), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n382), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n269), .A2(G264), .A3(G1698), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n269), .A2(G257), .A3(new_n272), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n350), .A2(G303), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n276), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n276), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n473), .A2(new_n472), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n474), .A2(G270), .B1(new_n475), .B2(new_n281), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n248), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n208), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n247), .A2(new_n480), .A3(new_n217), .A4(new_n249), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n249), .A2(new_n217), .B1(G20), .B2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n209), .C1(G33), .C2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT20), .B1(new_n482), .B2(new_n485), .ZN(new_n487));
  OAI221_X1 g0287(.A(new_n479), .B1(new_n478), .B2(new_n481), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n477), .A2(G169), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(G179), .A3(new_n470), .A4(new_n476), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n477), .A2(KEYINPUT21), .A3(new_n488), .A4(G169), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n488), .B1(new_n477), .B2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n289), .B2(new_n477), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n269), .A2(G238), .A3(new_n272), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n269), .A2(G244), .A3(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n276), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n208), .A2(G45), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n285), .A2(G250), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n285), .A2(G274), .A3(new_n472), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G169), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n503), .B2(new_n276), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n297), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n269), .A2(new_n209), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n209), .B1(new_n305), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n206), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n262), .B2(new_n484), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n250), .B1(new_n248), .B2(new_n370), .ZN(new_n520));
  INV_X1    g0320(.A(new_n481), .ZN(new_n521));
  INV_X1    g0321(.A(new_n370), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n511), .A2(new_n513), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(KEYINPUT84), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n510), .A2(G200), .ZN(new_n528));
  AOI211_X1 g0328(.A(new_n289), .B(new_n508), .C1(new_n276), .C2(new_n503), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(KEYINPUT85), .A3(G87), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT85), .ZN(new_n531));
  INV_X1    g0331(.A(G87), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n481), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n520), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g0337(.A(KEYINPUT88), .B(G294), .Z(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G33), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n269), .A2(G250), .A3(new_n272), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n276), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n475), .A2(new_n281), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n474), .A2(G264), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n294), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n542), .A2(new_n276), .B1(G264), .B2(new_n474), .ZN(new_n548));
  INV_X1    g0348(.A(G179), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(new_n544), .ZN(new_n550));
  INV_X1    g0350(.A(new_n250), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n269), .A2(new_n209), .A3(G87), .ZN(new_n552));
  AND2_X1   g0352(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT87), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n557), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT23), .ZN(new_n560));
  INV_X1    g0360(.A(G107), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(G20), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n269), .A2(new_n209), .A3(G87), .A4(new_n553), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n556), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n563), .A2(new_n566), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n564), .A4(new_n556), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n551), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT25), .B1(new_n248), .B2(new_n561), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n561), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n574), .A2(new_n575), .B1(G107), .B2(new_n521), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n547), .B(new_n550), .C1(new_n572), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n568), .A2(new_n571), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n250), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n548), .A2(G190), .A3(new_n544), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n546), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n580), .A2(new_n576), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n269), .A2(G244), .A3(new_n272), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(KEYINPUT4), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n269), .A2(new_n588), .A3(G244), .A4(new_n272), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n483), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n276), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n474), .A2(G257), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n544), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n595), .A3(new_n296), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n597), .A2(new_n484), .A3(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(G97), .B(G107), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n600), .A2(new_n209), .B1(new_n271), .B2(new_n260), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n561), .B1(new_n430), .B2(new_n431), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n250), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n247), .A2(G97), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n521), .B2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n594), .B1(new_n276), .B2(new_n591), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n596), .B(new_n606), .C1(new_n607), .C2(G169), .ZN(new_n608));
  INV_X1    g0408(.A(new_n605), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n484), .A2(new_n561), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n597), .B1(new_n610), .B2(new_n205), .ZN(new_n611));
  INV_X1    g0411(.A(new_n598), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n430), .A2(new_n431), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n561), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n609), .B1(new_n616), .B2(new_n250), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n592), .A2(new_n595), .A3(G190), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n618), .C1(new_n407), .C2(new_n607), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n578), .A2(new_n583), .A3(new_n608), .A4(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n465), .A2(new_n499), .A3(new_n537), .A4(new_n620), .ZN(G372));
  AOI21_X1  g0421(.A(new_n339), .B1(new_n324), .B2(new_n327), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n344), .B2(new_n381), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n443), .A2(new_n461), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n454), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n293), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n298), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(new_n608), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n537), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n296), .B(new_n508), .C1(new_n276), .C2(new_n503), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n294), .B1(new_n504), .B2(new_n509), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n524), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n592), .A2(new_n595), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n635), .A2(new_n294), .B1(new_n603), .B2(new_n605), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n512), .A2(G190), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n528), .A2(new_n637), .A3(new_n520), .A4(new_n534), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n636), .A2(new_n638), .A3(new_n596), .A4(new_n634), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n634), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n631), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n577), .B1(new_n579), .B2(new_n250), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n547), .A2(new_n550), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT89), .B1(new_n644), .B2(new_n494), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n638), .A2(new_n634), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n582), .A2(new_n581), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n619), .A2(new_n608), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n493), .A2(new_n492), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT89), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n578), .A2(new_n650), .A3(new_n651), .A4(new_n491), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n645), .A2(new_n648), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n628), .B1(new_n464), .B2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(G213), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n488), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n494), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n498), .B2(new_n662), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n661), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT90), .B1(new_n642), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n668), .B(new_n661), .C1(new_n572), .C2(new_n577), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n578), .A3(new_n583), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n644), .A2(new_n661), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n578), .A2(new_n661), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n583), .A2(new_n578), .A3(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n580), .A2(new_n576), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n676), .B2(new_n661), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n494), .A2(new_n666), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n674), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n212), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n208), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n685), .A2(new_n686), .B1(new_n216), .B2(new_n684), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT28), .Z(new_n688));
  INV_X1    g0488(.A(new_n646), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n630), .A3(new_n690), .A4(KEYINPUT26), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n689), .A2(new_n583), .A3(new_n608), .A4(new_n619), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n644), .A2(new_n494), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n691), .B(new_n634), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT26), .B1(new_n537), .B2(new_n630), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT92), .B1(new_n639), .B2(new_n629), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT29), .B(new_n666), .C1(new_n694), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n661), .B1(new_n641), .B2(new_n653), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(KEYINPUT29), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n499), .A2(new_n537), .A3(new_n620), .A4(new_n666), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n548), .A2(new_n512), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n470), .A2(new_n476), .A3(G179), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n705), .A3(KEYINPUT30), .A4(new_n607), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n297), .B1(new_n470), .B2(new_n476), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n635), .A2(new_n510), .A3(new_n546), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n592), .A2(new_n595), .A3(new_n512), .A4(new_n548), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n704), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT91), .B(new_n710), .C1(new_n711), .C2(new_n704), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n702), .B1(new_n716), .B2(new_n666), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n706), .A3(new_n708), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n701), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n700), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n688), .B1(new_n723), .B2(G1), .ZN(G364));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(G45), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n685), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n217), .B1(G20), .B2(new_n294), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n212), .A2(new_n269), .ZN(new_n741));
  INV_X1    g0541(.A(G355), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n212), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n683), .A2(new_n269), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n471), .B2(new_n216), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n242), .A2(new_n471), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n734), .B1(new_n740), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n407), .A2(G179), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n209), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(new_n289), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n750), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n269), .B1(new_n752), .B2(new_n561), .C1(new_n532), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n297), .A2(G20), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n296), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n753), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n758), .A2(new_n202), .B1(new_n201), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(new_n289), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n755), .B(new_n761), .C1(G50), .C2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(KEYINPUT97), .A2(G179), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT97), .B1(G179), .B2(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n289), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n209), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G97), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT96), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n759), .A2(new_n771), .A3(new_n751), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(new_n759), .B2(new_n751), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G77), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n209), .B(G190), .C1(new_n765), .C2(new_n766), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G159), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT32), .Z(new_n779));
  NAND4_X1  g0579(.A1(new_n763), .A2(new_n770), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n762), .B(KEYINPUT98), .Z(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G326), .ZN(new_n783));
  INV_X1    g0583(.A(new_n754), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n269), .B1(new_n784), .B2(G303), .ZN(new_n785));
  INV_X1    g0585(.A(G322), .ZN(new_n786));
  XOR2_X1   g0586(.A(KEYINPUT33), .B(G317), .Z(new_n787));
  OAI221_X1 g0587(.A(new_n785), .B1(new_n786), .B2(new_n760), .C1(new_n758), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n538), .B2(new_n769), .ZN(new_n789));
  INV_X1    g0589(.A(new_n752), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n777), .A2(G329), .B1(new_n790), .B2(G283), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n775), .A2(G311), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n783), .A2(new_n789), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n780), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n749), .B1(new_n795), .B2(new_n738), .ZN(new_n796));
  INV_X1    g0596(.A(new_n737), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n796), .B1(new_n664), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT100), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n664), .A2(G330), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n664), .A2(G330), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n733), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n799), .B1(new_n801), .B2(new_n803), .ZN(G396));
  XNOR2_X1  g0604(.A(new_n372), .B(new_n373), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n666), .B1(new_n805), .B2(new_n361), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n380), .B1(new_n377), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n376), .A2(new_n378), .A3(new_n379), .A4(new_n666), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n699), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n733), .B1(new_n811), .B2(new_n721), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n721), .C2(new_n811), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n738), .A2(new_n735), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n733), .B1(new_n271), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n810), .A2(new_n736), .ZN(new_n819));
  INV_X1    g0619(.A(new_n762), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n760), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G283), .B2(new_n757), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n775), .A2(G116), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n350), .B1(new_n752), .B2(new_n532), .C1(new_n561), .C2(new_n754), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G311), .B2(new_n777), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n770), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n350), .B1(new_n790), .B2(G68), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n333), .B2(new_n754), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G132), .B2(new_n777), .ZN(new_n831));
  INV_X1    g0631(.A(new_n760), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n762), .A2(G137), .B1(new_n832), .B2(G143), .ZN(new_n833));
  INV_X1    g0633(.A(G159), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n258), .B2(new_n758), .C1(new_n774), .C2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n831), .B1(new_n201), .B2(new_n768), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n828), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT101), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n738), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n818), .B(new_n819), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n815), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  NOR2_X1   g0647(.A1(new_n727), .A2(new_n208), .ZN(new_n848));
  INV_X1    g0648(.A(G330), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n850));
  OR3_X1    g0650(.A1(new_n716), .A2(new_n702), .A3(new_n666), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT105), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n852), .B(new_n702), .C1(new_n716), .C2(new_n666), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n850), .A2(new_n701), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n339), .A2(new_n666), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n341), .B2(new_n344), .ZN(new_n857));
  INV_X1    g0657(.A(new_n344), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n622), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n810), .B(new_n854), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n422), .A2(new_n425), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(new_n424), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n659), .B1(new_n863), .B2(new_n447), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n462), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n448), .A2(new_n451), .ZN(new_n868));
  INV_X1    g0668(.A(new_n659), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n448), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n411), .A2(new_n440), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n867), .A2(new_n868), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n863), .A2(new_n447), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n451), .B2(new_n869), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n867), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n866), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n871), .A2(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n868), .A2(new_n870), .A3(new_n871), .A4(new_n867), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n879), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT104), .B1(new_n878), .B2(new_n879), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n885), .B2(new_n865), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n861), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(new_n867), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n441), .A2(new_n442), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n870), .B1(new_n454), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n890), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n881), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n860), .A2(new_n888), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n465), .A2(new_n854), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n849), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n462), .A2(new_n864), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n876), .A2(new_n880), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n890), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n341), .A2(new_n661), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n454), .A2(new_n869), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n907), .A2(new_n881), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n341), .A2(new_n344), .A3(new_n856), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n855), .B1(new_n622), .B2(new_n858), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n699), .A2(new_n810), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n808), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n661), .B(new_n809), .C1(new_n641), .C2(new_n653), .ZN(new_n920));
  INV_X1    g0720(.A(new_n808), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT103), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n916), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n911), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n382), .A2(new_n463), .A3(new_n926), .A4(new_n698), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n628), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n925), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n848), .B1(new_n902), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n929), .B2(new_n902), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n613), .A2(KEYINPUT35), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n613), .A2(KEYINPUT35), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n932), .A2(G116), .A3(new_n218), .A4(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT36), .ZN(new_n935));
  OAI21_X1  g0735(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n215), .A2(new_n936), .B1(G50), .B2(new_n202), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(G1), .A3(new_n725), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n935), .A3(new_n938), .ZN(G367));
  NOR2_X1   g0739(.A1(new_n731), .A2(new_n208), .ZN(new_n940));
  INV_X1    g0740(.A(new_n673), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n606), .A2(new_n661), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n619), .A2(new_n608), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n630), .A2(new_n661), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n619), .A2(KEYINPUT107), .A3(new_n608), .A4(new_n942), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT44), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n681), .A2(new_n948), .B1(KEYINPUT110), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n670), .A2(new_n679), .B1(new_n578), .B2(new_n661), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(KEYINPUT110), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n949), .A2(KEYINPUT110), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT109), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n681), .A2(new_n958), .A3(new_n948), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT45), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT45), .B1(new_n957), .B2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n941), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n964), .A2(new_n673), .A3(new_n956), .A4(new_n960), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n671), .B(new_n679), .C1(new_n675), .C2(new_n677), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT111), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n678), .A2(new_n680), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n670), .A2(KEYINPUT111), .A3(new_n679), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n802), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n966), .A2(new_n967), .B1(new_n678), .B2(new_n680), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n665), .B1(new_n974), .B2(new_n971), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n976), .A2(new_n721), .A3(new_n700), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n963), .A2(new_n965), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n963), .A2(new_n965), .A3(new_n977), .A4(KEYINPUT112), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n722), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n684), .B(new_n983), .Z(new_n984));
  OAI21_X1  g0784(.A(new_n940), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n951), .A2(new_n969), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT42), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n578), .B1(new_n945), .B2(new_n947), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n666), .B1(new_n988), .B2(new_n630), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n535), .A2(new_n661), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n689), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n634), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n993), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(KEYINPUT43), .B2(new_n993), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n990), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n987), .A2(new_n989), .A3(new_n997), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n673), .A2(new_n951), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n985), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n744), .A2(new_n238), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n740), .B1(new_n683), .B2(new_n522), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n733), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n782), .A2(G143), .B1(G50), .B2(new_n775), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n269), .B1(new_n752), .B2(new_n271), .C1(new_n201), .C2(new_n754), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n758), .A2(new_n834), .B1(new_n258), .B2(new_n760), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G137), .C2(new_n777), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1008), .B(new_n1011), .C1(new_n202), .C2(new_n768), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n782), .A2(G311), .B1(G303), .B2(new_n832), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT113), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n784), .A2(G116), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n757), .A2(new_n538), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n561), .C2(new_n768), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n777), .A2(G317), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n350), .C1(new_n484), .C2(new_n752), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT114), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1021), .A2(new_n1022), .B1(new_n775), .B2(G283), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1015), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1012), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n1007), .B1(new_n797), .B2(new_n993), .C1(new_n1029), .C2(new_n843), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1004), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n366), .A2(new_n368), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n333), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1034), .A2(new_n686), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1032), .B2(new_n333), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n744), .B1(new_n1036), .B2(new_n1037), .C1(new_n235), .C2(new_n471), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(G107), .B2(new_n212), .C1(new_n686), .C2(new_n741), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n733), .B1(new_n1039), .B2(new_n739), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n672), .B2(new_n797), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n757), .A2(G311), .B1(new_n832), .B2(G317), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n821), .B2(new_n774), .C1(new_n781), .C2(new_n786), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n769), .A2(G283), .B1(new_n538), .B2(new_n784), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n350), .B1(new_n752), .B2(new_n478), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n777), .B2(G326), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n774), .A2(new_n202), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n758), .A2(new_n261), .B1(new_n333), .B2(new_n760), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G159), .B2(new_n762), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n769), .A2(new_n522), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n784), .A2(G77), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n269), .C1(new_n484), .C2(new_n752), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G150), .B2(new_n777), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1054), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1041), .B1(new_n1063), .B2(new_n738), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n940), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n976), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n977), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n684), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n723), .A2(new_n976), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n980), .A2(new_n981), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n684), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n963), .A2(new_n965), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n1067), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n963), .A2(new_n965), .A3(new_n1065), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n948), .A2(new_n797), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT116), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n350), .B1(new_n790), .B2(G87), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n202), .B2(new_n754), .C1(new_n758), .C2(new_n333), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G143), .B2(new_n777), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n775), .A2(new_n1032), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n769), .A2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n762), .A2(G150), .B1(new_n832), .B2(G159), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n777), .A2(G322), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n350), .B1(new_n752), .B2(new_n561), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G283), .B2(new_n784), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(new_n758), .C2(new_n821), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G116), .B2(new_n769), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n822), .B2(new_n774), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n762), .A2(G317), .B1(new_n832), .B2(G311), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1084), .A2(new_n1086), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n738), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n739), .B1(new_n484), .B2(new_n212), .C1(new_n745), .C2(new_n245), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1078), .A2(new_n734), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1076), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1075), .A2(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n922), .A2(new_n919), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n909), .B1(new_n1102), .B2(new_n915), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT39), .B1(new_n881), .B2(new_n895), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n666), .B(new_n807), .C1(new_n694), .C2(new_n697), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n808), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n909), .B1(new_n915), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n896), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n721), .A2(new_n809), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n915), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1107), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n915), .A2(new_n810), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n854), .A2(G330), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1103), .B1(new_n904), .B2(new_n908), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1111), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1114), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n382), .A2(G330), .A3(new_n463), .A4(new_n854), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n628), .A2(new_n927), .A3(new_n1122), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1115), .A2(new_n1116), .B1(new_n1112), .B2(new_n915), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1109), .B1(new_n1112), .B2(new_n915), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n916), .B1(new_n1116), .B2(new_n809), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1124), .A2(new_n1102), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1121), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1114), .A2(new_n1120), .A3(new_n1128), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n684), .A3(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1114), .A2(new_n1120), .A3(new_n1065), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n735), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n733), .B1(new_n261), .B2(new_n816), .ZN(new_n1135));
  INV_X1    g0935(.A(G137), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n269), .B1(new_n333), .B2(new_n752), .C1(new_n758), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G159), .B2(new_n769), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n775), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n784), .A2(G150), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G128), .B2(new_n762), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n832), .A2(G132), .B1(new_n777), .B2(G125), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1138), .A2(new_n1141), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(G283), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n820), .A2(new_n1147), .B1(new_n478), .B2(new_n760), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G107), .B2(new_n757), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n775), .A2(G97), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n350), .B1(new_n752), .B2(new_n202), .C1(new_n532), .C2(new_n754), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G294), .B2(new_n777), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1149), .A2(new_n1083), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1134), .B(new_n1135), .C1(new_n843), .C2(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1132), .A2(new_n1156), .ZN(G378));
  AND2_X1   g0957(.A1(new_n910), .A2(new_n924), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n267), .A2(new_n869), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n299), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n299), .A2(new_n1162), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1165), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1167), .A2(new_n1163), .A3(new_n1159), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT40), .B1(new_n912), .B2(new_n861), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n898), .A2(G330), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n849), .B1(new_n896), .B2(new_n897), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n860), .B1(new_n907), .B2(new_n881), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1169), .B(new_n1174), .C1(KEYINPUT40), .C2(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1158), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1173), .A2(new_n1176), .B1(new_n910), .B2(new_n924), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1123), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1131), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n684), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1176), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1169), .B1(new_n889), .B2(new_n1174), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n925), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1158), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1131), .A2(new_n1180), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1182), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1170), .A2(new_n735), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n816), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n734), .B1(G50), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n269), .A2(G41), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1194), .C1(new_n283), .C2(new_n284), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n820), .A2(new_n478), .B1(new_n561), .B2(new_n760), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G97), .B2(new_n757), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1059), .B(new_n1194), .C1(new_n201), .C2(new_n752), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n768), .A2(new_n202), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(G283), .C2(new_n777), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(new_n370), .C2(new_n774), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT58), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n762), .A2(G125), .B1(new_n832), .B2(G128), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n757), .A2(G132), .B1(new_n784), .B2(new_n1140), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1136), .B2(new_n774), .C1(new_n258), .C2(new_n768), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n283), .B(new_n284), .C1(new_n752), .C2(new_n834), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n777), .B2(G124), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1207), .A2(KEYINPUT59), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1203), .B1(new_n1202), .B2(new_n1201), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1193), .B1(new_n1213), .B2(new_n738), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1191), .A2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1187), .B2(new_n1065), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1216), .ZN(G375));
  INV_X1    g1017(.A(new_n984), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1129), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1127), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n916), .A2(new_n735), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n734), .B1(G68), .B2(new_n1192), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G132), .A2(new_n762), .B1(new_n757), .B2(new_n1140), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1136), .B2(new_n760), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT118), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n775), .A2(G150), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n777), .A2(G128), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n350), .B1(new_n790), .B2(G58), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n834), .C2(new_n754), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G50), .B2(new_n769), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .A4(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n350), .B1(new_n752), .B2(new_n271), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n820), .A2(new_n822), .B1(new_n1147), .B2(new_n760), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(G116), .C2(new_n757), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1237), .B(new_n1058), .C1(new_n561), .C2(new_n774), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n777), .A2(G303), .B1(G97), .B2(new_n784), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT117), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1234), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1223), .B1(new_n1241), .B2(new_n738), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1221), .A2(new_n1065), .B1(new_n1222), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1220), .A2(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(G375), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1030), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n985), .B2(new_n1003), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G393), .A2(G396), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n846), .A2(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G381), .A3(G390), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1245), .A2(new_n1247), .A3(new_n1248), .A4(new_n1251), .ZN(G407));
  NAND2_X1  g1052(.A1(new_n660), .A2(G213), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1245), .A2(new_n1248), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  INV_X1    g1056(.A(KEYINPUT124), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1187), .A2(new_n1188), .A3(new_n1218), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1215), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1185), .A2(KEYINPUT119), .A3(new_n1186), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1065), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT119), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1258), .B(new_n1259), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1248), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1216), .C1(new_n1182), .C2(new_n1189), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1219), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1129), .B(KEYINPUT120), .C1(new_n1267), .C2(KEYINPUT60), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT120), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT60), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1128), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1072), .B1(new_n1267), .B2(KEYINPUT60), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1243), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n846), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1273), .A2(G384), .A3(new_n1243), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1266), .A2(KEYINPUT63), .A3(new_n1253), .A4(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1254), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1277), .B(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1254), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1279), .B(new_n1280), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G387), .B(G390), .ZN(new_n1286));
  AND2_X1   g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1287), .A2(new_n1249), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1288), .B1(new_n1247), .B2(G390), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT121), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G390), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1075), .A2(KEYINPUT121), .A3(new_n1100), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT122), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(new_n1296), .A2(new_n1297), .A3(new_n1247), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT121), .B1(new_n1075), .B2(new_n1100), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n1293), .B(new_n1099), .C1(new_n1071), .C2(new_n1074), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT122), .B1(G387), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1292), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT123), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1297), .B1(new_n1296), .B2(new_n1247), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G387), .A2(new_n1301), .A3(KEYINPUT122), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT123), .B1(new_n1308), .B2(new_n1292), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1291), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1254), .B(new_n1277), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1310), .B1(new_n1311), .B2(KEYINPUT63), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1257), .B1(new_n1285), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(KEYINPUT123), .A3(new_n1292), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1290), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1266), .A2(new_n1253), .A3(new_n1278), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1284), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1277), .B(new_n1281), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1319), .A2(KEYINPUT124), .A3(new_n1322), .A4(new_n1279), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1322), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1326), .B(KEYINPUT62), .C1(new_n1284), .C2(new_n1278), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT125), .B1(new_n1318), .B2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1266), .A2(KEYINPUT62), .A3(new_n1253), .A4(new_n1278), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT126), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1284), .A2(new_n1333), .A3(KEYINPUT62), .A4(new_n1278), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1325), .B1(new_n1330), .B2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1324), .B1(new_n1336), .B2(new_n1310), .ZN(G405));
  NAND2_X1  g1137(.A1(G375), .A2(new_n1248), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1265), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1338), .A2(KEYINPUT127), .A3(new_n1265), .A4(new_n1278), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1310), .ZN(G402));
endmodule


