//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT76), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n187), .A2(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n191), .A2(KEYINPUT76), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n193), .B2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(G104), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n188), .B2(new_n190), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n197), .B1(new_n195), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(new_n205), .A3(KEYINPUT4), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(G113), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(KEYINPUT2), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n208), .B(new_n210), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n210), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n217), .A3(KEYINPUT67), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n217), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(G101), .C1(new_n193), .C2(new_n198), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n206), .A2(new_n218), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n188), .B2(new_n200), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n205), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n214), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT5), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(new_n211), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n232), .A3(new_n234), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT6), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G125), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT71), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(new_n248), .B2(G143), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G146), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n249), .A2(new_n252), .B1(G143), .B2(new_n248), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n241), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n242), .B(new_n247), .C1(new_n253), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n248), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(G146), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n250), .B1(new_n251), .B2(G146), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n248), .A2(KEYINPUT64), .A3(G143), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n258), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n262), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n257), .B1(new_n268), .B2(new_n247), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G224), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n269), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n233), .A2(new_n273), .A3(new_n235), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n238), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n276), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n257), .B(new_n278), .C1(new_n268), .C2(new_n247), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n237), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n234), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n228), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT80), .A4(KEYINPUT5), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n230), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n287), .A2(new_n214), .A3(new_n205), .A4(new_n225), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n288), .A2(KEYINPUT81), .B1(new_n226), .B2(new_n231), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n288), .A2(KEYINPUT81), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n281), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n275), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n293), .B(KEYINPUT82), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n275), .B2(new_n292), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G214), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(G221), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n239), .A2(new_n259), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n312), .A2(G128), .B1(new_n260), .B2(new_n261), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n266), .A2(new_n239), .A3(KEYINPUT77), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n205), .B(new_n225), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n205), .A2(new_n225), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n268), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT11), .A2(G134), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(G137), .ZN(new_n323));
  INV_X1    g137(.A(G137), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OR2_X1    g140(.A1(KEYINPUT65), .A2(G134), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT65), .A2(G134), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G137), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(G137), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n326), .B(new_n329), .C1(new_n330), .C2(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G131), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT65), .A2(G134), .ZN(new_n333));
  NOR2_X1   g147(.A1(KEYINPUT65), .A2(G134), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n326), .A4(new_n329), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT12), .B1(new_n320), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n310), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n320), .A2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT12), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n340), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT78), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n317), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n311), .B1(new_n253), .B2(new_n266), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n351), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n333), .A2(new_n334), .A3(new_n324), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n336), .B2(new_n335), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n338), .B1(new_n354), .B2(new_n326), .ZN(new_n355));
  INV_X1    g169(.A(new_n339), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n242), .B1(new_n253), .B2(new_n256), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n206), .A2(new_n359), .A3(new_n223), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n350), .A2(new_n352), .A3(new_n357), .A4(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G140), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n270), .A2(G227), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n343), .A2(new_n348), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n350), .A2(new_n360), .A3(new_n352), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n340), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n361), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G469), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n307), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n307), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n361), .B1(new_n341), .B2(new_n342), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n377), .A2(new_n364), .B1(new_n366), .B2(new_n369), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n378), .B2(G469), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n309), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT16), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n245), .A2(G125), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n243), .A2(KEYINPUT71), .ZN(new_n383));
  OAI21_X1  g197(.A(G140), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(G125), .A2(G140), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n381), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n244), .B2(new_n246), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n248), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n244), .B2(new_n246), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT16), .B1(new_n392), .B2(new_n385), .ZN(new_n393));
  INV_X1    g207(.A(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(G146), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G237), .A2(G953), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n251), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(G143), .A3(G214), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT17), .A3(G131), .ZN(new_n401));
  INV_X1    g215(.A(new_n399), .ZN(new_n402));
  AOI21_X1  g216(.A(G143), .B1(new_n396), .B2(G214), .ZN(new_n403));
  OAI21_X1  g217(.A(G131), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n338), .A3(new_n399), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n391), .A2(new_n395), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n187), .ZN(new_n410));
  XNOR2_X1  g224(.A(G125), .B(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n248), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT71), .B(G125), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n386), .B1(new_n413), .B2(new_n388), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(new_n248), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n400), .A2(KEYINPUT18), .A3(G131), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT18), .A2(G131), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n398), .A2(new_n399), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n408), .A2(new_n410), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n410), .B1(new_n408), .B2(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n307), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G475), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n410), .A3(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n404), .A2(new_n405), .ZN(new_n426));
  OAI211_X1 g240(.A(KEYINPUT19), .B(new_n386), .C1(new_n413), .C2(new_n388), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n411), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n248), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n395), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n419), .ZN(new_n432));
  INV_X1    g246(.A(new_n410), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(G475), .A2(G902), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT83), .Z(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n424), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g253(.A(KEYINPUT20), .B(new_n437), .C1(new_n425), .C2(new_n434), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n423), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT85), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n209), .B2(G122), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT84), .A3(G116), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n209), .A2(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n447), .A2(KEYINPUT14), .A3(G116), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G107), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n251), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n258), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n334), .B2(new_n333), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n333), .A2(new_n334), .ZN(new_n459));
  XNOR2_X1  g273(.A(G128), .B(G143), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n449), .A2(new_n196), .A3(new_n450), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G134), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n258), .A2(G143), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT13), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT13), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n468), .A2(new_n469), .B1(new_n459), .B2(new_n460), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n449), .A2(new_n196), .A3(new_n450), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n196), .B1(new_n449), .B2(new_n450), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n270), .A2(G217), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n304), .A2(new_n305), .A3(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n464), .B2(new_n473), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n307), .B(new_n444), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(new_n473), .ZN(new_n480));
  INV_X1    g294(.A(new_n475), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n478), .B(new_n479), .C1(new_n484), .C2(new_n443), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(KEYINPUT86), .A3(new_n444), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n270), .A2(G952), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(G234), .B2(G237), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n307), .B(new_n270), .C1(G234), .C2(G237), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(G898), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g307(.A1(new_n441), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n301), .A2(new_n380), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G217), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(G234), .B2(new_n307), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT22), .B(G137), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n270), .A2(G221), .A3(G234), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n207), .B2(G128), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(new_n503), .C1(G119), .C2(new_n258), .ZN(new_n504));
  XNOR2_X1  g318(.A(G119), .B(G128), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT24), .B(G110), .Z(new_n506));
  AOI22_X1  g320(.A1(new_n504), .A2(G110), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n248), .B(new_n390), .C1(new_n414), .C2(KEYINPUT16), .ZN(new_n508));
  AOI21_X1  g322(.A(G146), .B1(new_n393), .B2(new_n394), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n504), .A2(G110), .B1(new_n505), .B2(new_n506), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n395), .A2(new_n412), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n500), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  INV_X1    g332(.A(new_n500), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n518), .B(new_n519), .C1(new_n511), .C2(new_n513), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT25), .B1(new_n521), .B2(new_n307), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n517), .A2(new_n520), .A3(new_n523), .A4(G902), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n497), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n497), .A2(G902), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n391), .A2(new_n395), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n512), .B1(new_n528), .B2(new_n507), .ZN(new_n529));
  INV_X1    g343(.A(new_n513), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n516), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n519), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n518), .B1(new_n511), .B2(new_n513), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n500), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n532), .A2(KEYINPUT73), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n526), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  INV_X1    g352(.A(new_n218), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT67), .B1(new_n214), .B2(new_n217), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n324), .A2(G134), .ZN(new_n544));
  OAI21_X1  g358(.A(G131), .B1(new_n330), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n339), .A2(new_n351), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n542), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n358), .B1(new_n332), .B2(new_n339), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n339), .A2(new_n351), .A3(new_n545), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT30), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n541), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT69), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n548), .A2(new_n549), .A3(new_n541), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n396), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n552), .B1(new_n553), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n221), .A2(new_n218), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n543), .A2(new_n561), .A3(new_n546), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(KEYINPUT69), .A3(new_n558), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n551), .A2(new_n560), .A3(KEYINPUT31), .A4(new_n563), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n569), .B1(new_n562), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n553), .A2(KEYINPUT28), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n559), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT70), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT70), .B(new_n559), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n538), .B1(new_n568), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT32), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n566), .A2(new_n567), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n575), .A3(new_n576), .ZN(new_n582));
  INV_X1    g396(.A(new_n538), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n579), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n543), .A2(new_n542), .A3(new_n546), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT30), .B1(new_n548), .B2(new_n549), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n559), .B1(new_n587), .B2(new_n553), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n561), .B1(new_n543), .B2(new_n546), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT28), .B1(new_n590), .B2(new_n553), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n562), .A2(new_n569), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n588), .B(new_n589), .C1(new_n593), .C2(new_n559), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n591), .A2(KEYINPUT29), .A3(new_n558), .A4(new_n592), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n307), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n582), .A2(new_n584), .B1(new_n596), .B2(G472), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT74), .B(new_n537), .C1(new_n580), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT74), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n584), .B1(new_n568), .B2(new_n577), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n596), .A2(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT70), .B1(new_n593), .B2(new_n559), .ZN(new_n602));
  INV_X1    g416(.A(new_n576), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n583), .B1(new_n604), .B2(new_n581), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n600), .B(new_n601), .C1(new_n605), .C2(KEYINPUT32), .ZN(new_n606));
  INV_X1    g420(.A(new_n537), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n599), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n495), .B1(new_n598), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n582), .B2(new_n307), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n605), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n607), .A3(new_n380), .ZN(new_n614));
  XOR2_X1   g428(.A(new_n614), .B(KEYINPUT87), .Z(new_n615));
  NAND2_X1  g429(.A1(new_n275), .A2(new_n292), .ZN(new_n616));
  INV_X1    g430(.A(new_n293), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n275), .A2(new_n292), .A3(new_n293), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n299), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n482), .B2(KEYINPUT88), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n476), .B2(new_n477), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n482), .B(new_n483), .C1(KEYINPUT88), .C2(new_n622), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(G478), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n442), .A2(new_n307), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n484), .B2(new_n442), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n493), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n441), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT34), .B(G104), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  AOI21_X1  g450(.A(new_n300), .B1(new_n618), .B2(new_n619), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n435), .A2(new_n438), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT20), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n435), .A2(new_n424), .A3(new_n438), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(KEYINPUT89), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT89), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n439), .B2(new_n440), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n493), .B(KEYINPUT90), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n487), .B1(G475), .B2(new_n422), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n637), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n615), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT91), .ZN(new_n651));
  INV_X1    g465(.A(new_n497), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n521), .A2(KEYINPUT25), .A3(new_n307), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n532), .A2(new_n307), .A3(new_n534), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n523), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n533), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n526), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n651), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n525), .A2(KEYINPUT91), .A3(new_n660), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n495), .A3(new_n613), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT92), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n600), .A2(new_n601), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT32), .B1(new_n582), .B2(new_n538), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n380), .B(new_n637), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT93), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n491), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n490), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n644), .A2(new_n646), .A3(new_n672), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n641), .A2(new_n643), .A3(new_n676), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n488), .A2(new_n423), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT93), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n662), .A2(new_n663), .A3(new_n677), .A4(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT94), .B1(new_n671), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n375), .A2(new_n379), .ZN(new_n683));
  INV_X1    g497(.A(new_n309), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n637), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n580), .B2(new_n597), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT94), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n677), .A2(new_n680), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n687), .A3(new_n664), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XNOR2_X1  g506(.A(new_n676), .B(KEYINPUT39), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n380), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  AND2_X1   g509(.A1(new_n695), .A2(KEYINPUT96), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(KEYINPUT96), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n559), .B1(new_n590), .B2(new_n553), .ZN(new_n698));
  OR2_X1    g512(.A1(new_n698), .A2(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(KEYINPUT95), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n699), .A2(new_n564), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n611), .B1(new_n701), .B2(new_n307), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n582), .B2(new_n584), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n580), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n298), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n616), .A2(new_n295), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n619), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT38), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n653), .A2(new_n655), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n661), .B1(new_n712), .B2(new_n497), .ZN(new_n713));
  INV_X1    g527(.A(new_n441), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n487), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n299), .A3(new_n715), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n705), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n696), .A2(new_n697), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT97), .B(G143), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G45));
  NAND2_X1  g534(.A1(new_n630), .A2(new_n441), .ZN(new_n721));
  INV_X1    g535(.A(new_n676), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n662), .A2(new_n663), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n671), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n248), .ZN(G48));
  AOI21_X1  g540(.A(new_n374), .B1(new_n373), .B2(new_n307), .ZN(new_n727));
  AOI211_X1 g541(.A(G469), .B(G902), .C1(new_n367), .C2(new_n372), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n309), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n606), .A2(new_n607), .A3(new_n633), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT98), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n537), .B1(new_n580), .B2(new_n597), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT98), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n633), .A4(new_n729), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NAND3_X1  g551(.A1(new_n732), .A2(new_n647), .A3(new_n729), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  NAND2_X1  g553(.A1(new_n373), .A2(new_n307), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(G469), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n684), .A3(new_n375), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n621), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n664), .A2(new_n606), .A3(new_n494), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT99), .B(G119), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G21));
  AOI21_X1  g560(.A(new_n583), .B1(new_n581), .B2(new_n573), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n612), .A2(new_n537), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n637), .A2(new_n715), .ZN(new_n749));
  INV_X1    g563(.A(new_n645), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n742), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT100), .B(G122), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G24));
  INV_X1    g568(.A(KEYINPUT101), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n582), .A2(new_n307), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G472), .ZN(new_n757));
  INV_X1    g571(.A(new_n713), .ZN(new_n758));
  INV_X1    g572(.A(new_n747), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n729), .A2(new_n637), .A3(new_n723), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n755), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n612), .A2(new_n713), .A3(new_n747), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(KEYINPUT101), .A3(new_n723), .A4(new_n743), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n607), .B1(new_n669), .B2(new_n670), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n377), .A2(new_n364), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT102), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n366), .A2(new_n770), .A3(new_n369), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n366), .B2(new_n369), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n769), .B(G469), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n376), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n375), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n309), .A2(new_n300), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n708), .A2(new_n619), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n723), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n767), .B1(new_n768), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n781), .B1(new_n780), .B2(new_n783), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  NAND4_X1  g601(.A1(new_n677), .A2(new_n680), .A3(new_n776), .A4(new_n778), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT104), .B1(new_n768), .B2(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n677), .A2(new_n680), .A3(new_n776), .A4(new_n778), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT104), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n732), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(KEYINPUT43), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n630), .A2(new_n714), .A3(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n795), .A2(KEYINPUT43), .ZN(new_n799));
  OAI22_X1  g613(.A1(new_n629), .A2(new_n441), .B1(new_n799), .B2(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n758), .B(new_n801), .C1(new_n612), .C2(new_n605), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT44), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(KEYINPUT108), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n294), .A2(new_n297), .A3(new_n300), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n803), .B2(KEYINPUT44), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n805), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n361), .A2(new_n365), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT102), .B1(new_n370), .B2(new_n812), .ZN(new_n813));
  AOI221_X4 g627(.A(new_n811), .B1(new_n364), .B2(new_n377), .C1(new_n813), .C2(new_n771), .ZN(new_n814));
  OAI21_X1  g628(.A(G469), .B1(new_n378), .B2(KEYINPUT45), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT46), .B(new_n775), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT105), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n375), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n769), .B1(new_n370), .B2(new_n812), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n374), .B1(new_n819), .B2(new_n811), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n769), .B(KEYINPUT45), .C1(new_n772), .C2(new_n773), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n376), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT105), .B1(new_n822), .B2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT106), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n816), .A2(new_n817), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT106), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n825), .A2(new_n826), .A3(new_n827), .A4(new_n375), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n822), .A2(KEYINPUT46), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n684), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n693), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n810), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT109), .B(G137), .Z(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(G39));
  AND3_X1   g651(.A1(new_n830), .A2(KEYINPUT47), .A3(new_n684), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT47), .B1(new_n830), .B2(new_n684), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n537), .A2(new_n723), .A3(new_n807), .ZN(new_n841));
  OR3_X1    g655(.A1(new_n840), .A2(new_n606), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G140), .ZN(G42));
  NAND2_X1  g657(.A1(new_n741), .A2(new_n375), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT110), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT49), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n607), .A2(new_n714), .A3(new_n630), .A4(new_n777), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n705), .A3(new_n711), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n713), .A2(new_n684), .A3(new_n676), .ZN(new_n850));
  INV_X1    g664(.A(new_n776), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n851), .A3(new_n749), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n852), .B2(new_n704), .ZN(new_n853));
  INV_X1    g667(.A(new_n725), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n691), .A2(new_n765), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n725), .B1(new_n682), .B2(new_n690), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n765), .A4(new_n853), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n852), .A2(new_n704), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n691), .A2(new_n765), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n485), .A2(new_n486), .B1(new_n422), .B2(G475), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n641), .A2(new_n643), .A3(new_n866), .A4(new_n676), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n683), .A2(new_n807), .A3(new_n867), .A4(new_n684), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n580), .B2(new_n597), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n869), .A2(new_n664), .B1(new_n763), .B2(new_n782), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT112), .B1(new_n793), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n786), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n744), .A2(new_n738), .A3(new_n752), .A4(new_n665), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n441), .A2(new_n487), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n301), .A2(KEYINPUT111), .A3(new_n645), .A4(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n709), .A2(new_n299), .A3(new_n645), .ZN(new_n879));
  INV_X1    g693(.A(new_n876), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n877), .B(new_n881), .C1(new_n721), .C2(new_n879), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(new_n607), .A3(new_n380), .A4(new_n613), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n875), .A2(new_n609), .A3(new_n735), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n865), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n862), .B(KEYINPUT52), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n768), .A2(KEYINPUT104), .A3(new_n788), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n791), .B1(new_n732), .B2(new_n790), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n870), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n870), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n609), .A2(new_n883), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n731), .A2(new_n734), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n874), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n898), .A3(new_n786), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT53), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n887), .A2(new_n900), .A3(KEYINPUT54), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n886), .B1(new_n888), .B2(new_n899), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n886), .B1(new_n780), .B2(new_n783), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n871), .B2(new_n872), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n884), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n865), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n902), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n675), .B1(new_n798), .B2(new_n800), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n748), .A2(new_n743), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n489), .B(KEYINPUT118), .Z(new_n911));
  NOR3_X1   g725(.A1(new_n742), .A2(new_n808), .A3(new_n675), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n705), .A2(new_n607), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n911), .C1(new_n913), .C2(new_n721), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT116), .B1(new_n912), .B2(new_n801), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n808), .A2(new_n675), .ZN(new_n916));
  AND4_X1   g730(.A1(KEYINPUT116), .A2(new_n916), .A3(new_n729), .A4(new_n801), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n732), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT48), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(KEYINPUT48), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n757), .A2(new_n607), .A3(new_n909), .A4(new_n759), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n808), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n845), .A2(new_n309), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n840), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT50), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n711), .A2(new_n300), .A3(new_n729), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n922), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n300), .A2(new_n729), .A3(new_n710), .A4(new_n707), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT50), .A3(new_n748), .A4(new_n909), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n763), .B1(new_n915), .B2(new_n917), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n630), .A2(new_n441), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n705), .A2(new_n912), .A3(new_n607), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT117), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT117), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n932), .A2(new_n933), .A3(new_n935), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(KEYINPUT51), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n921), .B1(new_n926), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT47), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n831), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n830), .A2(KEYINPUT47), .A3(new_n684), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n925), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n923), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n933), .A2(new_n935), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n932), .A2(KEYINPUT115), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n932), .A2(KEYINPUT115), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT51), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n901), .A2(new_n908), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT119), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n901), .A2(new_n908), .A3(new_n952), .A4(KEYINPUT119), .ZN(new_n956));
  OR2_X1    g770(.A1(G952), .A2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n848), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT120), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n848), .C1(new_n955), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n238), .A2(new_n274), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(new_n272), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT55), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n902), .A2(new_n906), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n307), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(G210), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT56), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n270), .A2(G952), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n968), .A2(new_n307), .A3(new_n296), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n966), .A2(new_n971), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n972), .A2(new_n977), .ZN(G51));
  NOR2_X1   g792(.A1(new_n968), .A2(new_n907), .ZN(new_n979));
  INV_X1    g793(.A(new_n908), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n775), .B(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n373), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n969), .A2(new_n821), .A3(new_n820), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n973), .B1(new_n984), .B2(new_n985), .ZN(G54));
  NAND3_X1  g800(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n425), .A3(new_n434), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .A4(new_n435), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n988), .A2(new_n974), .A3(new_n989), .ZN(G60));
  XNOR2_X1  g804(.A(new_n627), .B(KEYINPUT59), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n901), .B2(new_n908), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n624), .A2(new_n625), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n974), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n624), .B2(new_n625), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n979), .B2(new_n980), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT122), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT122), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT60), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n967), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n527), .A2(new_n535), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n973), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n967), .A2(new_n659), .A3(new_n1001), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT61), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT124), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT124), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1004), .A2(new_n1009), .A3(KEYINPUT61), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1004), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1006), .A2(KEYINPUT123), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1011), .A2(new_n1016), .ZN(G66));
  NOR2_X1   g831(.A1(new_n898), .A2(G953), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT125), .ZN(new_n1019));
  INV_X1    g833(.A(G224), .ZN(new_n1020));
  OAI21_X1  g834(.A(G953), .B1(new_n492), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n964), .B1(G898), .B2(new_n270), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1022), .B(new_n1023), .ZN(G69));
  AOI211_X1 g838(.A(new_n808), .B(new_n694), .C1(new_n721), .C2(new_n880), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n608), .B2(new_n598), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n835), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n858), .A2(new_n765), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n718), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT62), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1027), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n842), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n547), .A2(new_n550), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(KEYINPUT126), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n427), .A2(new_n429), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1036), .B(new_n1037), .Z(new_n1038));
  NOR2_X1   g852(.A1(new_n1038), .A2(G953), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n833), .A2(new_n768), .A3(new_n749), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n786), .A2(new_n793), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(KEYINPUT127), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1028), .B1(new_n810), .B2(new_n834), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1044), .A2(new_n1045), .A3(new_n270), .A4(new_n842), .ZN(new_n1046));
  NAND2_X1  g860(.A1(G900), .A2(G953), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g862(.A1(new_n1034), .A2(new_n1039), .B1(new_n1048), .B2(new_n1038), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n270), .B1(G227), .B2(G900), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1049), .B(new_n1050), .ZN(G72));
  NOR2_X1   g865(.A1(new_n587), .A2(new_n553), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1033), .A2(new_n842), .A3(new_n898), .ZN(new_n1053));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  AOI211_X1 g869(.A(new_n559), .B(new_n1052), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1044), .A2(new_n842), .A3(new_n1045), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1055), .B1(new_n1057), .B2(new_n884), .ZN(new_n1058));
  AND3_X1   g872(.A1(new_n1058), .A2(new_n559), .A3(new_n1052), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n564), .A2(new_n588), .ZN(new_n1060));
  AND4_X1   g874(.A1(new_n900), .A2(new_n887), .A3(new_n1055), .A4(new_n1060), .ZN(new_n1061));
  NOR4_X1   g875(.A1(new_n1056), .A2(new_n1059), .A3(new_n973), .A4(new_n1061), .ZN(G57));
endmodule


