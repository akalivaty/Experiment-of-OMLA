//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT74), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT75), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n205), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n207), .A2(new_n211), .A3(new_n215), .A4(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G155gat), .B(G162gat), .Z(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n209), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT76), .B(G148gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n216), .B1(new_n224), .B2(new_n205), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT3), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n220), .A2(new_n221), .B1(new_n225), .B2(new_n223), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G127gat), .B(G134gat), .Z(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n228), .A2(new_n231), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT77), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n234), .A2(new_n238), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n222), .A2(new_n244), .A3(new_n226), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n240), .A2(new_n243), .A3(new_n247), .A4(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n229), .B(new_n239), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT5), .B1(new_n251), .B2(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n245), .B(KEYINPUT4), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT5), .A3(new_n243), .A4(new_n240), .ZN(new_n255));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256));
  XNOR2_X1  g055(.A(G57gat), .B(G85gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n253), .A2(new_n255), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n255), .A3(new_n260), .ZN(new_n264));
  INV_X1    g063(.A(new_n261), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n253), .B2(new_n255), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n263), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(G211gat), .ZN(new_n271));
  OR2_X1    g070(.A1(KEYINPUT71), .A2(G218gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(G218gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n274), .B2(KEYINPUT22), .ZN(new_n275));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n270), .B(new_n276), .C1(new_n274), .C2(KEYINPUT22), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n290), .B2(G190gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT67), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND4_X1   g094(.A1(new_n288), .A2(new_n291), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n300), .B1(new_n298), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n309), .A2(new_n310), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  AND4_X1   g113(.A1(KEYINPUT25), .A2(new_n302), .A3(new_n305), .A4(new_n304), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n307), .A2(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n296), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n307), .A2(new_n308), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n314), .A2(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n288), .A2(new_n291), .A3(new_n292), .A4(new_n295), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n281), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n324), .A3(new_n317), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n296), .A2(new_n316), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n280), .B(new_n328), .C1(new_n329), .C2(new_n320), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n319), .A2(new_n325), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT72), .A3(new_n280), .ZN(new_n333));
  XNOR2_X1  g132(.A(G8gat), .B(G36gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT73), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n331), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n336), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n331), .B2(new_n333), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT30), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OR2_X1    g141(.A1(new_n341), .A2(KEYINPUT30), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT85), .B1(new_n269), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT35), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n264), .A2(new_n265), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n262), .B1(new_n347), .B2(new_n267), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n342), .A4(new_n343), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n345), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n278), .B2(new_n279), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n227), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n353));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n231), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n280), .B1(new_n358), .B2(KEYINPUT81), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT29), .B1(new_n229), .B2(new_n230), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n356), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n281), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n364), .B2(new_n353), .ZN(new_n365));
  OAI21_X1  g164(.A(G22gat), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n353), .A2(new_n355), .ZN(new_n367));
  INV_X1    g166(.A(new_n362), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n281), .B1(new_n360), .B2(new_n361), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G22gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n353), .B1(new_n360), .B2(new_n280), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n354), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(KEYINPUT82), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT80), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT31), .B(G50gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n370), .A2(new_n380), .A3(new_n371), .A4(new_n373), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n375), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n366), .A2(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n358), .A2(KEYINPUT81), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n384), .A2(new_n362), .A3(new_n281), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n385), .A2(new_n367), .B1(new_n354), .B2(new_n372), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n379), .B1(new_n386), .B2(new_n371), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(G22gat), .C1(new_n363), .C2(new_n365), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n239), .B1(new_n296), .B2(new_n316), .ZN(new_n392));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n323), .A2(new_n244), .A3(new_n324), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n392), .A2(new_n394), .A3(new_n393), .A4(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n393), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n296), .A2(new_n316), .A3(new_n239), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n244), .B1(new_n323), .B2(new_n324), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT32), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(G15gat), .B(G43gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n404), .B(KEYINPUT32), .C1(new_n406), .C2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n400), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n400), .A3(new_n413), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT70), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n411), .A2(new_n400), .A3(new_n417), .A4(new_n413), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n391), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n202), .B1(new_n351), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n350), .A2(new_n346), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n391), .A2(new_n419), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n422), .A2(KEYINPUT86), .A3(new_n423), .A4(new_n345), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n269), .A2(new_n344), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n418), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n414), .B(KEYINPUT69), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n425), .A2(new_n391), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n424), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n426), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT36), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT36), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n331), .A2(new_n333), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n340), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n436), .A2(new_n437), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT38), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n326), .B2(new_n330), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n442), .A2(KEYINPUT38), .A3(new_n337), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n341), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n269), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n254), .A2(new_n240), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n242), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n447), .A2(KEYINPUT39), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n251), .A2(new_n243), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n242), .B2(new_n446), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n260), .ZN(new_n453));
  NOR2_X1   g252(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n448), .A2(new_n452), .A3(new_n453), .A4(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n453), .B1(new_n447), .B2(KEYINPUT39), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n454), .B1(new_n457), .B2(new_n451), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n344), .A2(new_n264), .A3(new_n456), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n445), .A2(new_n459), .A3(new_n391), .ZN(new_n460));
  INV_X1    g259(.A(new_n391), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n269), .B2(new_n344), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n435), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n430), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n465));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT16), .ZN(new_n467));
  AOI21_X1  g266(.A(G1gat), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G8gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(KEYINPUT89), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n466), .B2(KEYINPUT89), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(new_n468), .A3(new_n471), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  OR2_X1    g276(.A1(G43gat), .A2(G50gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479));
  NAND2_X1  g278(.A1(G43gat), .A2(G50gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(G43gat), .A2(G50gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(G43gat), .A2(G50gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT15), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n487));
  INV_X1    g286(.A(G29gat), .ZN(new_n488));
  INV_X1    g287(.A(G36gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(KEYINPUT87), .A2(G29gat), .A3(G36gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n486), .A2(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n495), .A2(new_n497), .A3(new_n484), .ZN(new_n498));
  INV_X1    g297(.A(new_n486), .ZN(new_n499));
  NOR3_X1   g298(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n494), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT87), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  OAI22_X1  g301(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n484), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT88), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n496), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT17), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n497), .B1(new_n495), .B2(new_n484), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(KEYINPUT88), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n496), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n477), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n474), .A2(new_n476), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n508), .A2(new_n509), .B1(new_n495), .B2(new_n485), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n465), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n514), .B(KEYINPUT13), .Z(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n477), .A2(new_n506), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n516), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI221_X4 g323(.A(KEYINPUT17), .B1(new_n485), .B2(new_n495), .C1(new_n508), .C2(new_n509), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n511), .B1(new_n510), .B2(new_n496), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n515), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n477), .A2(new_n506), .B1(G229gat), .B2(G233gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n518), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G197gat), .ZN(new_n532));
  XOR2_X1   g331(.A(KEYINPUT11), .B(G169gat), .Z(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT12), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n518), .A2(new_n524), .A3(new_n529), .A4(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G71gat), .B(G78gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT90), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(KEYINPUT90), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G71gat), .ZN(new_n548));
  INV_X1    g347(.A(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n544), .A2(new_n543), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n545), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G127gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n552), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT91), .B1(new_n550), .B2(new_n551), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n555), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT92), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n555), .B1(KEYINPUT90), .B2(new_n540), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n568), .A2(new_n569), .B1(new_n541), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n477), .B1(new_n571), .B2(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n562), .B(G127gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n572), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n212), .ZN(new_n579));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n573), .A2(new_n576), .A3(new_n581), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G99gat), .B(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n592), .A2(new_n593), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n595), .A3(new_n589), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(KEYINPUT94), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n595), .B1(new_n598), .B2(new_n589), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n525), .B2(new_n526), .ZN(new_n606));
  NAND2_X1  g405(.A1(G232gat), .A2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT93), .Z(new_n608));
  INV_X1    g407(.A(KEYINPUT41), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n604), .B2(new_n506), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n606), .A2(new_n615), .A3(new_n611), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n608), .A2(new_n609), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G134gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G162gat), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n615), .B1(new_n606), .B2(new_n611), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(KEYINPUT95), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n594), .A2(new_n596), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n601), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n627), .B(new_n545), .C1(new_n556), .C2(new_n557), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n628), .B(new_n629), .C1(new_n571), .C2(new_n604), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n600), .B2(new_n603), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n571), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n605), .A2(new_n558), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n636), .B2(new_n628), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  INV_X1    g442(.A(new_n634), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n630), .B2(new_n632), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n645), .B2(new_n637), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n585), .A2(new_n625), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n464), .A2(new_n539), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT96), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n464), .A2(new_n651), .A3(new_n539), .A4(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n269), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT97), .B(G1gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n344), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n658), .A2(KEYINPUT98), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n470), .B1(new_n653), .B2(new_n344), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT98), .ZN(new_n663));
  INV_X1    g462(.A(new_n344), .ZN(new_n664));
  INV_X1    g463(.A(new_n657), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n664), .B(new_n665), .C1(new_n650), .C2(new_n652), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n666), .B2(KEYINPUT42), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n662), .B2(new_n667), .ZN(G1325gat));
  INV_X1    g467(.A(new_n653), .ZN(new_n669));
  INV_X1    g468(.A(new_n419), .ZN(new_n670));
  OR3_X1    g469(.A1(new_n669), .A2(G15gat), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G15gat), .B1(new_n669), .B2(new_n435), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1326gat));
  NAND2_X1  g472(.A1(new_n653), .A2(new_n461), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  INV_X1    g475(.A(new_n647), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n585), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n623), .A2(new_n624), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n464), .A2(new_n539), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n488), .A3(new_n269), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AND4_X1   g483(.A1(new_n460), .A2(new_n432), .A3(new_n462), .A4(new_n434), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n423), .A2(new_n346), .A3(new_n345), .A4(new_n350), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n202), .B1(KEYINPUT35), .B2(new_n428), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n424), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n688), .B2(new_n679), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n464), .A2(KEYINPUT44), .A3(new_n625), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n537), .A2(KEYINPUT99), .A3(new_n538), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT99), .B1(new_n537), .B2(new_n538), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697), .B2(new_n348), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n698), .ZN(G1328gat));
  OAI21_X1  g498(.A(G36gat), .B1(new_n697), .B2(new_n664), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n489), .A3(new_n344), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT100), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT46), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n681), .A2(new_n704), .A3(new_n489), .A4(new_n344), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(new_n435), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n689), .A2(new_n709), .A3(new_n690), .A4(new_n696), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G43gat), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n670), .A2(G43gat), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n464), .A2(new_n539), .A3(new_n680), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(KEYINPUT47), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n710), .A2(KEYINPUT102), .A3(G43gat), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT102), .B1(new_n710), .B2(G43gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n713), .B(KEYINPUT103), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT101), .B(KEYINPUT47), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(G1330gat));
  NAND4_X1  g519(.A1(new_n689), .A2(new_n461), .A3(new_n690), .A4(new_n696), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G50gat), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT48), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n681), .A2(new_n725), .A3(new_n461), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n722), .B(new_n726), .C1(new_n723), .C2(KEYINPUT48), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1331gat));
  NOR4_X1   g529(.A1(new_n585), .A2(new_n625), .A3(new_n677), .A4(new_n694), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n464), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n348), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT105), .B(G57gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n664), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  OAI21_X1  g539(.A(new_n548), .B1(new_n732), .B2(new_n670), .ZN(new_n741));
  INV_X1    g540(.A(new_n732), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n435), .A2(new_n548), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(KEYINPUT106), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT106), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n391), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n549), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n688), .A2(new_n679), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n585), .A2(new_n695), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT51), .B1(new_n750), .B2(new_n753), .ZN(new_n754));
  AND4_X1   g553(.A1(KEYINPUT51), .A2(new_n753), .A3(new_n464), .A4(new_n625), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n587), .A3(new_n269), .A4(new_n647), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n752), .A2(new_n677), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n691), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n348), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n689), .A2(new_n690), .A3(new_n758), .A4(new_n344), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G92gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(KEYINPUT108), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n664), .A2(G92gat), .A3(new_n677), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n754), .B2(new_n755), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n764), .C1(KEYINPUT108), .C2(new_n762), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n759), .B2(new_n435), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n670), .A2(G99gat), .A3(new_n677), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n391), .A2(G106gat), .A3(new_n677), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n754), .B2(new_n755), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n689), .A2(new_n690), .A3(new_n758), .A4(new_n461), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT109), .B(G106gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g581(.A1(new_n645), .A2(new_n637), .A3(new_n643), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n634), .B1(new_n571), .B2(new_n631), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n630), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n635), .B2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n789));
  AOI21_X1  g588(.A(new_n641), .B1(new_n645), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n783), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n633), .A2(new_n634), .A3(new_n789), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n630), .A2(new_n786), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT54), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n643), .C1(new_n794), .C2(new_n645), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n784), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n521), .A2(new_n522), .A3(new_n520), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n521), .A2(new_n800), .A3(new_n522), .A4(new_n520), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n514), .B1(new_n527), .B2(new_n521), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n801), .C1(new_n802), .C2(KEYINPUT111), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n804), .B(new_n514), .C1(new_n527), .C2(new_n521), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n534), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n797), .A2(new_n625), .A3(new_n538), .A4(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n806), .A2(new_n538), .A3(new_n647), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n694), .B2(new_n797), .ZN(new_n809));
  OAI211_X1 g608(.A(KEYINPUT113), .B(new_n807), .C1(new_n809), .C2(new_n625), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n527), .A2(new_n528), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n523), .B1(new_n813), .B2(new_n465), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n535), .B1(new_n814), .B2(new_n529), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n535), .A2(new_n518), .A3(new_n529), .A4(new_n524), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n537), .A2(KEYINPUT99), .A3(new_n538), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n791), .A4(new_n796), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n806), .A2(new_n538), .A3(new_n647), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n625), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n791), .A2(new_n796), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n538), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n679), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n811), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n825), .A3(new_n585), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n583), .A2(new_n584), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n827), .A2(new_n679), .A3(new_n677), .A4(new_n695), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n269), .A3(new_n664), .A4(new_n423), .ZN(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n539), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n348), .B1(new_n826), .B2(new_n828), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n427), .A2(new_n391), .A3(new_n426), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n344), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n694), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n833), .B1(new_n839), .B2(new_n831), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n830), .A2(new_n841), .A3(new_n677), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n647), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n841), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n830), .B2(new_n585), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n563), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n845), .B1(new_n837), .B2(new_n846), .ZN(G1342gat));
  OR3_X1    g646(.A1(new_n837), .A2(G134gat), .A3(new_n679), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(KEYINPUT56), .ZN(new_n850));
  OAI21_X1  g649(.A(G134gat), .B1(new_n830), .B2(new_n679), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT114), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n849), .A2(new_n850), .A3(new_n854), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(G1343gat));
  NOR3_X1   g655(.A1(new_n709), .A2(new_n391), .A3(new_n344), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(new_n834), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n858), .A2(new_n205), .A3(new_n539), .ZN(new_n859));
  XNOR2_X1  g658(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n709), .A2(new_n348), .A3(new_n344), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n391), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n795), .ZN(new_n866));
  XNOR2_X1  g665(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n791), .B(new_n539), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(KEYINPUT116), .A3(new_n820), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n679), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT116), .B1(new_n868), .B2(new_n820), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n807), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n820), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n679), .A3(new_n869), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n585), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n865), .B1(new_n879), .B2(new_n828), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n391), .B1(new_n826), .B2(new_n828), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n862), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n883), .B2(new_n832), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n883), .A2(new_n695), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n859), .B1(new_n886), .B2(G141gat), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(new_n224), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n858), .A2(new_n890), .A3(new_n647), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT119), .Z(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(KEYINPUT59), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n883), .B2(new_n677), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n896), .B(new_n893), .C1(new_n883), .C2(new_n677), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n807), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n585), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n648), .A2(new_n832), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n391), .B1(new_n903), .B2(KEYINPUT121), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n900), .A2(new_n585), .B1(new_n648), .B2(new_n832), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n829), .A2(new_n864), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n647), .B(new_n862), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n899), .B1(new_n911), .B2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n892), .B1(new_n898), .B2(new_n912), .ZN(G1345gat));
  NAND2_X1  g712(.A1(new_n827), .A2(G155gat), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT122), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n883), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(G155gat), .B1(new_n858), .B2(new_n827), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  NOR3_X1   g717(.A1(new_n883), .A2(new_n213), .A3(new_n679), .ZN(new_n919));
  AOI21_X1  g718(.A(G162gat), .B1(new_n858), .B2(new_n625), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n664), .A2(new_n269), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n829), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n835), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n694), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n829), .A2(new_n423), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT123), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n829), .A2(new_n928), .A3(new_n423), .A4(new_n922), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n539), .A2(G169gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(G1348gat));
  NAND3_X1  g731(.A1(new_n930), .A2(G176gat), .A3(new_n647), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  AOI21_X1  g735(.A(G176gat), .B1(new_n924), .B2(new_n647), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(G1349gat));
  INV_X1    g737(.A(G183gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n930), .B2(new_n827), .ZN(new_n940));
  NOR4_X1   g739(.A1(new_n923), .A2(new_n290), .A3(new_n835), .A4(new_n585), .ZN(new_n941));
  OR3_X1    g740(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT60), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT60), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n294), .A3(new_n625), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n927), .A2(new_n625), .A3(new_n929), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n294), .B1(new_n947), .B2(KEYINPUT61), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n946), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT126), .B(new_n945), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1351gat));
  AND2_X1   g755(.A1(new_n435), .A2(new_n922), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n881), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n694), .ZN(new_n959));
  INV_X1    g758(.A(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n461), .B1(new_n905), .B2(new_n906), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n901), .A2(new_n906), .A3(new_n902), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n863), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n960), .B1(new_n963), .B2(new_n909), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n539), .A2(G197gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n959), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n967), .A3(new_n647), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n968), .B(KEYINPUT62), .Z(new_n969));
  AOI211_X1 g768(.A(new_n677), .B(new_n960), .C1(new_n963), .C2(new_n909), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n647), .B1(new_n908), .B2(new_n910), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(KEYINPUT127), .A3(new_n960), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n271), .A3(new_n827), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n827), .B(new_n957), .C1(new_n908), .C2(new_n910), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n977), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n977), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  AOI21_X1  g779(.A(G218gat), .B1(new_n958), .B2(new_n625), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n679), .B1(new_n272), .B2(new_n273), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n964), .B2(new_n982), .ZN(G1355gat));
endmodule


