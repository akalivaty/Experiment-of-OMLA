//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n569, new_n570, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT67), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  INV_X1    g046(.A(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(G2104), .ZN(new_n473));
  OAI22_X1  g048(.A1(new_n470), .A2(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT66), .B1(new_n478), .B2(new_n468), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(new_n469), .A3(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n475), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(new_n483), .A3(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n474), .B1(new_n479), .B2(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n487), .B1(new_n470), .B2(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT68), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  AND4_X1   g070(.A1(G2105), .A2(new_n464), .A3(new_n467), .A4(new_n469), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G126), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n467), .A3(new_n469), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NOR3_X1   g076(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n477), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n500), .A2(KEYINPUT4), .B1(new_n477), .B2(new_n502), .ZN(new_n507));
  INV_X1    g082(.A(new_n493), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(G114), .B2(new_n468), .ZN(new_n509));
  INV_X1    g084(.A(G126), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n490), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT69), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(G164));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT70), .B(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n514), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n514), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n527), .A2(G50), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n533), .B1(new_n524), .B2(new_n526), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT72), .B(G88), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  NAND3_X1  g116(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n543), .A2(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n537), .A2(G89), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n527), .A2(G51), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  XOR2_X1   g127(.A(KEYINPUT74), .B(G90), .Z(new_n553));
  NAND2_X1  g128(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n527), .A2(G52), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n525), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  NAND2_X1  g134(.A1(new_n537), .A2(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n527), .A2(G43), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n525), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  AOI21_X1  g146(.A(new_n517), .B1(new_n525), .B2(KEYINPUT6), .ZN(new_n572));
  AND4_X1   g147(.A1(KEYINPUT71), .A2(new_n519), .A3(new_n521), .A4(KEYINPUT6), .ZN(new_n573));
  OAI21_X1  g148(.A(G543), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n527), .A2(new_n577), .A3(G53), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n530), .B2(new_n531), .ZN(new_n582));
  OAI21_X1  g157(.A(G65), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G91), .B2(new_n537), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n579), .A2(new_n586), .ZN(G299));
  OAI211_X1 g162(.A(G49), .B(G543), .C1(new_n572), .C2(new_n573), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n532), .B1(new_n572), .B2(new_n573), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(G288));
  NAND2_X1  g169(.A1(new_n537), .A2(G86), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n527), .A2(G48), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n530), .B2(new_n531), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT78), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n598), .B2(KEYINPUT78), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n522), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n595), .A2(new_n596), .A3(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n537), .A2(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n527), .A2(G47), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n605), .B(new_n606), .C1(new_n525), .C2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n537), .A2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(G66), .B1(new_n580), .B2(new_n582), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n516), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G54), .B2(new_n527), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n579), .A2(new_n586), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n564), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n618), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n480), .A2(new_n469), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(new_n473), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2100), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n639), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n490), .B2(new_n641), .ZN(new_n642));
  AND4_X1   g217(.A1(new_n468), .A2(new_n464), .A3(new_n467), .A4(new_n469), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n642), .B1(G135), .B2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n638), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XOR2_X1   g225(.A(G2427), .B(G2430), .Z(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT83), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n671), .B1(new_n668), .B2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT18), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2096), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G227));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n686), .B(new_n687), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n687), .ZN(new_n694));
  MUX2_X1   g269(.A(new_n693), .B(new_n694), .S(new_n685), .Z(new_n695));
  AOI21_X1  g270(.A(new_n682), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n692), .A2(new_n682), .A3(new_n695), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n697), .A2(G1986), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(G1986), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT87), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n702), .B1(new_n699), .B2(new_n700), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(new_n704), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(G229));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G32), .ZN(new_n711));
  INV_X1    g286(.A(G129), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n490), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  INV_X1    g293(.A(G141), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n718), .C1(new_n719), .C2(new_n470), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n711), .B1(new_n721), .B2(new_n710), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT27), .B(G1996), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(KEYINPUT24), .A2(G34), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n710), .B1(KEYINPUT24), .B2(G34), .ZN(new_n726));
  OAI22_X1  g301(.A1(G160), .A2(new_n710), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G5), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G171), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n724), .B1(G2084), .B2(new_n727), .C1(new_n731), .C2(G1961), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT97), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n565), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G19), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n710), .A2(G26), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n643), .A2(G140), .ZN(new_n740));
  INV_X1    g315(.A(G128), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n468), .A2(G116), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n490), .A2(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(new_n710), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n722), .A2(new_n723), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n735), .A2(new_n736), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n737), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n710), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(new_n468), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n754), .B(new_n756), .C1(G139), .C2(new_n643), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n752), .B1(new_n757), .B2(new_n710), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G2072), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G11), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n762), .A2(KEYINPUT95), .A3(G28), .ZN(new_n763));
  AOI21_X1  g338(.A(KEYINPUT95), .B1(new_n762), .B2(G28), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n710), .B1(new_n762), .B2(G28), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n644), .A2(G29), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT94), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n758), .A2(G2072), .B1(KEYINPUT94), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n727), .A2(G2084), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n767), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n728), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n728), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G1966), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n751), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n619), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT90), .B(G1348), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n779), .C1(G4), .C2(G16), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(G1961), .B2(new_n731), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n728), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT100), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT23), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G27), .A2(G29), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G164), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2078), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G162), .A2(G29), .ZN(new_n794));
  OR2_X1    g369(.A1(G29), .A2(G35), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n776), .A2(new_n783), .A3(new_n793), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n733), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G24), .B(G290), .S(G16), .Z(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(G1986), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n710), .A2(G25), .ZN(new_n807));
  OR2_X1    g382(.A1(G95), .A2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n808), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n809));
  INV_X1    g384(.A(G119), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n490), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G131), .B2(new_n643), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(new_n710), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G1991), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n728), .A2(G22), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G166), .B2(new_n728), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1971), .ZN(new_n821));
  MUX2_X1   g396(.A(G6), .B(G305), .S(G16), .Z(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT32), .B(G1981), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n592), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G16), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n728), .A2(G23), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT89), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT33), .B(G1976), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT89), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n828), .A2(new_n833), .A3(new_n829), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n825), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n832), .B1(new_n831), .B2(new_n834), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n818), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n837), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n839), .A2(KEYINPUT34), .A3(new_n835), .A4(new_n825), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n817), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT36), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI211_X1 g418(.A(KEYINPUT36), .B(new_n817), .C1(new_n838), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n804), .B1(new_n843), .B2(new_n844), .ZN(G150));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n846));
  XNOR2_X1  g421(.A(G150), .B(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n537), .A2(G93), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n527), .A2(G55), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n848), .B(new_n849), .C1(new_n525), .C2(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n564), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n851), .A2(new_n564), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n619), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g437(.A(G860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n854), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(G162), .B(new_n644), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(G160), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n721), .B(new_n757), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n812), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n812), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n501), .A2(KEYINPUT104), .A3(new_n503), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT104), .B1(new_n501), .B2(new_n503), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n497), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n745), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n643), .A2(G142), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n496), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n468), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n635), .B(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n872), .A2(new_n878), .A3(new_n873), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n880), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n870), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(new_n870), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n892), .A2(KEYINPUT105), .A3(new_n893), .A4(new_n888), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n858), .A2(new_n630), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n855), .B(new_n857), .C1(G559), .C2(new_n618), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n618), .A2(new_n623), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n619), .A2(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n618), .A2(KEYINPUT107), .A3(new_n623), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n619), .B2(G299), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n906), .A2(new_n907), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT108), .B1(new_n900), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n901), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n898), .A2(new_n899), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n904), .A2(KEYINPUT106), .A3(new_n901), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n904), .B2(new_n901), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n900), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n910), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n827), .B(G290), .Z(new_n925));
  XNOR2_X1  g500(.A(G303), .B(G305), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n925), .B(new_n926), .Z(new_n927));
  AOI21_X1  g502(.A(new_n927), .B1(new_n922), .B2(KEYINPUT42), .ZN(new_n928));
  INV_X1    g503(.A(new_n923), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n910), .A2(new_n916), .A3(new_n929), .A4(new_n920), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n924), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n924), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n854), .A2(new_n628), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n934), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(G168), .A2(KEYINPUT110), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  NAND2_X1  g515(.A1(G286), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(G301), .A3(new_n941), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n855), .A3(new_n857), .A4(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n944), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n565), .B1(new_n852), .B2(new_n853), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n946), .A2(new_n942), .B1(new_n947), .B2(new_n856), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n913), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n904), .A2(new_n901), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n927), .A3(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n953), .A2(new_n895), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n952), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n925), .B(new_n926), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n938), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n908), .A2(new_n903), .A3(new_n905), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n907), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n945), .B(new_n948), .C1(new_n917), .C2(new_n918), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n956), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n953), .A2(new_n895), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n937), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n957), .A2(new_n938), .A3(new_n895), .A4(new_n953), .ZN(new_n968));
  AND4_X1   g543(.A1(KEYINPUT111), .A2(new_n967), .A3(new_n968), .A4(KEYINPUT44), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n937), .B1(new_n964), .B2(KEYINPUT43), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT111), .B1(new_n970), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(G397));
  NOR2_X1   g547(.A1(new_n473), .A2(new_n472), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n643), .B2(G137), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n483), .B1(new_n482), .B2(G2105), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT66), .B(new_n468), .C1(new_n481), .C2(new_n475), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n974), .B(G40), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(G160), .A2(KEYINPUT113), .A3(G40), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT112), .B(G1384), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n877), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(KEYINPUT114), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n745), .A2(new_n747), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n740), .A2(G2067), .A3(new_n744), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n721), .B2(new_n986), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n991), .A2(new_n721), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n812), .B(new_n814), .Z(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(G290), .B(G1986), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n999), .B1(new_n985), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n504), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n507), .A2(KEYINPUT104), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n511), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT50), .B1(new_n1006), .B2(G1384), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n506), .A2(new_n512), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n981), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n788), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT119), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1014), .A3(new_n788), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n506), .A2(new_n512), .A3(new_n1009), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n877), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT56), .B(G2072), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n981), .A2(new_n1019), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n623), .A2(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1002), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT120), .B(new_n1028), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n877), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n981), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT122), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n981), .A2(new_n1032), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n779), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1006), .A2(G1384), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n981), .A2(new_n1039), .A3(new_n747), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1031), .B(new_n619), .C1(new_n1038), .C2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n619), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1025), .A2(new_n1023), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1011), .A2(new_n1014), .A3(new_n788), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1014), .B1(new_n1011), .B2(new_n788), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1022), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1044), .A2(KEYINPUT123), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1030), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n981), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT124), .B(G1996), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT58), .B(G1341), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n981), .B2(new_n1039), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n565), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT59), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n565), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1045), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1026), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT61), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1048), .A2(new_n1045), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1035), .A2(new_n779), .A3(new_n1037), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(new_n619), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(KEYINPUT60), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1050), .B1(new_n1069), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1961), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1035), .A2(new_n1078), .A3(new_n1037), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1035), .A2(KEYINPUT125), .A3(new_n1078), .A4(new_n1037), .ZN(new_n1082));
  INV_X1    g657(.A(G2078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(new_n474), .C1(G2105), .C2(new_n482), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1020), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT126), .B1(new_n1086), .B2(new_n984), .ZN(new_n1087));
  INV_X1    g662(.A(new_n984), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1020), .A4(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n981), .A2(new_n1019), .A3(new_n1020), .A4(new_n1083), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1087), .A2(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1081), .A2(new_n1082), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT127), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT127), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1097), .A3(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1092), .A2(new_n1091), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1083), .A2(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1018), .B1(new_n1006), .B2(G1384), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1018), .A2(G1384), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n506), .A2(new_n512), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n981), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1079), .B(new_n1099), .C1(new_n1100), .C2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1096), .A2(KEYINPUT54), .A3(new_n1098), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1109));
  AND3_X1   g684(.A1(G303), .A2(G8), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(G303), .B2(G8), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1971), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1051), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1007), .A2(new_n981), .A3(new_n799), .A4(new_n1010), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G8), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1108), .B(new_n1112), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  OR2_X1    g693(.A1(G305), .A2(G1981), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G305), .A2(G1981), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT49), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1117), .B1(new_n981), .B2(new_n1039), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(KEYINPUT49), .A3(new_n1120), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n592), .A2(new_n826), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n592), .A2(new_n826), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(G1976), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT52), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1126), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1117), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1112), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT116), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1114), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1034), .A2(G2090), .ZN(new_n1140));
  OAI211_X1 g715(.A(G8), .B(new_n1137), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1118), .A2(new_n1135), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1034), .A2(G2084), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g719(.A(G1966), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1104), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n977), .A2(new_n978), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT113), .B1(G160), .B2(G40), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1103), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT45), .B1(new_n877), .B2(new_n1009), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(KEYINPUT117), .ZN(new_n1153));
  AOI21_X1  g728(.A(G168), .B1(new_n1147), .B2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1153), .A2(G168), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(G8), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT51), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT51), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1155), .A2(new_n1158), .A3(G8), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1142), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1105), .A2(G171), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1094), .B2(G171), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1107), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1077), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1153), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G286), .A2(new_n1117), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1168), .B1(new_n1142), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1169), .A2(KEYINPUT63), .A3(new_n1170), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(G8), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1112), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1173), .A2(new_n1175), .A3(KEYINPUT118), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1177), .A2(KEYINPUT63), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1172), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1141), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1185));
  INV_X1    g760(.A(G288), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1185), .A2(new_n1132), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1119), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1184), .A2(new_n1135), .B1(new_n1188), .B2(new_n1124), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1142), .A2(new_n1162), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1169), .A2(G286), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1191), .A2(G8), .A3(new_n1155), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1159), .B1(new_n1192), .B2(KEYINPUT51), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1190), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1157), .A2(new_n1160), .A3(new_n1194), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1183), .B(new_n1189), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1001), .B1(new_n1167), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT46), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n991), .B(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n994), .A2(new_n721), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n985), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT47), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n814), .B(new_n811), .C1(G131), .C2(new_n643), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n996), .A2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n985), .B1(new_n1206), .B2(new_n993), .ZN(new_n1207));
  NOR2_X1   g782(.A1(G290), .A2(G1986), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n985), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT48), .Z(new_n1210));
  OAI211_X1 g785(.A(new_n1204), .B(new_n1207), .C1(new_n999), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1198), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g788(.A1(new_n958), .A2(new_n965), .ZN(new_n1215));
  NOR3_X1   g789(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1216));
  OAI211_X1 g790(.A(new_n896), .B(new_n1216), .C1(new_n707), .C2(new_n708), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1215), .A2(new_n1217), .ZN(G308));
  OR2_X1    g792(.A1(new_n1215), .A2(new_n1217), .ZN(G225));
endmodule


