//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  OR3_X1    g005(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT28), .ZN(new_n211));
  NAND2_X1  g010(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT68), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(new_n212), .ZN(new_n220));
  AOI211_X1 g019(.A(new_n211), .B(G190gat), .C1(new_n215), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n212), .ZN(new_n222));
  INV_X1    g021(.A(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n206), .B(new_n210), .C1(new_n221), .C2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(new_n220), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n219), .B1(new_n218), .B2(new_n212), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(new_n211), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n206), .A4(new_n210), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n240));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  INV_X1    g045(.A(G176gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT23), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT23), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n248), .A2(new_n250), .A3(new_n208), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n245), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n248), .A2(new_n250), .A3(new_n208), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(new_n242), .B2(KEYINPUT64), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n242), .A2(new_n255), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(KEYINPUT25), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT66), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264));
  AOI211_X1 g063(.A(new_n264), .B(new_n261), .C1(new_n253), .C2(new_n258), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n237), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT1), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  OR3_X1    g070(.A1(new_n271), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT71), .B1(new_n271), .B2(G113gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274));
  INV_X1    g073(.A(G113gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(G120gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n272), .A2(new_n273), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G227gat), .ZN(new_n284));
  INV_X1    g083(.A(G233gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n237), .B(new_n281), .C1(new_n263), .C2(new_n265), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  XNOR2_X1  g088(.A(G15gat), .B(G43gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G71gat), .ZN(new_n291));
  INV_X1    g090(.A(G99gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n288), .B2(new_n294), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n289), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n283), .A2(new_n287), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT34), .B1(new_n298), .B2(new_n286), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n286), .B1(new_n283), .B2(new_n287), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT34), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n293), .A2(KEYINPUT33), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n288), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n297), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n303), .B1(new_n297), .B2(new_n305), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n204), .B(new_n205), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n297), .A2(new_n305), .ZN(new_n309));
  INV_X1    g108(.A(new_n303), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n297), .A2(new_n303), .A3(new_n305), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n311), .A2(new_n202), .A3(new_n203), .A4(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n318));
  OR2_X1    g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G197gat), .A2(G204gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n317), .B(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n257), .B1(new_n254), .B2(new_n256), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n262), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n228), .ZN(new_n326));
  NAND2_X1  g125(.A1(G226gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n264), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n262), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT29), .B1(new_n332), .B2(new_n237), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n327), .B(KEYINPUT75), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n322), .B(new_n329), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n322), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n332), .B2(new_n237), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n328), .B1(new_n326), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G8gat), .B(G36gat), .ZN(new_n343));
  INV_X1    g142(.A(G64gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(G92gat), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n342), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n346), .B(KEYINPUT76), .Z(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT77), .B1(new_n342), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n336), .A2(new_n341), .A3(new_n356), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n352), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G57gat), .ZN(new_n362));
  INV_X1    g161(.A(G85gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G162gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G162gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n368), .A3(G155gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G155gat), .B(G162gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(KEYINPUT2), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n377), .A2(new_n373), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(KEYINPUT79), .A3(new_n372), .A4(new_n373), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n281), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n376), .A2(new_n386), .A3(new_n378), .A4(new_n379), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n281), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n383), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n392), .B1(new_n396), .B2(new_n382), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n281), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n391), .B1(new_n382), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT81), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n381), .B1(new_n388), .B2(new_n383), .ZN(new_n404));
  INV_X1    g203(.A(new_n398), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n404), .A2(new_n392), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  NOR4_X1   g206(.A1(new_n406), .A2(new_n407), .A3(new_n395), .A4(new_n401), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n364), .B(new_n394), .C1(new_n403), .C2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n382), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n391), .A3(new_n398), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(KEYINPUT5), .A3(new_n402), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n407), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT81), .A3(new_n402), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n364), .B1(new_n417), .B2(new_n394), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n394), .B1(new_n403), .B2(new_n408), .ZN(new_n420));
  INV_X1    g219(.A(new_n364), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n359), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT31), .B(G50gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n386), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n380), .ZN(new_n429));
  AND2_X1   g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n429), .A2(G78gat), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(G78gat), .B1(new_n429), .B2(new_n430), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n380), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n387), .A2(new_n339), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n322), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G22gat), .ZN(new_n439));
  INV_X1    g238(.A(G106gat), .ZN(new_n440));
  INV_X1    g239(.A(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n441), .A3(new_n437), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G106gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n431), .A2(new_n426), .A3(new_n432), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n434), .A2(new_n443), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n443), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n431), .A2(new_n426), .A3(new_n432), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n433), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n424), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n314), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n420), .A2(new_n421), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n410), .A3(new_n409), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n422), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(new_n359), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n308), .A2(new_n313), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT83), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n352), .A2(new_n358), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n384), .A2(new_n389), .A3(new_n392), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n382), .A2(new_n391), .A3(new_n400), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(KEYINPUT84), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n463), .B(new_n466), .C1(KEYINPUT84), .C2(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(new_n364), .C1(KEYINPUT39), .C2(new_n463), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT40), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n456), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n336), .A2(KEYINPUT37), .A3(new_n341), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT86), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n346), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n342), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n471), .B2(new_n346), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n478), .A3(new_n422), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n329), .B1(new_n333), .B2(new_n335), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n474), .B1(new_n480), .B2(new_n337), .ZN(new_n481));
  OR3_X1    g280(.A1(new_n338), .A2(new_n340), .A3(new_n337), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n354), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT38), .B1(new_n342), .B2(new_n474), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(KEYINPUT85), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT85), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n348), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n455), .B(new_n470), .C1(new_n479), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n454), .A2(new_n461), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n462), .B1(new_n457), .B2(new_n422), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n306), .A2(new_n307), .A3(new_n451), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(KEYINPUT87), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n490), .B2(new_n491), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n499));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(G29gat), .ZN(new_n505));
  INV_X1    g304(.A(G36gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT89), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT91), .B(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G29gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OR3_X1    g313(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT90), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n503), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n507), .A2(new_n508), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(KEYINPUT92), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n501), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n503), .A3(new_n513), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n499), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  XOR2_X1   g322(.A(G15gat), .B(G22gat), .Z(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n526), .B2(KEYINPUT93), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(G1gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n527), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n511), .A3(new_n513), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n502), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT17), .A3(new_n520), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n531), .B1(new_n516), .B2(new_n521), .ZN(new_n537));
  NAND2_X1  g336(.A1(G229gat), .A2(G233gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(new_n534), .A3(new_n520), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n537), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n538), .B(KEYINPUT94), .Z(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT13), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n538), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n541), .A2(new_n547), .A3(new_n555), .A4(new_n548), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT97), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(KEYINPUT97), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(G71gat), .A2(G78gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n563), .B(new_n564), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT98), .B(G57gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(G64gat), .ZN(new_n571));
  INV_X1    g370(.A(G57gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(G64gat), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT99), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT99), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n569), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n344), .A2(G57gat), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n563), .B(new_n564), .C1(new_n573), .C2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n567), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n568), .B(KEYINPUT96), .Z(new_n583));
  AND3_X1   g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(KEYINPUT100), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n562), .B(KEYINPUT97), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n567), .A2(new_n568), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n577), .B1(new_n571), .B2(new_n574), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT99), .B(new_n573), .C1(new_n570), .C2(G64gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT19), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n585), .A2(KEYINPUT21), .A3(new_n594), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n604), .A2(new_n605), .A3(new_n532), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n604), .B2(new_n532), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n532), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT101), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n605), .A3(new_n532), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(KEYINPUT19), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT20), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n608), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n608), .B2(new_n612), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n602), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n614), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n608), .A2(new_n612), .A3(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n601), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OR2_X1    g424(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n626), .A2(G85gat), .A3(G92gat), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n629));
  NAND2_X1  g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(KEYINPUT8), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n628), .B(new_n632), .C1(G85gat), .C2(G92gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n522), .A2(new_n535), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n516), .B2(new_n521), .ZN(new_n638));
  NAND3_X1  g437(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(G134gat), .ZN(new_n641));
  INV_X1    g440(.A(G134gat), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n637), .A2(new_n642), .A3(new_n638), .A4(new_n639), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n625), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G162gat), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n641), .A2(new_n643), .A3(new_n625), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n647), .ZN(new_n650));
  INV_X1    g449(.A(new_n648), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n644), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n635), .B1(new_n585), .B2(new_n594), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n635), .A2(new_n591), .A3(new_n593), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n654), .A2(new_n656), .A3(KEYINPUT10), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n594), .A4(new_n635), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n653), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n653), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n654), .B2(new_n656), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n247), .ZN(new_n664));
  INV_X1    g463(.A(G204gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n660), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n660), .B2(new_n662), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n623), .A2(new_n649), .A3(new_n652), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n649), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n623), .A4(new_n671), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n498), .A2(new_n561), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n458), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n525), .ZN(G1324gat));
  AND3_X1   g480(.A1(new_n498), .A2(new_n561), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n462), .ZN(new_n683));
  NOR2_X1   g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n528), .A2(new_n523), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n523), .B1(new_n682), .B2(new_n462), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(G15gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n679), .A2(new_n691), .A3(new_n314), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n306), .A2(new_n307), .ZN(new_n693));
  AOI21_X1  g492(.A(G15gat), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(KEYINPUT104), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n455), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  AOI21_X1  g499(.A(new_n675), .B1(new_n489), .B2(new_n497), .ZN(new_n701));
  INV_X1    g500(.A(new_n561), .ZN(new_n702));
  INV_X1    g501(.A(new_n671), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n623), .A3(new_n703), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n458), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n505), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n498), .B2(new_n674), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n488), .A2(new_n314), .A3(new_n452), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n675), .B1(new_n497), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n715), .A2(new_n706), .A3(new_n704), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n708), .B1(new_n505), .B2(new_n716), .ZN(G1328gat));
  OAI211_X1 g516(.A(new_n462), .B(new_n704), .C1(new_n710), .C2(new_n714), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n718), .A2(new_n512), .ZN(new_n719));
  INV_X1    g518(.A(new_n512), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n701), .A2(new_n720), .A3(new_n462), .A4(new_n704), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT107), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n512), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n722), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n721), .A2(new_n722), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n724), .A2(new_n729), .ZN(G1329gat));
  NAND2_X1  g529(.A1(new_n705), .A2(new_n693), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n314), .A2(new_n732), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n704), .B(new_n734), .C1(new_n710), .C2(new_n714), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT47), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  OAI211_X1 g537(.A(new_n451), .B(new_n704), .C1(new_n710), .C2(new_n714), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  INV_X1    g540(.A(G50gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n705), .A2(new_n742), .A3(new_n451), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n741), .B1(new_n740), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1331gat));
  AOI21_X1  g545(.A(new_n561), .B1(new_n497), .B2(new_n711), .ZN(new_n747));
  INV_X1    g546(.A(new_n623), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n674), .A3(new_n671), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n458), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n570), .ZN(G1332gat));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n462), .A3(new_n749), .ZN(new_n753));
  AND2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT108), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1333gat));
  OAI21_X1  g557(.A(G71gat), .B1(new_n750), .B2(new_n314), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n693), .A2(new_n565), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g561(.A1(new_n750), .A2(new_n455), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT109), .B(G78gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n561), .A2(new_n623), .ZN(new_n767));
  AND3_X1   g566(.A1(new_n712), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n712), .B2(new_n767), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n768), .A2(new_n769), .A3(new_n671), .ZN(new_n770));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n706), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n561), .A2(new_n623), .A3(new_n671), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n715), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n458), .A2(new_n363), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(G1336gat));
  OAI211_X1 g574(.A(new_n462), .B(new_n772), .C1(new_n710), .C2(new_n714), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n359), .A2(G92gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT52), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1337gat));
  OAI211_X1 g583(.A(new_n460), .B(new_n772), .C1(new_n710), .C2(new_n714), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(G99gat), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n770), .A2(new_n292), .A3(new_n693), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1338gat));
  OAI211_X1 g590(.A(new_n451), .B(new_n772), .C1(new_n710), .C2(new_n714), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n768), .A2(new_n769), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n794), .A2(new_n440), .A3(new_n703), .A4(new_n451), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT53), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1339gat));
  AND3_X1   g599(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n592), .B1(new_n591), .B2(new_n593), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n636), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT10), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n655), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT54), .B(new_n661), .C1(new_n805), .C2(new_n658), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT112), .B1(new_n806), .B2(new_n667), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n661), .A3(new_n658), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT111), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n805), .A2(new_n810), .A3(new_n661), .A4(new_n658), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n809), .A2(new_n660), .A3(KEYINPUT54), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n653), .C1(new_n657), .C2(new_n659), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n666), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n807), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n561), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n807), .A2(new_n812), .A3(KEYINPUT55), .A4(new_n816), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT113), .B1(new_n821), .B2(new_n668), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(KEYINPUT113), .A3(new_n668), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n542), .A2(new_n537), .A3(new_n545), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n542), .A2(new_n537), .A3(new_n828), .A4(new_n545), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n538), .B1(new_n536), .B2(new_n537), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n554), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT115), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n558), .B(KEYINPUT95), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n703), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n674), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n823), .A2(new_n674), .A3(new_n824), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n833), .A2(new_n834), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n819), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n748), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n672), .A2(new_n561), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(new_n491), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n458), .A2(new_n462), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n702), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(new_n275), .ZN(G1340gat));
  INV_X1    g649(.A(new_n848), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n703), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n271), .A2(KEYINPUT116), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n271), .A2(KEYINPUT116), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n852), .B2(new_n853), .ZN(G1341gat));
  NOR2_X1   g655(.A1(new_n848), .A2(new_n748), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(G127gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n857), .B2(G127gat), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n857), .A2(G127gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1342gat));
  NAND2_X1  g661(.A1(new_n851), .A2(new_n674), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT56), .B1(new_n863), .B2(G134gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(G134gat), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n863), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n868), .B(KEYINPUT56), .C1(new_n863), .C2(G134gat), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n865), .A2(new_n866), .A3(new_n867), .A4(new_n869), .ZN(G1343gat));
  NOR3_X1   g669(.A1(new_n460), .A2(new_n458), .A3(new_n462), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n817), .A2(KEYINPUT119), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n807), .A2(new_n812), .A3(new_n873), .A4(new_n816), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n818), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n821), .A2(new_n668), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n561), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n674), .B1(new_n836), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n748), .B1(new_n879), .B2(new_n841), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n455), .B1(new_n880), .B2(new_n844), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n871), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n821), .A2(new_n668), .A3(KEYINPUT113), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n822), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n674), .A3(new_n839), .A4(new_n819), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n835), .B1(new_n885), .B2(new_n820), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n674), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n843), .B1(new_n888), .B2(new_n748), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n455), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n883), .A2(new_n890), .A3(new_n702), .ZN(new_n891));
  INV_X1    g690(.A(G141gat), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT120), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n845), .A2(new_n451), .A3(new_n871), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n892), .A3(new_n561), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n891), .B2(new_n892), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n893), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1344gat));
  INV_X1    g699(.A(G148gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n901), .A3(new_n703), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT57), .B1(new_n889), .B2(new_n455), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n836), .A2(new_n878), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n675), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n623), .B1(new_n906), .B2(new_n886), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n673), .A2(new_n677), .A3(new_n702), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n673), .A2(new_n677), .A3(new_n910), .A4(new_n702), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n882), .B(new_n451), .C1(new_n907), .C2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n904), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n703), .A3(new_n871), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n903), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n883), .A2(new_n890), .ZN(new_n917));
  AOI211_X1 g716(.A(KEYINPUT59), .B(new_n901), .C1(new_n917), .C2(new_n703), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n902), .B1(new_n916), .B2(new_n918), .ZN(G1345gat));
  AOI21_X1  g718(.A(G155gat), .B1(new_n894), .B2(new_n623), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n623), .A2(G155gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n917), .B2(new_n921), .ZN(G1346gat));
  NAND2_X1  g721(.A1(new_n366), .A2(new_n368), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n894), .A2(new_n923), .A3(new_n674), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n883), .A2(new_n890), .A3(new_n675), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n923), .B2(new_n926), .ZN(G1347gat));
  NAND3_X1  g726(.A1(new_n458), .A2(new_n693), .A3(new_n462), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT124), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n845), .A2(new_n455), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n702), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n889), .A2(new_n932), .A3(new_n706), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n845), .B2(new_n458), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n462), .B(new_n491), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n561), .A2(new_n246), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(G1348gat));
  NOR3_X1   g736(.A1(new_n930), .A2(new_n247), .A3(new_n671), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n247), .B1(new_n935), .B2(new_n671), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n930), .B2(new_n748), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n623), .B1(new_n233), .B2(new_n232), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n930), .B2(new_n675), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n674), .A2(new_n223), .ZN(new_n951));
  OAI22_X1  g750(.A1(new_n949), .A2(new_n950), .B1(new_n935), .B2(new_n951), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n460), .A2(new_n706), .A3(new_n359), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n914), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n561), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G197gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n359), .A2(new_n455), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n314), .B(new_n957), .C1(new_n934), .C2(new_n933), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n702), .A2(G197gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  NAND3_X1  g759(.A1(new_n845), .A2(KEYINPUT123), .A3(new_n458), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n932), .B1(new_n889), .B2(new_n706), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n460), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n963), .A2(new_n665), .A3(new_n703), .A4(new_n957), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n914), .A2(new_n703), .A3(new_n953), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n965), .A2(new_n966), .B1(G204gat), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n964), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT126), .B1(new_n964), .B2(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G1353gat));
  OR3_X1    g770(.A1(new_n958), .A2(G211gat), .A3(new_n748), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n904), .A2(new_n623), .A3(new_n913), .A4(new_n953), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n914), .A2(new_n974), .A3(new_n623), .A4(new_n953), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n978));
  AND4_X1   g777(.A1(KEYINPUT63), .A2(new_n977), .A3(G211gat), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n972), .B1(new_n976), .B2(new_n979), .ZN(G1354gat));
  INV_X1    g779(.A(G218gat), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n675), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n674), .A3(new_n957), .ZN(new_n983));
  AOI22_X1  g782(.A1(new_n954), .A2(new_n982), .B1(new_n983), .B2(new_n981), .ZN(G1355gat));
endmodule


