

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747;

  AND2_X1 U376 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U377 ( .A1(n555), .A2(n556), .ZN(n377) );
  INV_X2 U378 ( .A(G953), .ZN(n734) );
  XNOR2_X1 U379 ( .A(n528), .B(KEYINPUT35), .ZN(n745) );
  AND2_X4 U380 ( .A1(n610), .A2(n681), .ZN(n710) );
  NOR2_X2 U381 ( .A1(n662), .A2(n659), .ZN(n373) );
  XNOR2_X2 U382 ( .A(n433), .B(n512), .ZN(n687) );
  XNOR2_X2 U383 ( .A(n487), .B(n466), .ZN(n512) );
  XNOR2_X2 U384 ( .A(n583), .B(KEYINPUT1), .ZN(n641) );
  XNOR2_X2 U385 ( .A(n513), .B(G469), .ZN(n583) );
  NAND2_X1 U386 ( .A1(n656), .A2(n655), .ZN(n662) );
  NOR2_X1 U387 ( .A1(n589), .A2(n588), .ZN(n591) );
  XNOR2_X1 U388 ( .A(n373), .B(n558), .ZN(n674) );
  NAND2_X1 U389 ( .A1(n562), .A2(n638), .ZN(n642) );
  XNOR2_X1 U390 ( .A(n404), .B(n401), .ZN(n711) );
  XNOR2_X1 U391 ( .A(n504), .B(n405), .ZN(n404) );
  XNOR2_X1 U392 ( .A(n462), .B(KEYINPUT4), .ZN(n730) );
  XNOR2_X1 U393 ( .A(n471), .B(n403), .ZN(n498) );
  XOR2_X1 U394 ( .A(G146), .B(G125), .Z(n471) );
  XNOR2_X2 U395 ( .A(n584), .B(n547), .ZN(n656) );
  NAND2_X1 U396 ( .A1(n494), .A2(n393), .ZN(n392) );
  INV_X1 U397 ( .A(G902), .ZN(n393) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U399 ( .A(G131), .B(G134), .ZN(n727) );
  NOR2_X1 U400 ( .A1(n631), .A2(n421), .ZN(n586) );
  NAND2_X1 U401 ( .A1(n422), .A2(n585), .ZN(n421) );
  XNOR2_X1 U402 ( .A(n623), .B(n398), .ZN(n422) );
  XNOR2_X1 U403 ( .A(n566), .B(n374), .ZN(n589) );
  INV_X1 U404 ( .A(KEYINPUT46), .ZN(n374) );
  NOR2_X1 U405 ( .A1(n744), .A2(n742), .ZN(n566) );
  INV_X1 U406 ( .A(n394), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n730), .B(n463), .ZN(n487) );
  XNOR2_X1 U408 ( .A(KEYINPUT65), .B(G101), .ZN(n463) );
  XNOR2_X1 U409 ( .A(n468), .B(n467), .ZN(n488) );
  XNOR2_X1 U410 ( .A(n427), .B(KEYINPUT3), .ZN(n468) );
  XNOR2_X1 U411 ( .A(G113), .B(KEYINPUT69), .ZN(n427) );
  INV_X1 U412 ( .A(n729), .ZN(n401) );
  XNOR2_X1 U413 ( .A(n501), .B(n406), .ZN(n405) );
  XNOR2_X1 U414 ( .A(n727), .B(G146), .ZN(n507) );
  XNOR2_X1 U415 ( .A(n372), .B(n523), .ZN(n676) );
  NOR2_X1 U416 ( .A1(n534), .A2(n540), .ZN(n372) );
  XNOR2_X1 U417 ( .A(n377), .B(n557), .ZN(n596) );
  INV_X1 U418 ( .A(KEYINPUT39), .ZN(n557) );
  INV_X1 U419 ( .A(n745), .ZN(n369) );
  INV_X1 U420 ( .A(n437), .ZN(n390) );
  INV_X1 U421 ( .A(G472), .ZN(n492) );
  XNOR2_X1 U422 ( .A(KEYINPUT5), .B(KEYINPUT96), .ZN(n380) );
  INV_X1 U423 ( .A(KEYINPUT10), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n365), .B(n471), .ZN(n435) );
  XNOR2_X1 U425 ( .A(n470), .B(n436), .ZN(n365) );
  INV_X1 U426 ( .A(KEYINPUT76), .ZN(n436) );
  XOR2_X1 U427 ( .A(KEYINPUT75), .B(KEYINPUT89), .Z(n470) );
  XNOR2_X1 U428 ( .A(n648), .B(n425), .ZN(n540) );
  XNOR2_X1 U429 ( .A(n426), .B(KEYINPUT99), .ZN(n425) );
  INV_X1 U430 ( .A(KEYINPUT6), .ZN(n426) );
  XNOR2_X1 U431 ( .A(KEYINPUT16), .B(G122), .ZN(n469) );
  XNOR2_X1 U432 ( .A(n452), .B(n409), .ZN(n503) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n452) );
  XNOR2_X1 U434 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U435 ( .A(KEYINPUT67), .ZN(n410) );
  XOR2_X1 U436 ( .A(G134), .B(G122), .Z(n454) );
  XNOR2_X1 U437 ( .A(G107), .B(G116), .ZN(n453) );
  XNOR2_X1 U438 ( .A(n462), .B(n457), .ZN(n413) );
  XOR2_X1 U439 ( .A(G122), .B(G113), .Z(n441) );
  XNOR2_X1 U440 ( .A(G140), .B(G104), .ZN(n440) );
  XOR2_X1 U441 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n445) );
  XNOR2_X1 U442 ( .A(G143), .B(G131), .ZN(n447) );
  XOR2_X1 U443 ( .A(G137), .B(G140), .Z(n510) );
  XNOR2_X1 U444 ( .A(KEYINPUT68), .B(KEYINPUT48), .ZN(n590) );
  NOR2_X1 U445 ( .A1(n524), .A2(n676), .ZN(n526) );
  NOR2_X1 U446 ( .A1(n560), .A2(n659), .ZN(n460) );
  NOR2_X1 U447 ( .A1(n554), .A2(n559), .ZN(n582) );
  NAND2_X1 U448 ( .A1(n381), .A2(n355), .ZN(n554) );
  NAND2_X1 U449 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n506), .B(n505), .ZN(n562) );
  NOR2_X1 U451 ( .A1(n708), .A2(G902), .ZN(n458) );
  XNOR2_X1 U452 ( .A(n408), .B(n407), .ZN(n533) );
  XNOR2_X1 U453 ( .A(KEYINPUT13), .B(G475), .ZN(n407) );
  NOR2_X1 U454 ( .A1(n702), .A2(G902), .ZN(n408) );
  INV_X1 U455 ( .A(n540), .ZN(n578) );
  XNOR2_X1 U456 ( .A(n491), .B(n419), .ZN(n611) );
  XNOR2_X1 U457 ( .A(n420), .B(n488), .ZN(n419) );
  XNOR2_X1 U458 ( .A(n507), .B(n378), .ZN(n420) );
  INV_X1 U459 ( .A(KEYINPUT83), .ZN(n398) );
  OR2_X1 U460 ( .A1(G902), .A2(G237), .ZN(n477) );
  XNOR2_X1 U461 ( .A(G110), .B(KEYINPUT92), .ZN(n499) );
  XOR2_X1 U462 ( .A(KEYINPUT24), .B(KEYINPUT84), .Z(n500) );
  XNOR2_X1 U463 ( .A(n502), .B(KEYINPUT23), .ZN(n406) );
  XNOR2_X1 U464 ( .A(G119), .B(G128), .ZN(n502) );
  XNOR2_X1 U465 ( .A(n498), .B(n402), .ZN(n729) );
  INV_X1 U466 ( .A(n510), .ZN(n402) );
  NAND2_X1 U467 ( .A1(n734), .A2(G234), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n371), .B(n546), .ZN(n604) );
  NAND2_X1 U469 ( .A1(G237), .A2(G234), .ZN(n479) );
  NAND2_X1 U470 ( .A1(n386), .A2(n385), .ZN(n389) );
  NAND2_X1 U471 ( .A1(n388), .A2(n437), .ZN(n387) );
  INV_X1 U472 ( .A(n655), .ZN(n388) );
  NAND2_X1 U473 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U474 ( .A1(n397), .A2(G902), .ZN(n395) );
  NAND2_X1 U475 ( .A1(n611), .A2(n397), .ZN(n396) );
  XNOR2_X1 U476 ( .A(n379), .B(n358), .ZN(n378) );
  XNOR2_X1 U477 ( .A(n489), .B(n380), .ZN(n379) );
  XNOR2_X1 U478 ( .A(G137), .B(KEYINPUT95), .ZN(n489) );
  XNOR2_X1 U479 ( .A(G110), .B(G104), .ZN(n464) );
  XNOR2_X1 U480 ( .A(n718), .B(n434), .ZN(n433) );
  XNOR2_X1 U481 ( .A(n435), .B(n474), .ZN(n434) );
  AND2_X1 U482 ( .A1(n605), .A2(n597), .ZN(n732) );
  NOR2_X1 U483 ( .A1(n583), .A2(n642), .ZN(n548) );
  OR2_X2 U484 ( .A1(n391), .A2(n394), .ZN(n648) );
  XNOR2_X1 U485 ( .A(n456), .B(n412), .ZN(n708) );
  XNOR2_X1 U486 ( .A(n455), .B(n413), .ZN(n412) );
  XNOR2_X1 U487 ( .A(n450), .B(n449), .ZN(n702) );
  XNOR2_X1 U488 ( .A(n509), .B(n370), .ZN(n511) );
  XNOR2_X1 U489 ( .A(n510), .B(n508), .ZN(n370) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n742) );
  INV_X1 U491 ( .A(KEYINPUT42), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n376), .B(n375), .ZN(n744) );
  INV_X1 U493 ( .A(KEYINPUT40), .ZN(n375) );
  AND2_X1 U494 ( .A1(n424), .A2(n423), .ZN(n631) );
  XNOR2_X1 U495 ( .A(n579), .B(KEYINPUT36), .ZN(n424) );
  INV_X1 U496 ( .A(KEYINPUT34), .ZN(n525) );
  XNOR2_X1 U497 ( .A(n515), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U498 ( .A1(n367), .A2(n366), .ZN(n515) );
  AND2_X1 U499 ( .A1(n357), .A2(n514), .ZN(n366) );
  NAND2_X1 U500 ( .A1(n361), .A2(n399), .ZN(n623) );
  NOR2_X1 U501 ( .A1(n583), .A2(n400), .ZN(n399) );
  NAND2_X1 U502 ( .A1(n431), .A2(n693), .ZN(n430) );
  XNOR2_X1 U503 ( .A(n432), .B(n364), .ZN(n431) );
  INV_X1 U504 ( .A(KEYINPUT120), .ZN(n414) );
  NAND2_X1 U505 ( .A1(n416), .A2(n693), .ZN(n415) );
  XNOR2_X1 U506 ( .A(n418), .B(n417), .ZN(n416) );
  AND2_X1 U507 ( .A1(n389), .A2(n387), .ZN(n355) );
  INV_X1 U508 ( .A(n641), .ZN(n423) );
  XOR2_X1 U509 ( .A(KEYINPUT80), .B(KEYINPUT90), .Z(n356) );
  XOR2_X1 U510 ( .A(KEYINPUT77), .B(n540), .Z(n357) );
  AND2_X1 U511 ( .A1(n490), .A2(G210), .ZN(n358) );
  XOR2_X1 U512 ( .A(n475), .B(n356), .Z(n359) );
  OR2_X1 U513 ( .A1(n391), .A2(n390), .ZN(n360) );
  INV_X1 U514 ( .A(n584), .ZN(n400) );
  AND2_X1 U515 ( .A1(n582), .A2(n581), .ZN(n361) );
  INV_X1 U516 ( .A(n494), .ZN(n397) );
  XNOR2_X1 U517 ( .A(n493), .B(n492), .ZN(n494) );
  OR2_X1 U518 ( .A1(n551), .A2(n483), .ZN(n362) );
  NAND2_X1 U519 ( .A1(n390), .A2(n655), .ZN(n363) );
  XOR2_X1 U520 ( .A(n611), .B(KEYINPUT62), .Z(n364) );
  XNOR2_X1 U521 ( .A(n488), .B(n469), .ZN(n718) );
  NOR2_X1 U522 ( .A1(G952), .A2(n734), .ZN(n712) );
  INV_X1 U523 ( .A(n516), .ZN(n367) );
  AND2_X1 U524 ( .A1(n567), .A2(n362), .ZN(n484) );
  NAND2_X1 U525 ( .A1(n369), .A2(n368), .ZN(n530) );
  INV_X1 U526 ( .A(KEYINPUT44), .ZN(n368) );
  NAND2_X1 U527 ( .A1(n545), .A2(n544), .ZN(n371) );
  NOR2_X2 U528 ( .A1(n580), .A2(n527), .ZN(n528) );
  XNOR2_X1 U529 ( .A(n732), .B(KEYINPUT73), .ZN(n598) );
  NAND2_X1 U530 ( .A1(n596), .A2(n626), .ZN(n376) );
  NAND2_X1 U531 ( .A1(n394), .A2(n363), .ZN(n382) );
  NAND2_X1 U532 ( .A1(n384), .A2(n360), .ZN(n383) );
  NOR2_X1 U533 ( .A1(n611), .A2(n392), .ZN(n391) );
  NOR2_X1 U534 ( .A1(n363), .A2(n392), .ZN(n385) );
  INV_X1 U535 ( .A(n611), .ZN(n386) );
  OR2_X2 U536 ( .A1(n642), .A2(n641), .ZN(n534) );
  NOR2_X2 U537 ( .A1(n705), .A2(n712), .ZN(n706) );
  XNOR2_X1 U538 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U539 ( .A(n415), .B(n414), .ZN(G66) );
  INV_X1 U540 ( .A(n711), .ZN(n417) );
  NAND2_X1 U541 ( .A1(n710), .A2(G217), .ZN(n418) );
  INV_X1 U542 ( .A(n648), .ZN(n535) );
  NAND2_X1 U543 ( .A1(n674), .A2(n568), .ZN(n429) );
  XNOR2_X2 U544 ( .A(n476), .B(n359), .ZN(n584) );
  XNOR2_X1 U545 ( .A(n430), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U546 ( .A1(n710), .A2(G472), .ZN(n432) );
  XNOR2_X1 U547 ( .A(n511), .B(n512), .ZN(n698) );
  NOR2_X2 U548 ( .A1(n600), .A2(n687), .ZN(n476) );
  XNOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n437) );
  XNOR2_X1 U550 ( .A(n518), .B(KEYINPUT86), .ZN(n519) );
  XNOR2_X1 U551 ( .A(n520), .B(n519), .ZN(n529) );
  INV_X1 U552 ( .A(KEYINPUT70), .ZN(n465) );
  INV_X1 U553 ( .A(n487), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n719), .B(n465), .ZN(n466) );
  INV_X1 U555 ( .A(KEYINPUT41), .ZN(n558) );
  INV_X1 U556 ( .A(KEYINPUT45), .ZN(n546) );
  XNOR2_X1 U557 ( .A(G902), .B(KEYINPUT15), .ZN(n461) );
  NAND2_X1 U558 ( .A1(n461), .A2(G234), .ZN(n438) );
  XNOR2_X1 U559 ( .A(n438), .B(KEYINPUT20), .ZN(n495) );
  NAND2_X1 U560 ( .A1(G221), .A2(n495), .ZN(n439) );
  XOR2_X1 U561 ( .A(KEYINPUT21), .B(n439), .Z(n638) );
  INV_X1 U562 ( .A(n638), .ZN(n560) );
  INV_X1 U563 ( .A(n498), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U565 ( .A(n443), .B(n442), .Z(n450) );
  NAND2_X1 U566 ( .A1(G214), .A2(n490), .ZN(n444) );
  XNOR2_X1 U567 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U568 ( .A(n446), .B(KEYINPUT98), .Z(n448) );
  XNOR2_X1 U569 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U570 ( .A(n533), .ZN(n459) );
  XNOR2_X2 U571 ( .A(G128), .B(KEYINPUT79), .ZN(n451) );
  XNOR2_X2 U572 ( .A(n451), .B(G143), .ZN(n462) );
  XNOR2_X1 U573 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n457) );
  NAND2_X1 U574 ( .A1(G217), .A2(n503), .ZN(n456) );
  XNOR2_X1 U575 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U576 ( .A(G478), .B(n458), .ZN(n532) );
  NAND2_X1 U577 ( .A1(n459), .A2(n532), .ZN(n659) );
  XNOR2_X1 U578 ( .A(KEYINPUT100), .B(n460), .ZN(n485) );
  INV_X1 U579 ( .A(n461), .ZN(n600) );
  XNOR2_X1 U580 ( .A(n464), .B(G107), .ZN(n719) );
  XNOR2_X1 U581 ( .A(G119), .B(G116), .ZN(n467) );
  XOR2_X1 U582 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n473) );
  NAND2_X1 U583 ( .A1(G224), .A2(n734), .ZN(n472) );
  XNOR2_X1 U584 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U585 ( .A1(G210), .A2(n477), .ZN(n475) );
  NAND2_X1 U586 ( .A1(G214), .A2(n477), .ZN(n655) );
  NAND2_X1 U587 ( .A1(n584), .A2(n655), .ZN(n478) );
  XNOR2_X1 U588 ( .A(n478), .B(KEYINPUT19), .ZN(n567) );
  XNOR2_X1 U589 ( .A(KEYINPUT14), .B(n479), .ZN(n481) );
  NAND2_X1 U590 ( .A1(n481), .A2(G952), .ZN(n480) );
  XOR2_X1 U591 ( .A(KEYINPUT91), .B(n480), .Z(n673) );
  NOR2_X1 U592 ( .A1(G953), .A2(n673), .ZN(n551) );
  AND2_X1 U593 ( .A1(G953), .A2(n481), .ZN(n482) );
  NAND2_X1 U594 ( .A1(G902), .A2(n482), .ZN(n549) );
  NOR2_X1 U595 ( .A1(G898), .A2(n549), .ZN(n483) );
  XNOR2_X2 U596 ( .A(n484), .B(KEYINPUT0), .ZN(n522) );
  NAND2_X1 U597 ( .A1(n485), .A2(n522), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n486), .B(KEYINPUT22), .ZN(n516) );
  XNOR2_X1 U599 ( .A(KEYINPUT97), .B(KEYINPUT71), .ZN(n493) );
  XOR2_X1 U600 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n497) );
  NAND2_X1 U601 ( .A1(n495), .A2(G217), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n497), .B(n496), .ZN(n506) );
  XNOR2_X1 U603 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U604 ( .A1(G221), .A2(n503), .ZN(n504) );
  NOR2_X1 U605 ( .A1(G902), .A2(n711), .ZN(n505) );
  XOR2_X1 U606 ( .A(n562), .B(KEYINPUT101), .Z(n637) );
  XOR2_X1 U607 ( .A(n507), .B(KEYINPUT74), .Z(n509) );
  NAND2_X1 U608 ( .A1(G227), .A2(n734), .ZN(n508) );
  NOR2_X1 U609 ( .A1(G902), .A2(n698), .ZN(n513) );
  NOR2_X1 U610 ( .A1(n637), .A2(n641), .ZN(n514) );
  NOR2_X1 U611 ( .A1(n648), .A2(n562), .ZN(n517) );
  NOR2_X1 U612 ( .A1(n516), .A2(n423), .ZN(n541) );
  NAND2_X1 U613 ( .A1(n517), .A2(n541), .ZN(n620) );
  NAND2_X1 U614 ( .A1(n747), .A2(n620), .ZN(n520) );
  NOR2_X1 U615 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n518) );
  INV_X1 U616 ( .A(n532), .ZN(n521) );
  NAND2_X1 U617 ( .A1(n533), .A2(n521), .ZN(n580) );
  INV_X1 U618 ( .A(n522), .ZN(n524) );
  XNOR2_X1 U619 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n523) );
  NAND2_X1 U620 ( .A1(n529), .A2(n745), .ZN(n531) );
  NAND2_X1 U621 ( .A1(n531), .A2(n530), .ZN(n545) );
  NAND2_X1 U622 ( .A1(n532), .A2(n533), .ZN(n576) );
  INV_X1 U623 ( .A(n576), .ZN(n626) );
  NOR2_X1 U624 ( .A1(n533), .A2(n532), .ZN(n628) );
  NOR2_X1 U625 ( .A1(n626), .A2(n628), .ZN(n661) );
  NOR2_X1 U626 ( .A1(n535), .A2(n534), .ZN(n651) );
  NAND2_X1 U627 ( .A1(n651), .A2(n522), .ZN(n536) );
  XNOR2_X1 U628 ( .A(KEYINPUT31), .B(n536), .ZN(n629) );
  AND2_X1 U629 ( .A1(n522), .A2(n548), .ZN(n537) );
  XOR2_X1 U630 ( .A(KEYINPUT94), .B(n537), .Z(n538) );
  NOR2_X1 U631 ( .A1(n648), .A2(n538), .ZN(n615) );
  NOR2_X1 U632 ( .A1(n629), .A2(n615), .ZN(n539) );
  NOR2_X1 U633 ( .A1(n661), .A2(n539), .ZN(n543) );
  NAND2_X1 U634 ( .A1(n541), .A2(n637), .ZN(n542) );
  NOR2_X1 U635 ( .A1(n578), .A2(n542), .ZN(n612) );
  NOR2_X1 U636 ( .A1(n543), .A2(n612), .ZN(n544) );
  INV_X1 U637 ( .A(KEYINPUT38), .ZN(n547) );
  NAND2_X1 U638 ( .A1(n656), .A2(n548), .ZN(n556) );
  XNOR2_X1 U639 ( .A(n549), .B(KEYINPUT102), .ZN(n550) );
  NOR2_X1 U640 ( .A1(G900), .A2(n550), .ZN(n552) );
  NOR2_X1 U641 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U642 ( .A(n553), .B(KEYINPUT81), .Z(n559) );
  INV_X1 U643 ( .A(n582), .ZN(n555) );
  OR2_X1 U644 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U645 ( .A1(n562), .A2(n561), .ZN(n574) );
  AND2_X1 U646 ( .A1(n648), .A2(n574), .ZN(n564) );
  XNOR2_X1 U647 ( .A(KEYINPUT28), .B(KEYINPUT105), .ZN(n563) );
  XNOR2_X1 U648 ( .A(n564), .B(n563), .ZN(n565) );
  NOR2_X1 U649 ( .A1(n565), .A2(n583), .ZN(n568) );
  INV_X1 U650 ( .A(KEYINPUT72), .ZN(n573) );
  NOR2_X1 U651 ( .A1(n573), .A2(KEYINPUT47), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U653 ( .A(KEYINPUT78), .B(n569), .Z(n624) );
  INV_X1 U654 ( .A(n661), .ZN(n570) );
  NAND2_X1 U655 ( .A1(n624), .A2(n570), .ZN(n571) );
  XNOR2_X1 U656 ( .A(n572), .B(n571), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n573), .A2(KEYINPUT47), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n574), .A2(n655), .ZN(n575) );
  NOR2_X1 U659 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n592) );
  NOR2_X1 U661 ( .A1(n400), .A2(n592), .ZN(n579) );
  NOR2_X1 U662 ( .A1(n642), .A2(n580), .ZN(n581) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n591), .B(n590), .ZN(n605) );
  XNOR2_X1 U665 ( .A(KEYINPUT103), .B(n592), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n593), .A2(n641), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT43), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n595), .A2(n400), .ZN(n636) );
  NAND2_X1 U669 ( .A1(n628), .A2(n596), .ZN(n634) );
  AND2_X1 U670 ( .A1(n636), .A2(n634), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n604), .A2(n598), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n599), .A2(n600), .ZN(n603) );
  NAND2_X1 U673 ( .A1(KEYINPUT2), .A2(n600), .ZN(n601) );
  XNOR2_X1 U674 ( .A(n601), .B(KEYINPUT64), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(n610) );
  INV_X1 U676 ( .A(n604), .ZN(n713) );
  NAND2_X1 U677 ( .A1(n605), .A2(n636), .ZN(n608) );
  NAND2_X1 U678 ( .A1(KEYINPUT2), .A2(n634), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT82), .B(n606), .ZN(n607) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n713), .A2(n609), .ZN(n681) );
  XOR2_X1 U682 ( .A(G101), .B(n612), .Z(G3) );
  NAND2_X1 U683 ( .A1(n615), .A2(n626), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT106), .ZN(n614) );
  XNOR2_X1 U685 ( .A(G104), .B(n614), .ZN(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n617) );
  NAND2_X1 U687 ( .A1(n615), .A2(n628), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(G107), .B(n618), .ZN(G9) );
  XOR2_X1 U690 ( .A(G110), .B(KEYINPUT107), .Z(n619) );
  XNOR2_X1 U691 ( .A(n620), .B(n619), .ZN(G12) );
  XOR2_X1 U692 ( .A(G128), .B(KEYINPUT29), .Z(n622) );
  NAND2_X1 U693 ( .A1(n628), .A2(n624), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(G30) );
  XNOR2_X1 U695 ( .A(G143), .B(n623), .ZN(G45) );
  NAND2_X1 U696 ( .A1(n624), .A2(n626), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n625), .B(G146), .ZN(G48) );
  NAND2_X1 U698 ( .A1(n629), .A2(n626), .ZN(n627) );
  XNOR2_X1 U699 ( .A(n627), .B(G113), .ZN(G15) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(G116), .ZN(G18) );
  XNOR2_X1 U702 ( .A(n631), .B(KEYINPUT108), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT37), .ZN(n633) );
  XNOR2_X1 U704 ( .A(G125), .B(n633), .ZN(G27) );
  INV_X1 U705 ( .A(n634), .ZN(n635) );
  XOR2_X1 U706 ( .A(G134), .B(n635), .Z(G36) );
  XNOR2_X1 U707 ( .A(G140), .B(n636), .ZN(G42) );
  NOR2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U709 ( .A(KEYINPUT49), .B(n639), .Z(n640) );
  XNOR2_X1 U710 ( .A(KEYINPUT109), .B(n640), .ZN(n646) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT50), .ZN(n644) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(n644), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U716 ( .A(KEYINPUT111), .B(n649), .Z(n650) );
  NOR2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U718 ( .A(n652), .B(KEYINPUT51), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT112), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n654), .A2(n674), .ZN(n669) );
  NOR2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U722 ( .A(KEYINPUT113), .B(n657), .Z(n658) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U724 ( .A(n660), .B(KEYINPUT114), .ZN(n664) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n665), .Z(n666) );
  NOR2_X1 U728 ( .A1(n676), .A2(n666), .ZN(n667) );
  XOR2_X1 U729 ( .A(KEYINPUT116), .B(n667), .Z(n668) );
  NAND2_X1 U730 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U731 ( .A(n670), .B(KEYINPUT117), .ZN(n671) );
  XNOR2_X1 U732 ( .A(n671), .B(KEYINPUT52), .ZN(n672) );
  NOR2_X1 U733 ( .A1(n673), .A2(n672), .ZN(n678) );
  INV_X1 U734 ( .A(n674), .ZN(n675) );
  NOR2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n684) );
  NAND2_X1 U737 ( .A1(n713), .A2(n732), .ZN(n680) );
  INV_X1 U738 ( .A(KEYINPUT2), .ZN(n679) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U742 ( .A1(n685), .A2(G953), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n686), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U744 ( .A(n712), .ZN(n693) );
  NAND2_X1 U745 ( .A1(n710), .A2(G210), .ZN(n691) );
  XOR2_X1 U746 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n689) );
  XNOR2_X1 U747 ( .A(n687), .B(KEYINPUT87), .ZN(n688) );
  XNOR2_X1 U748 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U750 ( .A(KEYINPUT56), .B(n694), .ZN(G51) );
  XOR2_X1 U751 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n696) );
  XNOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n695) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(n697) );
  XOR2_X1 U754 ( .A(n698), .B(n697), .Z(n700) );
  NAND2_X1 U755 ( .A1(n710), .A2(G469), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n712), .A2(n701), .ZN(G54) );
  XOR2_X1 U758 ( .A(n702), .B(KEYINPUT59), .Z(n704) );
  NAND2_X1 U759 ( .A1(n710), .A2(G475), .ZN(n703) );
  XNOR2_X1 U760 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U762 ( .A1(G478), .A2(n710), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n712), .A2(n709), .ZN(G63) );
  NAND2_X1 U765 ( .A1(n734), .A2(n713), .ZN(n717) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n714) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n714), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n715), .A2(G898), .ZN(n716) );
  NAND2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n724) );
  XOR2_X1 U770 ( .A(G101), .B(n719), .Z(n720) );
  XNOR2_X1 U771 ( .A(n718), .B(n720), .ZN(n722) );
  NOR2_X1 U772 ( .A1(G898), .A2(n734), .ZN(n721) );
  NOR2_X1 U773 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U774 ( .A(n724), .B(n723), .ZN(n725) );
  XOR2_X1 U775 ( .A(KEYINPUT121), .B(n725), .Z(G69) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n726) );
  XNOR2_X1 U777 ( .A(n727), .B(n726), .ZN(n728) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n730), .B(n731), .ZN(n736) );
  XOR2_X1 U780 ( .A(n732), .B(KEYINPUT124), .Z(n733) );
  XNOR2_X1 U781 ( .A(n736), .B(n733), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n741) );
  XNOR2_X1 U783 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(G900), .ZN(n738) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n738), .Z(n739) );
  NAND2_X1 U786 ( .A1(G953), .A2(n739), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G137), .B(KEYINPUT127), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(n742), .ZN(G39) );
  XOR2_X1 U790 ( .A(n744), .B(G131), .Z(G33) );
  XNOR2_X1 U791 ( .A(G122), .B(KEYINPUT126), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n746), .B(n745), .ZN(G24) );
  XNOR2_X1 U793 ( .A(G119), .B(n747), .ZN(G21) );
endmodule

