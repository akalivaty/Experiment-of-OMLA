//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n461), .B2(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n467), .B1(new_n470), .B2(new_n462), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n468), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n471), .B2(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n473), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2105), .B1(KEYINPUT68), .B2(G114), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT68), .A2(G114), .ZN(new_n490));
  OAI211_X1 g065(.A(G2104), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n461), .A2(G138), .A3(new_n462), .A4(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n462), .C1(new_n472), .C2(new_n473), .ZN(new_n497));
  INV_X1    g072(.A(new_n495), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n496), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n508), .A2(G50), .B1(G651), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(new_n507), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n502), .A2(new_n505), .B1(KEYINPUT6), .B2(new_n501), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT71), .A3(new_n516), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n508), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n526), .B(new_n531), .C1(new_n522), .C2(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND3_X1  g109(.A1(new_n519), .A2(G90), .A3(new_n521), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n512), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n508), .A2(G52), .B1(G651), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n535), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND3_X1  g116(.A1(new_n519), .A2(G81), .A3(new_n521), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n512), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n508), .A2(G43), .B1(G651), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT72), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n506), .A2(G543), .A3(new_n507), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n520), .A2(KEYINPUT73), .A3(G53), .A4(G543), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n555), .B(new_n561), .C1(new_n556), .C2(new_n557), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  INV_X1    g139(.A(G543), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n512), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n568), .B1(new_n564), .B2(new_n565), .C1(new_n512), .C2(new_n563), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(G651), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n519), .A2(G91), .A3(new_n521), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n560), .A2(new_n562), .A3(new_n570), .A4(new_n571), .ZN(G299));
  NAND3_X1  g147(.A1(new_n519), .A2(G87), .A3(new_n521), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n516), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n508), .A2(G49), .B1(new_n574), .B2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n519), .A2(G86), .A3(new_n521), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n512), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n508), .A2(G48), .B1(G651), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G305));
  NAND3_X1  g157(.A1(new_n519), .A2(G85), .A3(new_n521), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n512), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n508), .A2(G47), .B1(G651), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n519), .A2(G92), .A3(new_n521), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n519), .A2(new_n592), .A3(new_n521), .A4(G92), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n512), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n556), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n591), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n548), .ZN(G323));
  XOR2_X1   g188(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n614));
  XNOR2_X1  g189(.A(G323), .B(new_n614), .ZN(G282));
  NAND2_X1  g190(.A1(new_n461), .A2(new_n464), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n482), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n480), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n462), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT76), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT79), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT78), .B(G2438), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(new_n632), .ZN(new_n637));
  INV_X1    g212(.A(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n658), .A2(new_n653), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n655), .ZN(new_n661));
  INV_X1    g236(.A(new_n654), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n653), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n671), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n671), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT82), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n675), .B(KEYINPUT20), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n684));
  NAND4_X1  g259(.A1(new_n683), .A2(new_n684), .A3(new_n680), .A4(new_n679), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n668), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n682), .A2(new_n685), .A3(new_n668), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n690), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n688), .B1(new_n692), .B2(new_n686), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT83), .B(G16), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n705), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G6), .A2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G305), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(G16), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n713), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(KEYINPUT34), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT34), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n713), .A2(new_n720), .A3(new_n725), .A4(new_n721), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n701), .A2(G24), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n583), .A2(new_n587), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n701), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n482), .A2(G131), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n480), .A2(G119), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n462), .A2(G107), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  MUX2_X1   g310(.A(G25), .B(new_n735), .S(G29), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT35), .B(G1991), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n699), .B1(new_n724), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n723), .A2(new_n726), .A3(new_n740), .A4(new_n698), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G27), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT97), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n499), .A2(new_n496), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n491), .A2(new_n492), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n747), .B1(new_n750), .B2(G29), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT98), .Z(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NOR2_X1   g328(.A1(G5), .A2(G16), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT96), .Z(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G301), .B2(new_n706), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n752), .A2(G2078), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n548), .B2(new_n700), .ZN(new_n759));
  INV_X1    g334(.A(G1966), .ZN(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n706), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n706), .B2(G21), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n757), .B1(G1341), .B2(new_n759), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n760), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n745), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n482), .A2(G139), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT88), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(new_n462), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT25), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n775), .A2(new_n776), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n767), .B1(new_n780), .B2(new_n745), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n766), .B1(new_n781), .B2(G2072), .ZN(new_n782));
  OR3_X1    g357(.A1(new_n781), .A2(new_n766), .A3(G2072), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n763), .B(new_n765), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT30), .B(G28), .ZN(new_n785));
  OR2_X1    g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  NAND2_X1  g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n785), .A2(new_n745), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n626), .B2(new_n745), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G35), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G162), .B2(G29), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n793));
  INV_X1    g368(.A(G2090), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n792), .B(new_n795), .Z(new_n796));
  INV_X1    g371(.A(G2084), .ZN(new_n797));
  NAND2_X1  g372(.A1(G160), .A2(G29), .ZN(new_n798));
  AND2_X1   g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NOR2_X1   g374(.A1(KEYINPUT24), .A2(G34), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n745), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT91), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n790), .B(new_n796), .C1(new_n797), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n753), .B2(new_n756), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n781), .A2(G2072), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n482), .A2(G140), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n480), .A2(G128), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n462), .A2(G116), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n807), .B(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G29), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n745), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT87), .ZN(new_n816));
  INV_X1    g391(.A(G2067), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n752), .A2(G2078), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n759), .A2(G1341), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n806), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n700), .A2(G20), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT100), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT23), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n606), .B2(new_n706), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n803), .A2(new_n797), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n745), .A2(G32), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n480), .A2(G129), .ZN(new_n830));
  NAND3_X1  g405(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT26), .Z(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n828), .B1(new_n837), .B2(new_n745), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT27), .B(G1996), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT93), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n827), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n840), .B2(new_n838), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n805), .A2(new_n821), .A3(new_n826), .A4(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(G4), .A2(G16), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n602), .B2(G16), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT86), .ZN(new_n846));
  INV_X1    g421(.A(G1348), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND4_X1   g423(.A1(new_n744), .A2(new_n784), .A3(new_n843), .A4(new_n848), .ZN(G311));
  NAND4_X1  g424(.A1(new_n744), .A2(new_n784), .A3(new_n843), .A4(new_n848), .ZN(G150));
  NAND3_X1  g425(.A1(new_n519), .A2(G93), .A3(new_n521), .ZN(new_n851));
  OAI21_X1  g426(.A(G67), .B1(new_n510), .B2(new_n511), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n501), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n508), .B2(G55), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n602), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n547), .A2(new_n856), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n542), .A2(new_n851), .A3(new_n546), .A4(new_n855), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n860), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n858), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(G145));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n493), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n748), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n835), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n748), .A2(new_n876), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n834), .A2(new_n881), .A3(new_n835), .A4(new_n875), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n811), .B(KEYINPUT103), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n873), .B(new_n780), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n882), .ZN(new_n887));
  INV_X1    g462(.A(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT104), .B1(new_n778), .B2(new_n779), .ZN(new_n890));
  INV_X1    g465(.A(new_n779), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n873), .A3(new_n777), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n889), .A2(new_n890), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n482), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n480), .A2(G130), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n462), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n900), .B(new_n617), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n735), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n886), .A2(new_n894), .A3(new_n902), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G162), .B(new_n626), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G160), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G37), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n886), .A2(new_n894), .A3(new_n902), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n902), .B1(new_n886), .B2(new_n894), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT105), .B1(new_n913), .B2(new_n908), .ZN(new_n914));
  AND4_X1   g489(.A1(KEYINPUT105), .A2(new_n904), .A3(new_n908), .A4(new_n905), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g492(.A(G868), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n856), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(G288), .A2(G290), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n922));
  NAND2_X1  g497(.A1(G288), .A2(G290), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT107), .B1(new_n925), .B2(new_n920), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n715), .B(G303), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(G303), .B(G305), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n922), .A3(new_n923), .A4(new_n921), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n931), .A2(KEYINPUT108), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n930), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(KEYINPUT108), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n601), .A2(G299), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n601), .A2(G299), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n611), .B(new_n863), .Z(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT41), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n941), .B2(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n602), .A2(new_n606), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n940), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n947), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n939), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n919), .B1(new_n955), .B2(new_n918), .ZN(G295));
  OAI21_X1  g531(.A(new_n919), .B1(new_n955), .B2(new_n918), .ZN(G331));
  AOI21_X1  g532(.A(G286), .B1(G171), .B2(KEYINPUT109), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n960));
  NAND2_X1  g535(.A1(G301), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n861), .A2(new_n961), .A3(new_n862), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n861), .B2(new_n862), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT109), .B1(new_n535), .B2(new_n539), .ZN(new_n966));
  AND4_X1   g541(.A1(new_n542), .A2(new_n851), .A3(new_n546), .A4(new_n855), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n542), .A2(new_n546), .B1(new_n851), .B2(new_n855), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n962), .A3(new_n958), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n943), .A3(new_n970), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n969), .A2(new_n962), .A3(new_n958), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n958), .B1(new_n969), .B2(new_n962), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n974), .B2(new_n952), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(new_n934), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n975), .B2(new_n934), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(KEYINPUT110), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n949), .B(new_n951), .C1(new_n972), .C2(new_n973), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n931), .B1(new_n980), .B2(new_n971), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n981), .B2(G37), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT43), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n945), .A2(new_n974), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n931), .B1(new_n984), .B2(new_n980), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n985), .A2(new_n976), .A3(new_n986), .A4(G37), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT44), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n978), .B2(new_n982), .ZN(new_n990));
  NOR4_X1   g565(.A1(new_n985), .A2(new_n976), .A3(KEYINPUT43), .A4(G37), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(G397));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n877), .A2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n995), .B2(KEYINPUT111), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n466), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n467), .B(new_n462), .C1(new_n474), .C2(new_n468), .ZN(new_n1001));
  OAI211_X1 g576(.A(G40), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n811), .B(new_n817), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n836), .B2(G1996), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n836), .A2(G1996), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT112), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OR4_X1    g584(.A1(KEYINPUT112), .A2(new_n998), .A3(new_n1008), .A4(new_n1002), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n735), .B(new_n738), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT113), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1003), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G290), .B(G1986), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1003), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n750), .B2(new_n994), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n1002), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n994), .A2(KEYINPUT45), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT114), .B1(new_n877), .B2(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n877), .A2(KEYINPUT114), .A3(new_n1021), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1019), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1956), .ZN(new_n1025));
  INV_X1    g600(.A(G40), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1026), .B(new_n466), .C1(new_n471), .C2(new_n476), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n748), .B2(new_n749), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n877), .B2(new_n994), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1025), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1024), .A2(new_n1033), .ZN(new_n1034));
  OR2_X1    g609(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n877), .A2(new_n1029), .A3(new_n994), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1027), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n995), .A2(new_n1002), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1041), .A2(new_n847), .B1(new_n1042), .B2(new_n817), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n1043), .B2(new_n601), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1028), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1002), .B1(new_n1046), .B2(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1348), .B1(new_n1047), .B2(new_n1039), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n995), .A2(new_n1002), .A3(G2067), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1045), .B(new_n602), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1038), .A2(new_n1044), .A3(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1024), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(KEYINPUT120), .A3(new_n1052), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1043), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n601), .B1(new_n1043), .B2(KEYINPUT60), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1057), .A2(new_n1058), .B1(KEYINPUT60), .B2(new_n1043), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n877), .A2(new_n1021), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n877), .A2(KEYINPUT114), .A3(new_n1021), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1996), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n1019), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n995), .B2(new_n1002), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n548), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1072), .B2(new_n548), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1059), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT61), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1052), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1024), .A2(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1038), .A2(KEYINPUT61), .A3(new_n1052), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1055), .B(new_n1056), .C1(new_n1076), .C2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n573), .A2(new_n575), .A3(G1976), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1084), .B(G8), .C1(new_n995), .C2(new_n1002), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(KEYINPUT115), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n995), .B2(new_n1002), .ZN(new_n1092));
  INV_X1    g667(.A(G1981), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n577), .A2(new_n581), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n577), .B2(new_n581), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1096), .B2(KEYINPUT49), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT116), .B(new_n1098), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1097), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1086), .A2(new_n1104), .A3(new_n1088), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1091), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(G303), .A2(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1971), .B1(new_n1064), .B2(new_n1019), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1041), .A2(G2090), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1109), .B(G8), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1032), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(new_n794), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1115));
  OAI211_X1 g690(.A(G160), .B(G40), .C1(KEYINPUT45), .C2(new_n1028), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1117), .B2(G1971), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1113), .B(new_n1109), .C1(new_n1118), .C2(G8), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1031), .A2(G2090), .A3(new_n1032), .ZN(new_n1120));
  OAI21_X1  g695(.A(G8), .B1(new_n1110), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1109), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT117), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1106), .B(new_n1112), .C1(new_n1119), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1064), .A2(new_n1019), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(G2078), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n750), .A2(new_n1021), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(G160), .A3(G40), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT45), .B1(new_n877), .B2(new_n994), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1125), .A2(G2078), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1041), .A2(new_n753), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1127), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(G301), .B(KEYINPUT54), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1138));
  OAI21_X1  g713(.A(new_n760), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1039), .A2(new_n1027), .A3(new_n797), .A4(new_n1040), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G286), .A2(G8), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT123), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n1144));
  NAND3_X1  g719(.A1(G286), .A2(new_n1144), .A3(G8), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(G8), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G8), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(G286), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1138), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1141), .A2(G8), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1142), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n475), .A2(G2105), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n999), .A2(G40), .A3(new_n1153), .A4(new_n1132), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1136), .B1(new_n998), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1127), .A2(new_n1156), .A3(new_n1134), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1137), .A2(new_n1149), .A3(new_n1152), .A4(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1124), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1083), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1091), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G288), .A2(G1976), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1094), .B1(new_n1103), .B2(new_n1162), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1161), .A2(new_n1112), .B1(new_n1163), .B2(new_n1092), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1148), .B(KEYINPUT118), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1122), .B1(new_n1166), .B2(new_n1147), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1106), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1168), .B2(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1160), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1149), .A2(KEYINPUT62), .A3(new_n1152), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1173), .A2(G171), .A3(new_n1174), .A4(new_n1135), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1165), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1124), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1017), .B1(new_n1170), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n1180));
  INV_X1    g755(.A(G1986), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1003), .A2(new_n1181), .A3(new_n728), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT48), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1183), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1003), .A2(KEYINPUT46), .A3(new_n1065), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT124), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1003), .A2(new_n1187), .A3(KEYINPUT46), .A4(new_n1065), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(KEYINPUT46), .B1(new_n1003), .B2(new_n1065), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n837), .A2(new_n1004), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1003), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT47), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1184), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n735), .A2(new_n738), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1011), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n811), .A2(G2067), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1007), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1180), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT47), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1189), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1197), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n1207), .B(new_n1006), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1003), .B1(new_n1208), .B2(new_n1199), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1206), .A2(new_n1209), .A3(KEYINPUT125), .A4(new_n1184), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1202), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1179), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g787(.A1(G227), .A2(new_n459), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1214), .B1(new_n649), .B2(new_n651), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n1215), .B1(new_n695), .B2(new_n696), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(KEYINPUT126), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n1215), .B(new_n1218), .C1(new_n695), .C2(new_n696), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g794(.A(new_n916), .B(new_n1220), .C1(new_n990), .C2(new_n991), .ZN(G225));
  INV_X1    g795(.A(G225), .ZN(G308));
endmodule


