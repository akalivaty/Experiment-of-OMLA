//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n548, new_n550, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT65), .B(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(KEYINPUT65), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n468), .B(G2104), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n467), .A2(new_n462), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n463), .B(new_n464), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  INV_X1    g055(.A(G136), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n467), .A2(G2105), .A3(new_n473), .A4(new_n474), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n480), .B1(new_n475), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n485), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n475), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n460), .A2(new_n498), .A3(G138), .A4(new_n462), .ZN(new_n499));
  XNOR2_X1  g074(.A(new_n499), .B(KEYINPUT68), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G62), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  INV_X1    g092(.A(new_n506), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n518), .A3(new_n514), .ZN(new_n519));
  OAI221_X1 g094(.A(new_n509), .B1(new_n515), .B2(new_n516), .C1(new_n517), .C2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n515), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n510), .ZN(new_n534));
  INV_X1    g109(.A(new_n519), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n510), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(G81), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT71), .B(G43), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n528), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT72), .Z(G188));
  AND2_X1   g128(.A1(new_n513), .A2(new_n514), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n554), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n515), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n556), .A2(new_n558), .B1(G91), .B2(new_n535), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n506), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G651), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n559), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n535), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n528), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n506), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(KEYINPUT75), .A3(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n519), .A2(new_n582), .B1(new_n515), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n510), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT76), .B(G85), .Z(new_n589));
  NAND2_X1  g164(.A1(new_n535), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n528), .A2(G47), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n506), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT10), .B1(new_n519), .B2(new_n601), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G280));
  XNOR2_X1  g186(.A(KEYINPUT78), .B(G559), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(G860), .B2(new_n605), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(G148));
  INV_X1    g190(.A(new_n613), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n622), .B(new_n623), .C1(G111), .C2(new_n462), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n475), .B2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n483), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT13), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT15), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2435), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2435), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n646), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n638), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n637), .A3(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n656), .A3(G14), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT83), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n677), .A2(new_n681), .A3(new_n684), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  INV_X1    g267(.A(G1981), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n585), .B2(new_n697), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT88), .B1(G16), .B2(G23), .ZN(new_n708));
  OR3_X1    g283(.A1(KEYINPUT88), .A2(G16), .A3(G23), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n708), .B(new_n709), .C1(G288), .C2(new_n697), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  OR3_X1    g288(.A1(new_n702), .A2(new_n703), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n703), .B1(new_n702), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G25), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G131), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n462), .A2(G107), .ZN(new_n720));
  OAI22_X1  g295(.A1(new_n475), .A2(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G119), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT87), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT35), .B(G1991), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G24), .B(G290), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1986), .Z(new_n731));
  NAND3_X1  g306(.A1(new_n716), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT36), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n716), .A2(new_n734), .A3(new_n729), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n697), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n697), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2090), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n743), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n741), .A2(G26), .ZN(new_n747));
  OR2_X1    g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n749));
  INV_X1    g324(.A(G140), .ZN(new_n750));
  INV_X1    g325(.A(G128), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n749), .B1(new_n475), .B2(new_n750), .C1(new_n751), .C2(new_n483), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n747), .B1(new_n756), .B2(new_n741), .ZN(new_n757));
  MUX2_X1   g332(.A(new_n747), .B(new_n757), .S(KEYINPUT28), .Z(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G2067), .ZN(new_n759));
  NAND2_X1  g334(.A1(G164), .A2(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G27), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2078), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n758), .A2(G2067), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n759), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n768));
  INV_X1    g343(.A(G20), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G16), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n770), .C1(new_n609), .C2(new_n697), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT95), .B(G1956), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT24), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n774), .A2(new_n741), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G160), .B2(new_n741), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT31), .B(G11), .Z(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G28), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n780), .B(new_n783), .C1(new_n629), .C2(G29), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(new_n462), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  INV_X1    g363(.A(G139), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n788), .C1(new_n475), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2072), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n773), .A2(new_n779), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G29), .A2(G32), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT26), .Z(new_n797));
  INV_X1    g372(.A(G141), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n795), .B(new_n797), .C1(new_n475), .C2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G129), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n483), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n799), .A2(KEYINPUT92), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n794), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT27), .B(G1996), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n605), .A2(G16), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G4), .B2(G16), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT90), .B(G1348), .Z(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G1341), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n546), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G16), .B2(G19), .ZN(new_n817));
  NOR2_X1   g392(.A1(G5), .A2(G16), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G171), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(G1961), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n815), .A2(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n811), .A2(new_n813), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n817), .A2(new_n815), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n814), .A2(new_n822), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n766), .A2(new_n793), .A3(new_n809), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n736), .A2(new_n740), .A3(new_n746), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n820), .A2(new_n821), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(G311));
  OR2_X1    g404(.A1(new_n827), .A2(new_n828), .ZN(G150));
  XNOR2_X1  g405(.A(KEYINPUT98), .B(G55), .ZN(new_n831));
  AOI22_X1  g406(.A1(G93), .A2(new_n535), .B1(new_n528), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n506), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT97), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(KEYINPUT97), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(G651), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n545), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n605), .A2(G559), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT39), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n844), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n841), .B1(new_n847), .B2(G860), .ZN(G145));
  INV_X1    g423(.A(G37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n756), .A2(G164), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n754), .A2(new_n755), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n497), .A2(new_n500), .ZN(new_n852));
  INV_X1    g427(.A(new_n495), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n790), .B1(new_n804), .B2(new_n805), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n803), .A2(new_n790), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n850), .B(new_n855), .C1(new_n857), .C2(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n865));
  INV_X1    g440(.A(G142), .ZN(new_n866));
  INV_X1    g441(.A(G130), .ZN(new_n867));
  OAI221_X1 g442(.A(new_n865), .B1(new_n475), .B2(new_n866), .C1(new_n867), .C2(new_n483), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n724), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n633), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n486), .A2(KEYINPUT99), .A3(new_n487), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n486), .B2(new_n487), .ZN(new_n875));
  OAI21_X1  g450(.A(G160), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n488), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n477), .A3(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n629), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n879), .ZN(new_n881));
  INV_X1    g456(.A(new_n629), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n861), .A2(new_n862), .A3(new_n870), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n872), .A2(new_n880), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n871), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n863), .A2(new_n888), .B1(new_n883), .B2(new_n880), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n861), .A2(new_n871), .A3(new_n862), .A4(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n863), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(new_n880), .ZN(new_n893));
  AND4_X1   g468(.A1(new_n886), .A2(new_n892), .A3(new_n893), .A4(new_n890), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n849), .B(new_n885), .C1(new_n891), .C2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g471(.A1(new_n839), .A2(G868), .ZN(new_n897));
  INV_X1    g472(.A(G288), .ZN(new_n898));
  NAND2_X1  g473(.A1(G290), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(G288), .B(new_n588), .C1(new_n593), .C2(new_n594), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n585), .B(G303), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(KEYINPUT103), .A3(new_n900), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n903), .B2(new_n904), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n842), .B(new_n616), .ZN(new_n914));
  NAND3_X1  g489(.A1(G299), .A2(KEYINPUT102), .A3(new_n604), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n559), .A2(new_n567), .A3(new_n564), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n567), .B1(new_n559), .B2(new_n564), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT102), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n566), .A2(new_n919), .A3(new_n568), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n920), .A3(new_n605), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n914), .A2(new_n915), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n915), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n928), .B2(new_n914), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n912), .A2(new_n913), .A3(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n913), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n912), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n897), .B1(new_n932), .B2(G868), .ZN(G295));
  AOI21_X1  g508(.A(new_n897), .B1(new_n932), .B2(G868), .ZN(G331));
  INV_X1    g509(.A(new_n907), .ZN(new_n935));
  NAND2_X1  g510(.A1(G286), .A2(G171), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(G301), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n936), .A2(new_n842), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n842), .B1(new_n936), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n926), .B2(new_n927), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n924), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n915), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT41), .B1(new_n921), .B2(new_n915), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n945), .A2(new_n946), .B1(new_n938), .B2(new_n939), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n907), .A3(new_n942), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n849), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n944), .A2(new_n951), .A3(new_n948), .A4(new_n849), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n952), .A2(KEYINPUT107), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(KEYINPUT44), .A3(new_n950), .A4(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n958), .ZN(G397));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n851), .B(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1996), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n806), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n961), .B(new_n963), .C1(new_n962), .C2(new_n802), .ZN(new_n964));
  XOR2_X1   g539(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G164), .B2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(G40), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n477), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT111), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n728), .A3(new_n725), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n756), .A2(new_n960), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n972), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n971), .B1(new_n961), .B2(new_n802), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n979), .B(KEYINPUT126), .Z(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n962), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n724), .B(new_n728), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n972), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n974), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n971), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT48), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n978), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT68), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n499), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n471), .A2(KEYINPUT65), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n468), .B1(new_n998), .B2(G2104), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT66), .B(new_n466), .C1(new_n996), .C2(new_n997), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1001), .A2(G138), .A3(new_n462), .A4(new_n474), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n995), .B1(new_n1002), .B2(KEYINPUT4), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n993), .C1(new_n1003), .C2(new_n495), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n967), .A2(new_n1004), .A3(new_n970), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n701), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n477), .A2(new_n969), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1384), .B1(new_n852), .B2(new_n853), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(G2090), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1007), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(G8), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n584), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n577), .B1(new_n584), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g605(.A(G1981), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n585), .A2(new_n693), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT118), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  AOI211_X1 g610(.A(KEYINPUT118), .B(new_n1035), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1009), .A2(new_n970), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(G8), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1037), .B2(G8), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1034), .A2(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n898), .A2(G1976), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT52), .B1(G288), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1043), .B(new_n1045), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1041), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1048), .A2(new_n1039), .B1(G1976), .B2(new_n898), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1042), .B(new_n1046), .C1(new_n1047), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1027), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1042), .A2(new_n1044), .A3(new_n898), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1032), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1053), .A2(new_n1054), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1026), .A2(KEYINPUT63), .A3(new_n1051), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1025), .B1(new_n1017), .B2(G8), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(G164), .B2(G1384), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n854), .A2(new_n993), .A3(new_n965), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n970), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n739), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1011), .A2(new_n1012), .A3(new_n778), .A4(new_n1014), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G168), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1056), .A2(new_n1057), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1052), .B(new_n1055), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  OAI211_X1 g644(.A(G168), .B(new_n1065), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT123), .ZN(new_n1074));
  NAND2_X1  g649(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1077), .A2(G8), .A3(G286), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1065), .A2(KEYINPUT51), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(G168), .A3(new_n1074), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT62), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n967), .A2(new_n1004), .A3(new_n762), .A4(new_n970), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1015), .A2(new_n821), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(G2078), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1060), .A2(new_n1061), .A3(new_n970), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1077), .A2(G8), .A3(G286), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1063), .A2(new_n1064), .A3(KEYINPUT123), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT123), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1075), .B1(new_n1095), .B2(G168), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1091), .B(new_n1092), .C1(new_n1096), .C2(new_n1079), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1082), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n1010), .A3(new_n993), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1100), .A3(new_n970), .ZN(new_n1101));
  INV_X1    g676(.A(G1956), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n565), .B(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n967), .A2(new_n1004), .A3(new_n970), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1110), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(G1956), .B1(new_n1011), .B2(new_n1099), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n967), .A2(new_n1004), .A3(new_n970), .A4(new_n1106), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT120), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1105), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1103), .A2(new_n1117), .A3(new_n1107), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT121), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .A4(new_n1116), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1037), .A2(G2067), .ZN(new_n1124));
  INV_X1    g699(.A(G1348), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1015), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1126), .A2(new_n604), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1112), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1116), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1109), .A2(new_n1111), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n967), .A2(new_n1004), .A3(new_n962), .A4(new_n970), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1037), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT122), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1138), .A3(new_n1135), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1139), .A3(new_n546), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .A4(new_n546), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1126), .A2(KEYINPUT60), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1015), .A2(new_n1125), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1124), .ZN(new_n1147));
  AND4_X1   g722(.A1(KEYINPUT60), .A2(new_n1146), .A3(new_n604), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n604), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1132), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1128), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1015), .A2(new_n821), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1154), .A2(G301), .A3(new_n1155), .A4(new_n1087), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n967), .A2(new_n1004), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT124), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n463), .A2(G40), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(new_n1086), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1154), .A2(new_n1162), .A3(new_n1155), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G171), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1085), .A2(new_n1165), .A3(G301), .A4(new_n1087), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1157), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1167), .A2(KEYINPUT54), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1163), .A2(G171), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1090), .A2(KEYINPUT54), .A3(new_n1169), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1168), .A2(new_n1170), .B1(new_n1081), .B2(new_n1078), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1070), .B(new_n1098), .C1(new_n1153), .C2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1006), .B1(G2090), .B2(new_n1101), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1025), .B1(G8), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1027), .A2(new_n1050), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1069), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n988), .A2(KEYINPUT110), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n972), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n987), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT112), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT112), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n987), .A2(new_n1183), .A3(new_n1180), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n992), .B1(new_n1176), .B2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n950), .A2(new_n952), .ZN(new_n1189));
  INV_X1    g763(.A(G401), .ZN(new_n1190));
  INV_X1    g764(.A(G229), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g766(.A1(new_n895), .A2(G319), .A3(new_n673), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g768(.A(G401), .B(G229), .C1(new_n950), .C2(new_n952), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n895), .A2(G319), .A3(new_n673), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n1195), .A2(KEYINPUT127), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1194), .A2(new_n1197), .ZN(G308));
  NAND2_X1  g772(.A1(new_n1195), .A2(new_n1196), .ZN(G225));
endmodule


