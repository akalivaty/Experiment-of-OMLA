//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  AND4_X1   g007(.A1(new_n187), .A2(new_n191), .A3(new_n193), .A4(KEYINPUT16), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n190), .A3(G125), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n195), .A2(KEYINPUT75), .A3(G146), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(new_n193), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT74), .B1(new_n199), .B2(new_n196), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n188), .A2(new_n187), .A3(KEYINPUT16), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n200), .A2(G146), .A3(new_n201), .A4(new_n197), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n200), .A2(new_n197), .A3(new_n201), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n198), .A2(new_n204), .A3(new_n207), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  XNOR2_X1  g023(.A(G119), .B(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n214), .B(new_n216), .C1(G119), .C2(new_n215), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G110), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n208), .A2(new_n211), .A3(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(KEYINPUT76), .B(G110), .Z(new_n220));
  OAI22_X1  g034(.A1(new_n217), .A2(new_n220), .B1(new_n210), .B2(new_n209), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n202), .B(new_n221), .C1(G146), .C2(new_n199), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT77), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n219), .A2(new_n225), .A3(new_n222), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT22), .B(G137), .Z(new_n227));
  INV_X1    g041(.A(G221), .ZN(new_n228));
  INV_X1    g042(.A(G234), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n228), .A2(new_n229), .A3(G953), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n227), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n219), .A2(new_n225), .A3(new_n222), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G902), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g052(.A(G217), .B1(new_n229), .B2(G902), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(KEYINPUT73), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n235), .A2(new_n241), .A3(new_n236), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n240), .A2(G902), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT32), .ZN(new_n247));
  INV_X1    g061(.A(G472), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n236), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n206), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n215), .A2(KEYINPUT0), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT0), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n261), .A3(KEYINPUT65), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n215), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n253), .A2(new_n262), .B1(new_n251), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n268), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(KEYINPUT66), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n276), .A3(G131), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT68), .B1(new_n275), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n264), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n282), .A2(new_n254), .A3(new_n256), .ZN(new_n283));
  AOI21_X1  g097(.A(G128), .B1(new_n254), .B2(new_n256), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n255), .A2(KEYINPUT1), .A3(G146), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n283), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n268), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n266), .A2(G137), .ZN(new_n289));
  OAI21_X1  g103(.A(G131), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n274), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n295), .B(new_n264), .C1(new_n278), .C2(new_n279), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n294), .A4(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT2), .B(G113), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(G116), .A2(G119), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(G116), .A2(G119), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n275), .A2(new_n277), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n264), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n291), .B(KEYINPUT67), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n287), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n297), .A2(new_n307), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G237), .A2(G953), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G210), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g135(.A(new_n307), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n281), .A2(new_n322), .A3(new_n294), .A4(new_n296), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n315), .A2(KEYINPUT31), .A3(new_n321), .A4(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n312), .A2(new_n307), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n308), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n292), .B1(new_n335), .B2(new_n264), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT28), .B1(new_n336), .B2(new_n322), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n321), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n249), .B1(new_n328), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n247), .B1(new_n341), .B2(KEYINPUT72), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n326), .A2(new_n327), .B1(new_n338), .B2(new_n339), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n343), .B(KEYINPUT32), .C1(new_n344), .C2(new_n249), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n338), .A2(new_n339), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n321), .B1(new_n315), .B2(new_n323), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(KEYINPUT29), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n281), .A2(new_n294), .A3(new_n296), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n307), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n352), .B2(new_n323), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n337), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT29), .A3(new_n321), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n236), .ZN(new_n356));
  OAI21_X1  g170(.A(G472), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n246), .B1(new_n346), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT9), .B(G234), .Z(new_n359));
  AOI21_X1  g173(.A(new_n228), .B1(new_n359), .B2(new_n236), .ZN(new_n360));
  INV_X1    g174(.A(G469), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n236), .ZN(new_n362));
  INV_X1    g176(.A(G104), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(new_n363), .B2(G107), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(G101), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(G101), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n364), .A2(new_n367), .A3(new_n318), .A4(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n264), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n376));
  XNOR2_X1  g190(.A(G104), .B(G107), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT78), .B1(new_n377), .B2(new_n318), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT78), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n363), .A2(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n366), .A2(G104), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n379), .B(G101), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n373), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n376), .B1(new_n383), .B2(new_n287), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n382), .A2(new_n373), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n282), .A2(new_n254), .A3(new_n256), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n285), .C1(G128), .C2(new_n251), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(KEYINPUT10), .A3(new_n387), .A4(new_n378), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n375), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n335), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n335), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n335), .B2(new_n389), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G110), .B(G140), .ZN(new_n396));
  INV_X1    g210(.A(G953), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G227), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n396), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT12), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n278), .A2(new_n279), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n383), .B(new_n387), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n383), .B(new_n287), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT12), .A3(new_n309), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n375), .A2(new_n384), .A3(new_n388), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n409), .B2(new_n403), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n362), .B1(new_n412), .B2(new_n361), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n410), .B1(new_n393), .B2(new_n394), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n390), .B1(new_n405), .B2(new_n407), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(G469), .C1(new_n415), .C2(new_n399), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n360), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n418));
  AOI21_X1  g232(.A(G143), .B1(new_n316), .B2(G214), .ZN(new_n419));
  OAI21_X1  g233(.A(G131), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n316), .A2(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n255), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n273), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n420), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT17), .A3(G131), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n429), .A2(new_n207), .A3(new_n198), .A4(new_n204), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n188), .B(G146), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n420), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n427), .A2(KEYINPUT83), .A3(KEYINPUT18), .A4(G131), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n422), .B(new_n423), .C1(new_n433), .C2(new_n273), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(G104), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n206), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n420), .A2(new_n424), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n202), .A3(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n449), .A2(new_n443), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n441), .A2(new_n444), .B1(new_n440), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT85), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT20), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n443), .B1(new_n430), .B2(new_n440), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n450), .A2(new_n440), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n458));
  NOR4_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n453), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n441), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n461), .B2(new_n441), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G475), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n359), .A2(G217), .A3(new_n397), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G116), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(G116), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n469), .A2(new_n470), .A3(G107), .ZN(new_n471));
  XNOR2_X1  g285(.A(G128), .B(G143), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(G134), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n468), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT87), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n470), .A2(new_n474), .ZN(new_n478));
  OAI211_X1 g292(.A(KEYINPUT87), .B(new_n468), .C1(new_n470), .C2(new_n474), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n471), .B(new_n473), .C1(G107), .C2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n366), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n472), .A2(new_n266), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n266), .B1(new_n472), .B2(KEYINPUT13), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n255), .A2(G128), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(KEYINPUT13), .B2(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n466), .B1(new_n481), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n471), .B1(new_n480), .B2(G107), .ZN(new_n490));
  INV_X1    g304(.A(new_n473), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(new_n466), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI211_X1 g309(.A(KEYINPUT88), .B(G902), .C1(new_n489), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G478), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n489), .A2(new_n495), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n236), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n498), .B1(new_n502), .B2(new_n496), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n397), .A2(G952), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(G237), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n236), .B(new_n397), .C1(G234), .C2(G237), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT21), .B(G898), .Z(new_n510));
  OAI21_X1  g324(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT89), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n465), .A2(new_n504), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G214), .B1(G237), .B2(G902), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(KEYINPUT5), .A2(G119), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n300), .A2(KEYINPUT5), .B1(G116), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n518), .A2(G113), .B1(new_n299), .B2(new_n300), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT80), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n378), .A4(new_n385), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n213), .A3(G116), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(G113), .C1(new_n305), .C2(new_n522), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n301), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT80), .B1(new_n525), .B2(new_n383), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n374), .A2(new_n307), .A3(new_n371), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(G110), .B(G122), .Z(new_n529));
  OR2_X1    g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n529), .B(KEYINPUT8), .Z(new_n531));
  AND2_X1   g345(.A1(new_n525), .A2(new_n383), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n525), .A2(new_n383), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n264), .A2(G125), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n387), .A2(new_n192), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n538));
  INV_X1    g352(.A(G224), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n538), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n535), .B2(new_n536), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n530), .B(new_n534), .C1(new_n541), .C2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n529), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT81), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT6), .B1(new_n528), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n528), .A2(new_n529), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n540), .B(KEYINPUT82), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n537), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n236), .B(new_n544), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G210), .B1(G237), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n528), .A2(new_n546), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT6), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n528), .A2(KEYINPUT6), .A3(new_n546), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n530), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(G902), .B1(new_n562), .B2(new_n552), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n555), .A3(new_n544), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n516), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n417), .A2(new_n514), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n358), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  INV_X1    g382(.A(new_n246), .ZN(new_n569));
  INV_X1    g383(.A(new_n341), .ZN(new_n570));
  OAI21_X1  g384(.A(G472), .B1(new_n344), .B2(G902), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n417), .A4(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n501), .A2(KEYINPUT33), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n501), .A2(KEYINPUT33), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(G478), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n497), .A2(new_n236), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n501), .A2(new_n497), .A3(new_n236), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n465), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n564), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT90), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n554), .A2(new_n582), .A3(new_n556), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n515), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n512), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n572), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT34), .B(G104), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G6));
  INV_X1    g403(.A(new_n465), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n572), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G107), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n592), .B(new_n595), .ZN(G9));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n219), .A2(new_n597), .A3(new_n222), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n219), .B2(new_n222), .ZN(new_n600));
  OAI22_X1  g414(.A1(new_n599), .A2(new_n600), .B1(KEYINPUT36), .B2(new_n233), .ZN(new_n601));
  INV_X1    g415(.A(new_n600), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n598), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n604), .A3(new_n244), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT94), .A4(new_n244), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n243), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n566), .A2(new_n570), .A3(new_n571), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT95), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(G12));
  NAND2_X1  g428(.A1(new_n346), .A2(new_n357), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n610), .A2(new_n417), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT96), .B(G900), .Z(new_n617));
  AOI21_X1  g431(.A(new_n506), .B1(new_n508), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n591), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n585), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  XNOR2_X1  g435(.A(new_n618), .B(KEYINPUT39), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n417), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT40), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n625), .A2(new_n516), .A3(new_n610), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n557), .A2(new_n564), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT38), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n460), .A2(new_n464), .B1(new_n499), .B2(new_n503), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n352), .A2(new_n339), .A3(new_n323), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n630), .A2(new_n236), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n315), .A2(new_n323), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n321), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n248), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n342), .B2(new_n345), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n626), .A2(new_n628), .A3(new_n629), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G143), .ZN(G45));
  NOR2_X1   g452(.A1(new_n580), .A2(new_n618), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n615), .A2(new_n585), .A3(new_n616), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G146), .ZN(G48));
  NOR2_X1   g455(.A1(new_n586), .A2(new_n580), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n412), .B(new_n361), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n360), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n615), .A2(new_n569), .A3(new_n642), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT97), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT41), .B(G113), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  NOR2_X1   g462(.A1(new_n586), .A2(new_n591), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n615), .A2(new_n569), .A3(new_n649), .A4(new_n644), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G116), .ZN(G18));
  AND3_X1   g465(.A1(new_n644), .A2(new_n585), .A3(new_n610), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n615), .A2(new_n514), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G119), .ZN(G21));
  NAND4_X1  g468(.A1(new_n581), .A2(new_n629), .A3(new_n515), .A4(new_n583), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n339), .B1(new_n353), .B2(new_n337), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n249), .B1(new_n328), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n328), .B2(new_n340), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n248), .ZN(new_n663));
  OAI211_X1 g477(.A(KEYINPUT98), .B(G472), .C1(new_n344), .C2(G902), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n643), .A2(new_n513), .A3(new_n360), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(new_n665), .A3(new_n569), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n652), .A3(new_n639), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G125), .ZN(G27));
  OAI21_X1  g484(.A(KEYINPUT79), .B1(new_n409), .B2(new_n403), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n335), .A2(new_n389), .A3(new_n392), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n399), .B1(new_n673), .B2(new_n391), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n408), .A2(new_n410), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n361), .B(new_n236), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n416), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n362), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT12), .B1(new_n335), .B2(new_n406), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n404), .A2(new_n402), .A3(new_n308), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n400), .B1(new_n682), .B2(new_n390), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT100), .A3(G469), .A4(new_n414), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n676), .A2(new_n678), .A3(new_n679), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n688));
  INV_X1    g502(.A(new_n360), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n627), .A2(new_n516), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n413), .A2(new_n686), .A3(new_n678), .A4(new_n684), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n685), .A2(KEYINPUT101), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n689), .A4(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n358), .A2(new_n696), .A3(new_n639), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n570), .A2(new_n247), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n341), .A2(KEYINPUT32), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n357), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n569), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(KEYINPUT42), .A3(new_n696), .A4(new_n639), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  NAND3_X1  g520(.A1(new_n358), .A2(new_n696), .A3(new_n619), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G134), .ZN(G36));
  NAND2_X1  g522(.A1(new_n590), .A2(new_n579), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT43), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n571), .A2(new_n570), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n610), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n713), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(KEYINPUT105), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n683), .A2(new_n414), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(KEYINPUT45), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(G469), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n679), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT103), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n722), .A2(new_n727), .A3(KEYINPUT46), .A4(new_n679), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n726), .A3(new_n676), .A4(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n689), .A3(new_n623), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n690), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n717), .B2(KEYINPUT105), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n715), .A2(new_n718), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G137), .ZN(G39));
  NAND2_X1  g549(.A1(new_n729), .A2(new_n689), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT47), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n615), .A2(new_n569), .A3(new_n732), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n639), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G140), .ZN(G42));
  XOR2_X1   g555(.A(new_n505), .B(KEYINPUT115), .Z(new_n742));
  AND3_X1   g556(.A1(new_n665), .A2(new_n569), .A3(new_n506), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n644), .A3(new_n710), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n628), .A2(new_n515), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n744), .A2(new_n748), .A3(new_n515), .A4(new_n628), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n732), .A2(new_n643), .A3(new_n507), .A4(new_n360), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n710), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT113), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n607), .A2(new_n608), .ZN(new_n754));
  AOI21_X1  g568(.A(G902), .B1(new_n232), .B2(new_n234), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT25), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n756), .B2(new_n240), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n757), .B(new_n660), .C1(new_n663), .C2(new_n664), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n635), .A2(new_n569), .A3(new_n751), .ZN(new_n760));
  INV_X1    g574(.A(new_n579), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n590), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n750), .A2(KEYINPUT114), .A3(new_n759), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n643), .B(KEYINPUT112), .Z(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n737), .B1(new_n689), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n690), .A3(new_n710), .A4(new_n743), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n759), .B(new_n762), .C1(new_n747), .C2(new_n749), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n774));
  INV_X1    g588(.A(new_n767), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n768), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n753), .A2(new_n703), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT48), .ZN(new_n778));
  INV_X1    g592(.A(new_n580), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n745), .A2(new_n585), .B1(new_n779), .B2(new_n760), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n742), .A2(new_n771), .A3(new_n776), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT107), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n696), .A2(new_n758), .A3(new_n639), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n732), .A2(new_n504), .A3(new_n465), .A4(new_n618), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n615), .A2(new_n616), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n707), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n705), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n591), .A2(new_n580), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n512), .A3(new_n565), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n572), .A2(new_n790), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n567), .A2(new_n653), .A3(new_n791), .A4(new_n611), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n645), .A2(new_n650), .A3(new_n667), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n783), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n610), .B2(new_n618), .ZN(new_n798));
  INV_X1    g612(.A(new_n618), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n243), .A2(new_n609), .A3(KEYINPUT108), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n798), .A2(new_n689), .A3(new_n687), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT99), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n655), .B(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT109), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n801), .A2(new_n635), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n634), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n346), .A2(new_n806), .B1(new_n656), .B2(new_n657), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n687), .A2(new_n689), .A3(new_n800), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT108), .B1(new_n757), .B2(new_n799), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT109), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n620), .A2(new_n640), .A3(new_n669), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n796), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n807), .A2(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n804), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n807), .A2(new_n810), .A3(KEYINPUT109), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n620), .A2(new_n640), .A3(new_n669), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n567), .A2(new_n653), .A3(new_n791), .A4(new_n611), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n645), .A2(new_n650), .A3(new_n667), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(KEYINPUT107), .A3(new_n705), .A4(new_n787), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n795), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n705), .A2(new_n787), .A3(new_n792), .A4(new_n793), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n795), .A2(KEYINPUT53), .A3(new_n821), .A4(new_n825), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n828), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n821), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n827), .B2(new_n826), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(KEYINPUT110), .A3(new_n829), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n782), .A2(new_n834), .A3(new_n837), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT116), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n840), .A2(new_n834), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n837), .A4(new_n782), .ZN(new_n845));
  NOR2_X1   g659(.A1(G952), .A2(G953), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT117), .Z(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n246), .A2(new_n709), .A3(new_n360), .A4(new_n516), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT106), .Z(new_n850));
  XNOR2_X1  g664(.A(new_n643), .B(KEYINPUT49), .ZN(new_n851));
  OR4_X1    g665(.A1(new_n628), .A2(new_n850), .A3(new_n636), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(G75));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n839), .B2(new_n236), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n828), .A2(new_n831), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT118), .A3(G902), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n556), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n562), .B(new_n553), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT55), .Z(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n397), .A2(G952), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(G210), .A3(G902), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n867), .B2(new_n860), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n863), .A2(KEYINPUT120), .A3(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(G51));
  NAND2_X1  g687(.A1(new_n855), .A2(new_n857), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n874), .A2(new_n722), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(new_n832), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n362), .B(KEYINPUT57), .Z(new_n878));
  OAI22_X1  g692(.A1(new_n877), .A2(new_n878), .B1(new_n674), .B2(new_n675), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n864), .B1(new_n875), .B2(new_n879), .ZN(G54));
  NAND2_X1  g694(.A1(KEYINPUT58), .A2(G475), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n882), .A2(new_n451), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n451), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n864), .ZN(G60));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n876), .A2(new_n832), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n573), .A2(new_n574), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n577), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n864), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n840), .A2(new_n834), .A3(new_n837), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n894), .A2(new_n890), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n886), .B(new_n893), .C1(new_n895), .C2(new_n888), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n888), .B1(new_n894), .B2(new_n890), .ZN(new_n897));
  INV_X1    g711(.A(new_n864), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n877), .B2(new_n891), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(G63));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n828), .B2(new_n831), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n905), .B2(new_n235), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n601), .A2(new_n604), .ZN(new_n907));
  INV_X1    g721(.A(new_n904), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n856), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(KEYINPUT124), .A3(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n906), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n856), .A2(new_n907), .A3(new_n908), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n916), .B(new_n898), .C1(new_n235), .C2(new_n905), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n913), .B1(new_n917), .B2(new_n902), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(G66));
  INV_X1    g734(.A(new_n510), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n921), .B2(new_n539), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n824), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n550), .B1(G898), .B2(new_n397), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G69));
  NAND2_X1  g739(.A1(new_n297), .A2(new_n314), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT126), .B(KEYINPUT127), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n445), .A2(new_n446), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT125), .Z(new_n930));
  XOR2_X1   g744(.A(new_n928), .B(new_n930), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n740), .A2(new_n734), .A3(new_n819), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n731), .A2(new_n658), .A3(new_n703), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n705), .A3(new_n707), .A4(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n935), .B2(new_n397), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n397), .A2(G900), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n819), .A2(new_n637), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n624), .A2(new_n732), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n358), .A2(new_n789), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n734), .A3(new_n740), .A4(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n931), .A2(G953), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n936), .A2(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n397), .B1(G227), .B2(G900), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G72));
  NAND2_X1  g760(.A1(G472), .A2(G902), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT63), .Z(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n942), .B2(new_n794), .ZN(new_n949));
  INV_X1    g763(.A(new_n633), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n864), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n935), .B2(new_n794), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n632), .A2(new_n321), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n948), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n950), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n836), .B2(new_n957), .ZN(G57));
endmodule


