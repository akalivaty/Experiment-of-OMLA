

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  XNOR2_X1 U322 ( .A(n469), .B(KEYINPUT48), .ZN(n470) );
  XNOR2_X1 U323 ( .A(n426), .B(n378), .ZN(n519) );
  XOR2_X1 U324 ( .A(n379), .B(KEYINPUT27), .Z(n290) );
  XOR2_X1 U325 ( .A(G64GAT), .B(KEYINPUT72), .Z(n291) );
  INV_X1 U326 ( .A(KEYINPUT94), .ZN(n371) );
  XNOR2_X1 U327 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U328 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U329 ( .A(n442), .B(n373), .ZN(n374) );
  XNOR2_X1 U330 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n476) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U333 ( .A(n471), .B(n470), .ZN(n546) );
  NOR2_X1 U334 ( .A1(n516), .A2(n486), .ZN(n451) );
  INV_X1 U335 ( .A(G43GAT), .ZN(n452) );
  XNOR2_X1 U336 ( .A(n451), .B(KEYINPUT38), .ZN(n502) );
  XNOR2_X1 U337 ( .A(n479), .B(KEYINPUT58), .ZN(n480) );
  XNOR2_X1 U338 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U339 ( .A(n481), .B(n480), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n293) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(n294), .B(KEYINPUT87), .Z(n296) );
  XOR2_X1 U345 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XNOR2_X1 U346 ( .A(G15GAT), .B(n447), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U348 ( .A(KEYINPUT86), .B(G176GAT), .Z(n298) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U351 ( .A(n300), .B(n299), .Z(n306) );
  XNOR2_X1 U352 ( .A(G127GAT), .B(KEYINPUT85), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(KEYINPUT84), .ZN(n302) );
  XOR2_X1 U354 ( .A(n302), .B(KEYINPUT0), .Z(n304) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n343) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(n343), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(G190GAT), .Z(n308) );
  XNOR2_X1 U360 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U362 ( .A(KEYINPUT17), .B(n309), .Z(n375) );
  XOR2_X2 U363 ( .A(n310), .B(n375), .Z(n531) );
  XOR2_X1 U364 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n412) );
  XOR2_X1 U365 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n312) );
  XNOR2_X1 U366 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n311) );
  XNOR2_X1 U367 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U368 ( .A(n313), .B(KEYINPUT11), .Z(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT75), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U370 ( .A(G218GAT), .B(n353), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n321) );
  XNOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .ZN(n446) );
  XOR2_X1 U373 ( .A(G29GAT), .B(G43GAT), .Z(n317) );
  XNOR2_X1 U374 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U375 ( .A(n317), .B(n316), .ZN(n414) );
  XNOR2_X1 U376 ( .A(n446), .B(n414), .ZN(n319) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U379 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U380 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n323) );
  XNOR2_X1 U381 ( .A(G190GAT), .B(G92GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U383 ( .A(G106GAT), .B(G134GAT), .Z(n325) );
  XNOR2_X1 U384 ( .A(G50GAT), .B(G36GAT), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n555) );
  INV_X1 U388 ( .A(n555), .ZN(n539) );
  XNOR2_X1 U389 ( .A(KEYINPUT36), .B(n539), .ZN(n585) );
  XOR2_X1 U390 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n331) );
  XNOR2_X1 U391 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n347) );
  XOR2_X1 U393 ( .A(G85GAT), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U394 ( .A(G29GAT), .B(G120GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U396 ( .A(G57GAT), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U397 ( .A(G141GAT), .B(G1GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U399 ( .A(n337), .B(n336), .Z(n345) );
  XOR2_X1 U400 ( .A(G155GAT), .B(KEYINPUT3), .Z(n339) );
  XNOR2_X1 U401 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n361) );
  XOR2_X1 U403 ( .A(n361), .B(KEYINPUT4), .Z(n341) );
  NAND2_X1 U404 ( .A1(G225GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n543) );
  XNOR2_X1 U409 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n367) );
  XNOR2_X1 U410 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n348), .B(KEYINPUT89), .ZN(n349) );
  XOR2_X1 U412 ( .A(n349), .B(KEYINPUT90), .Z(n351) );
  XNOR2_X1 U413 ( .A(G204GAT), .B(G218GAT), .ZN(n350) );
  XOR2_X1 U414 ( .A(n351), .B(n350), .Z(n376) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n352), .B(G148GAT), .ZN(n434) );
  XOR2_X1 U417 ( .A(n434), .B(KEYINPUT22), .Z(n355) );
  XNOR2_X1 U418 ( .A(G197GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U420 ( .A(n376), .B(n356), .Z(n365) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n358) );
  NAND2_X1 U422 ( .A1(G228GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(n359), .B(KEYINPUT92), .Z(n363) );
  XNOR2_X1 U425 ( .A(G50GAT), .B(G22GAT), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n360), .B(G141GAT), .ZN(n427) );
  XNOR2_X1 U427 ( .A(n427), .B(n361), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n475) );
  NOR2_X1 U430 ( .A1(n531), .A2(n475), .ZN(n366) );
  XOR2_X1 U431 ( .A(n367), .B(n366), .Z(n569) );
  XOR2_X1 U432 ( .A(G8GAT), .B(G197GAT), .Z(n369) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(G36GAT), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n426) );
  XNOR2_X1 U435 ( .A(G176GAT), .B(G92GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n291), .B(n370), .ZN(n442) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n519), .B(KEYINPUT95), .ZN(n379) );
  AND2_X1 U441 ( .A1(n569), .A2(n290), .ZN(n544) );
  NAND2_X1 U442 ( .A1(n531), .A2(n519), .ZN(n380) );
  NAND2_X1 U443 ( .A1(n475), .A2(n380), .ZN(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT25), .B(n381), .ZN(n382) );
  NOR2_X1 U445 ( .A1(n544), .A2(n382), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n383), .B(KEYINPUT98), .ZN(n384) );
  NOR2_X1 U447 ( .A1(n543), .A2(n384), .ZN(n389) );
  INV_X1 U448 ( .A(n543), .ZN(n385) );
  XOR2_X1 U449 ( .A(n475), .B(KEYINPUT28), .Z(n524) );
  NOR2_X1 U450 ( .A1(n385), .A2(n524), .ZN(n386) );
  NAND2_X1 U451 ( .A1(n386), .A2(n290), .ZN(n529) );
  NOR2_X1 U452 ( .A1(n531), .A2(n529), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n387), .B(KEYINPUT96), .ZN(n388) );
  NOR2_X1 U454 ( .A1(n389), .A2(n388), .ZN(n483) );
  NOR2_X1 U455 ( .A1(n585), .A2(n483), .ZN(n410) );
  XOR2_X1 U456 ( .A(G155GAT), .B(G211GAT), .Z(n391) );
  XNOR2_X1 U457 ( .A(G22GAT), .B(G127GAT), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U459 ( .A(KEYINPUT83), .B(G64GAT), .Z(n393) );
  XNOR2_X1 U460 ( .A(G8GAT), .B(G78GAT), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U462 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U463 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n397) );
  NAND2_X1 U464 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U466 ( .A(KEYINPUT12), .B(n398), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n400), .B(n399), .ZN(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n402) );
  XNOR2_X1 U469 ( .A(KEYINPUT82), .B(KEYINPUT79), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n407) );
  XNOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n403), .B(KEYINPUT71), .ZN(n443) );
  XOR2_X1 U473 ( .A(n443), .B(G71GAT), .Z(n405) );
  XOR2_X1 U474 ( .A(G15GAT), .B(G1GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(n419), .B(G183GAT), .ZN(n404) );
  XNOR2_X1 U476 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U477 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n567) );
  NAND2_X1 U479 ( .A1(n410), .A2(n567), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U481 ( .A(KEYINPUT102), .B(n413), .Z(n516) );
  XOR2_X1 U482 ( .A(n414), .B(KEYINPUT67), .Z(n416) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n418) );
  INV_X1 U485 ( .A(KEYINPUT68), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n421) );
  XNOR2_X1 U487 ( .A(G113GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U489 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n423) );
  XNOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n422) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n571) );
  XOR2_X1 U495 ( .A(n571), .B(KEYINPUT70), .Z(n558) );
  XOR2_X1 U496 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n431) );
  XNOR2_X1 U497 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n434), .B(KEYINPUT31), .ZN(n432) );
  AND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  NAND2_X1 U501 ( .A1(n432), .A2(n435), .ZN(n439) );
  INV_X1 U502 ( .A(KEYINPUT31), .ZN(n433) );
  XNOR2_X1 U503 ( .A(n434), .B(n433), .ZN(n437) );
  INV_X1 U504 ( .A(n435), .ZN(n436) );
  NAND2_X1 U505 ( .A1(n437), .A2(n436), .ZN(n438) );
  NAND2_X1 U506 ( .A1(n439), .A2(n438), .ZN(n440) );
  XOR2_X1 U507 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n445), .B(n444), .ZN(n449) );
  INV_X1 U510 ( .A(n456), .ZN(n576) );
  NOR2_X1 U511 ( .A1(n558), .A2(n576), .ZN(n450) );
  XOR2_X1 U512 ( .A(KEYINPUT74), .B(n450), .Z(n486) );
  NAND2_X1 U513 ( .A1(n531), .A2(n502), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(n549) );
  NAND2_X1 U517 ( .A1(n549), .A2(n571), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT114), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n460), .A2(n567), .ZN(n461) );
  NOR2_X1 U521 ( .A1(n555), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT47), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n585), .A2(n567), .ZN(n463) );
  XNOR2_X1 U524 ( .A(KEYINPUT45), .B(n463), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n464), .A2(n456), .ZN(n465) );
  XNOR2_X1 U526 ( .A(KEYINPUT115), .B(n465), .ZN(n466) );
  NAND2_X1 U527 ( .A1(n466), .A2(n558), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n468), .A2(n467), .ZN(n471) );
  INV_X1 U529 ( .A(KEYINPUT116), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n519), .B(KEYINPUT121), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n546), .A2(n472), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT54), .B(n473), .Z(n474) );
  NOR2_X1 U533 ( .A1(n543), .A2(n474), .ZN(n570) );
  NAND2_X1 U534 ( .A1(n570), .A2(n475), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n478), .A2(n531), .ZN(n566) );
  NOR2_X1 U536 ( .A1(n539), .A2(n566), .ZN(n481) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n489) );
  NOR2_X1 U539 ( .A1(n555), .A2(n567), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT16), .ZN(n485) );
  INV_X1 U541 ( .A(n483), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n485), .A2(n484), .ZN(n505) );
  NOR2_X1 U543 ( .A1(n486), .A2(n505), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(n487), .Z(n494) );
  NAND2_X1 U545 ( .A1(n494), .A2(n543), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U547 ( .A(G1GAT), .B(n490), .Z(G1324GAT) );
  NAND2_X1 U548 ( .A1(n494), .A2(n519), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .Z(n493) );
  NAND2_X1 U551 ( .A1(n494), .A2(n531), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  XOR2_X1 U553 ( .A(G22GAT), .B(KEYINPUT101), .Z(n496) );
  NAND2_X1 U554 ( .A1(n494), .A2(n524), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  NAND2_X1 U557 ( .A1(n502), .A2(n543), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n500) );
  NAND2_X1 U560 ( .A1(n519), .A2(n502), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U564 ( .A1(n524), .A2(n502), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n507) );
  INV_X1 U567 ( .A(n549), .ZN(n562) );
  OR2_X1 U568 ( .A1(n571), .A2(n562), .ZN(n515) );
  NOR2_X1 U569 ( .A1(n505), .A2(n515), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n543), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U573 ( .A1(n512), .A2(n519), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT109), .Z(n511) );
  NAND2_X1 U576 ( .A1(n512), .A2(n531), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n524), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n518) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n543), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  XOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U586 ( .A1(n525), .A2(n519), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n531), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n546), .A2(n529), .ZN(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U597 ( .A1(n558), .A2(n538), .ZN(n532) );
  XOR2_X1 U598 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U599 ( .A1(n562), .A2(n538), .ZN(n534) );
  XNOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n535), .Z(G1341GAT) );
  NOR2_X1 U603 ( .A1(n567), .A2(n538), .ZN(n536) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(n536), .Z(n537) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n541) );
  XNOR2_X1 U607 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT119), .Z(n548) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n556), .A2(n571), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U617 ( .A1(n556), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  INV_X1 U620 ( .A(n567), .ZN(n580) );
  NAND2_X1 U621 ( .A1(n556), .A2(n580), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n566), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n566), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n573) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n584) );
  INV_X1 U637 ( .A(n584), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n575) );
  XOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .Z(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U643 ( .A1(n581), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

