

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n634), .A2(G651), .ZN(n650) );
  BUF_X1 U550 ( .A(n682), .Z(n610) );
  AND2_X2 U551 ( .A1(n536), .A2(G2104), .ZN(n680) );
  NAND2_X1 U552 ( .A1(n751), .A2(n514), .ZN(n762) );
  INV_X1 U553 ( .A(G2105), .ZN(n536) );
  XOR2_X1 U554 ( .A(n691), .B(KEYINPUT27), .Z(n693) );
  AND2_X1 U555 ( .A1(n755), .A2(n516), .ZN(n756) );
  NOR2_X1 U556 ( .A1(n536), .A2(G2104), .ZN(n537) );
  AND2_X1 U557 ( .A1(n774), .A2(n773), .ZN(n776) );
  NOR2_X2 U558 ( .A1(n634), .A2(n524), .ZN(n586) );
  OR2_X1 U559 ( .A1(n750), .A2(n749), .ZN(n514) );
  AND2_X1 U560 ( .A1(n768), .A2(n771), .ZN(n515) );
  NOR2_X1 U561 ( .A1(n771), .A2(n754), .ZN(n516) );
  NOR2_X1 U562 ( .A1(n792), .A2(n791), .ZN(n517) );
  NOR2_X2 U563 ( .A1(n688), .A2(n687), .ZN(G160) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n518) );
  INV_X1 U565 ( .A(KEYINPUT92), .ZN(n696) );
  XNOR2_X1 U566 ( .A(n697), .B(n696), .ZN(n711) );
  INV_X1 U567 ( .A(KEYINPUT95), .ZN(n735) );
  XNOR2_X1 U568 ( .A(n736), .B(n735), .ZN(n742) );
  INV_X1 U569 ( .A(n957), .ZN(n754) );
  XNOR2_X1 U570 ( .A(n744), .B(KEYINPUT32), .ZN(n751) );
  NOR2_X1 U571 ( .A1(n766), .A2(n765), .ZN(n767) );
  INV_X1 U572 ( .A(KEYINPUT98), .ZN(n775) );
  INV_X1 U573 ( .A(KEYINPUT71), .ZN(n591) );
  AND2_X1 U574 ( .A1(n517), .A2(n815), .ZN(n812) );
  XNOR2_X1 U575 ( .A(n591), .B(KEYINPUT15), .ZN(n592) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n519), .Z(n644) );
  INV_X1 U577 ( .A(G651), .ZN(n524) );
  NOR2_X1 U578 ( .A1(G543), .A2(n524), .ZN(n519) );
  NAND2_X1 U579 ( .A1(G63), .A2(n644), .ZN(n521) );
  XNOR2_X1 U580 ( .A(KEYINPUT68), .B(n518), .ZN(n634) );
  NAND2_X1 U581 ( .A1(G51), .A2(n650), .ZN(n520) );
  NAND2_X1 U582 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n522), .ZN(n530) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n645) );
  NAND2_X1 U585 ( .A1(n645), .A2(G89), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(KEYINPUT4), .ZN(n526) );
  NAND2_X1 U587 ( .A1(G76), .A2(n586), .ZN(n525) );
  NAND2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U589 ( .A(KEYINPUT72), .B(n527), .Z(n528) );
  XNOR2_X1 U590 ( .A(KEYINPUT5), .B(n528), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT7), .B(n531), .Z(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n533) );
  NOR2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(n682) );
  NAND2_X1 U597 ( .A1(G138), .A2(n682), .ZN(n535) );
  NAND2_X1 U598 ( .A1(G102), .A2(n680), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n541) );
  AND2_X1 U600 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U601 ( .A1(n886), .A2(G114), .ZN(n539) );
  XNOR2_X2 U602 ( .A(n537), .B(KEYINPUT66), .ZN(n888) );
  NAND2_X1 U603 ( .A1(G126), .A2(n888), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(G164) );
  XOR2_X1 U606 ( .A(G2430), .B(G2443), .Z(n543) );
  XNOR2_X1 U607 ( .A(KEYINPUT101), .B(G2451), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n550) );
  XOR2_X1 U609 ( .A(G2435), .B(G2427), .Z(n545) );
  XNOR2_X1 U610 ( .A(G2446), .B(G2454), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(n546), .B(G2438), .Z(n548) );
  XNOR2_X1 U613 ( .A(G1341), .B(G1348), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U616 ( .A1(n551), .A2(G14), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  INV_X1 U619 ( .A(G82), .ZN(G220) );
  NAND2_X1 U620 ( .A1(G88), .A2(n645), .ZN(n553) );
  NAND2_X1 U621 ( .A1(G75), .A2(n586), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U623 ( .A1(G62), .A2(n644), .ZN(n555) );
  NAND2_X1 U624 ( .A1(G50), .A2(n650), .ZN(n554) );
  NAND2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U626 ( .A1(n557), .A2(n556), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G78), .A2(n586), .ZN(n559) );
  NAND2_X1 U628 ( .A1(G53), .A2(n650), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G65), .A2(n644), .ZN(n561) );
  NAND2_X1 U631 ( .A1(G91), .A2(n645), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n564), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n831) );
  NAND2_X1 U638 ( .A1(n831), .A2(G567), .ZN(n566) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n644), .ZN(n567) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n567), .Z(n573) );
  NAND2_X1 U642 ( .A1(n645), .A2(G81), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U644 ( .A1(G68), .A2(n586), .ZN(n569) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U647 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n650), .A2(G43), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n938) );
  INV_X1 U650 ( .A(n938), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n576), .A2(G860), .ZN(G153) );
  NAND2_X1 U652 ( .A1(G64), .A2(n644), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G52), .A2(n650), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G90), .A2(n645), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G77), .A2(n586), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U658 ( .A(KEYINPUT9), .B(n581), .Z(n582) );
  NOR2_X1 U659 ( .A1(n583), .A2(n582), .ZN(G171) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G66), .A2(n644), .ZN(n585) );
  NAND2_X1 U663 ( .A1(G92), .A2(n645), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U665 ( .A1(G79), .A2(n586), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n650), .A2(G54), .ZN(n587) );
  NAND2_X1 U667 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n593) );
  XNOR2_X2 U669 ( .A(n593), .B(n592), .ZN(n941) );
  INV_X1 U670 ( .A(G868), .ZN(n660) );
  NAND2_X1 U671 ( .A1(n941), .A2(n660), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(G284) );
  XNOR2_X1 U673 ( .A(KEYINPUT73), .B(G868), .ZN(n596) );
  NOR2_X1 U674 ( .A1(G286), .A2(n596), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT74), .ZN(n599) );
  NOR2_X1 U676 ( .A1(G299), .A2(G868), .ZN(n598) );
  NOR2_X1 U677 ( .A1(n599), .A2(n598), .ZN(G297) );
  INV_X1 U678 ( .A(G559), .ZN(n600) );
  NOR2_X1 U679 ( .A1(G860), .A2(n600), .ZN(n601) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(n601), .ZN(n602) );
  INV_X1 U681 ( .A(n941), .ZN(n620) );
  NAND2_X1 U682 ( .A1(n602), .A2(n620), .ZN(n603) );
  XNOR2_X1 U683 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n938), .ZN(n604) );
  XNOR2_X1 U685 ( .A(KEYINPUT76), .B(n604), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G868), .A2(n620), .ZN(n605) );
  NOR2_X1 U687 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U689 ( .A1(n888), .A2(G123), .ZN(n608) );
  XOR2_X1 U690 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  XNOR2_X1 U691 ( .A(n609), .B(KEYINPUT77), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G135), .A2(n610), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U694 ( .A(KEYINPUT78), .B(n613), .ZN(n617) );
  NAND2_X1 U695 ( .A1(G99), .A2(n680), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G111), .A2(n886), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n978) );
  XNOR2_X1 U699 ( .A(G2096), .B(n978), .ZN(n619) );
  INV_X1 U700 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U702 ( .A1(G559), .A2(n620), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n938), .B(n621), .ZN(n658) );
  NOR2_X1 U704 ( .A1(n658), .A2(G860), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G67), .A2(n644), .ZN(n623) );
  NAND2_X1 U706 ( .A1(G93), .A2(n645), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G80), .A2(n586), .ZN(n624) );
  XNOR2_X1 U709 ( .A(KEYINPUT79), .B(n624), .ZN(n625) );
  NOR2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n650), .A2(G55), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n661) );
  XOR2_X1 U713 ( .A(n661), .B(KEYINPUT80), .Z(n629) );
  XNOR2_X1 U714 ( .A(n630), .B(n629), .ZN(G145) );
  NAND2_X1 U715 ( .A1(G49), .A2(n650), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n644), .A2(n633), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G61), .A2(n644), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G86), .A2(n645), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n586), .A2(G73), .ZN(n639) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n650), .A2(G48), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(G305) );
  AND2_X1 U729 ( .A1(n644), .A2(G60), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G85), .A2(n645), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G72), .A2(n586), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n650), .A2(G47), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(G290) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(G288), .ZN(n657) );
  XOR2_X1 U737 ( .A(G299), .B(G305), .Z(n653) );
  XNOR2_X1 U738 ( .A(n661), .B(n653), .ZN(n654) );
  XNOR2_X1 U739 ( .A(G166), .B(n654), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U741 ( .A(n657), .B(n656), .ZN(n841) );
  XOR2_X1 U742 ( .A(n658), .B(n841), .Z(n659) );
  NOR2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n663) );
  NOR2_X1 U744 ( .A1(G868), .A2(n661), .ZN(n662) );
  NOR2_X1 U745 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT81), .B(n664), .Z(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n666) );
  XOR2_X1 U748 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n665) );
  XNOR2_X1 U749 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U754 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U755 ( .A1(G219), .A2(G220), .ZN(n670) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U757 ( .A1(G218), .A2(n671), .ZN(n672) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(n672), .Z(n673) );
  NAND2_X1 U759 ( .A1(G96), .A2(n673), .ZN(n838) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n838), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U762 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U763 ( .A1(G108), .A2(n675), .ZN(n837) );
  NAND2_X1 U764 ( .A1(G567), .A2(n837), .ZN(n676) );
  NAND2_X1 U765 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U766 ( .A(KEYINPUT84), .B(n678), .ZN(n864) );
  NAND2_X1 U767 ( .A1(G661), .A2(G483), .ZN(n679) );
  NOR2_X1 U768 ( .A1(n864), .A2(n679), .ZN(n836) );
  NAND2_X1 U769 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NAND2_X1 U771 ( .A1(G101), .A2(n680), .ZN(n681) );
  XOR2_X1 U772 ( .A(KEYINPUT23), .B(n681), .Z(n684) );
  NAND2_X1 U773 ( .A1(n682), .A2(G137), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n684), .A2(n683), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n886), .A2(G113), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n888), .A2(G125), .ZN(n685) );
  NAND2_X1 U777 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G40), .A2(G160), .ZN(n777) );
  XNOR2_X1 U779 ( .A(n777), .B(KEYINPUT85), .ZN(n689) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n779) );
  NAND2_X2 U781 ( .A1(n689), .A2(n779), .ZN(n737) );
  INV_X1 U782 ( .A(n737), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n690), .A2(G2072), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G1956), .A2(n737), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U786 ( .A1(G299), .A2(n695), .ZN(n694) );
  XOR2_X1 U787 ( .A(KEYINPUT28), .B(n694), .Z(n718) );
  NOR2_X1 U788 ( .A1(G299), .A2(n695), .ZN(n697) );
  INV_X1 U789 ( .A(G1341), .ZN(n999) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n941), .ZN(n944) );
  NAND2_X1 U791 ( .A1(n999), .A2(n944), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n737), .A2(n698), .ZN(n701) );
  INV_X1 U793 ( .A(n737), .ZN(n720) );
  NAND2_X1 U794 ( .A1(n720), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U795 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n699), .A2(n703), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n938), .A2(n702), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n941), .A2(G2067), .ZN(n706) );
  INV_X1 U800 ( .A(n703), .ZN(n704) );
  NAND2_X1 U801 ( .A1(G1996), .A2(n704), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n707), .A2(n720), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G1348), .A2(n737), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G2067), .A2(n720), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n941), .A2(n714), .ZN(n715) );
  NOR2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U812 ( .A(n719), .B(KEYINPUT29), .ZN(n724) );
  XOR2_X1 U813 ( .A(G2078), .B(KEYINPUT25), .Z(n919) );
  NOR2_X1 U814 ( .A1(n919), .A2(n737), .ZN(n722) );
  XOR2_X1 U815 ( .A(KEYINPUT91), .B(G1961), .Z(n1010) );
  NOR2_X1 U816 ( .A1(n720), .A2(n1010), .ZN(n721) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n729) );
  OR2_X1 U818 ( .A1(G301), .A2(n729), .ZN(n723) );
  NAND2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n734) );
  NAND2_X1 U820 ( .A1(G8), .A2(n737), .ZN(n771) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n771), .ZN(n750) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n737), .ZN(n746) );
  NOR2_X1 U823 ( .A1(n750), .A2(n746), .ZN(n725) );
  NAND2_X1 U824 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U826 ( .A1(G168), .A2(n727), .ZN(n728) );
  XNOR2_X1 U827 ( .A(n728), .B(KEYINPUT93), .ZN(n731) );
  NAND2_X1 U828 ( .A1(n729), .A2(G301), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U830 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n745), .A2(G286), .ZN(n736) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n771), .ZN(n739) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n737), .ZN(n738) );
  NOR2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U836 ( .A1(G303), .A2(n740), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U839 ( .A(n745), .B(KEYINPUT94), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n746), .A2(G8), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n960) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n960), .A2(n752), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n762), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n957) );
  XNOR2_X1 U847 ( .A(n756), .B(KEYINPUT64), .ZN(n757) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n757), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n960), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U850 ( .A1(n758), .A2(n771), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n952) );
  NAND2_X1 U853 ( .A1(n761), .A2(n952), .ZN(n774) );
  INV_X1 U854 ( .A(n762), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G8), .A2(G166), .ZN(n763) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n763), .ZN(n764) );
  XNOR2_X1 U857 ( .A(n764), .B(KEYINPUT96), .ZN(n765) );
  XNOR2_X1 U858 ( .A(n767), .B(KEYINPUT97), .ZN(n768) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n769) );
  XOR2_X1 U860 ( .A(n769), .B(KEYINPUT24), .Z(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U862 ( .A1(n515), .A2(n772), .ZN(n773) );
  XNOR2_X1 U863 ( .A(n776), .B(n775), .ZN(n813) );
  XNOR2_X1 U864 ( .A(G1986), .B(G290), .ZN(n943) );
  XOR2_X1 U865 ( .A(KEYINPUT85), .B(n777), .Z(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n826) );
  AND2_X1 U867 ( .A1(n943), .A2(n826), .ZN(n792) );
  NAND2_X1 U868 ( .A1(G140), .A2(n610), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G104), .A2(n680), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n782), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n886), .A2(G116), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT86), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G128), .A2(n888), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U876 ( .A(n786), .B(KEYINPUT35), .Z(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U878 ( .A(KEYINPUT36), .B(n789), .Z(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT87), .B(n790), .ZN(n904) );
  XNOR2_X1 U880 ( .A(KEYINPUT37), .B(G2067), .ZN(n824) );
  NOR2_X1 U881 ( .A1(n904), .A2(n824), .ZN(n971) );
  NAND2_X1 U882 ( .A1(n826), .A2(n971), .ZN(n822) );
  INV_X1 U883 ( .A(n822), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G141), .A2(n610), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G129), .A2(n888), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G105), .A2(n680), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT89), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT38), .ZN(n797) );
  NOR2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n886), .A2(G117), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n874) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n874), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT90), .B(n801), .Z(n810) );
  NAND2_X1 U895 ( .A1(G95), .A2(n680), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G107), .A2(n886), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n888), .A2(G119), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT88), .B(n804), .Z(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n610), .A2(G131), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n903) );
  AND2_X1 U903 ( .A1(G1991), .A2(n903), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n980) );
  INV_X1 U905 ( .A(n980), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n811), .A2(n826), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n829) );
  XOR2_X1 U908 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n814) );
  XNOR2_X1 U909 ( .A(KEYINPUT99), .B(n814), .ZN(n821) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n874), .ZN(n974) );
  INV_X1 U911 ( .A(n815), .ZN(n818) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n903), .ZN(n982) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U914 ( .A1(n982), .A2(n816), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n974), .A2(n819), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n821), .B(n820), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n904), .A2(n824), .ZN(n970) );
  NAND2_X1 U920 ( .A1(n825), .A2(n970), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  INV_X1 U925 ( .A(G661), .ZN(n833) );
  NAND2_X1 U926 ( .A1(G2), .A2(G15), .ZN(n832) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT102), .B(n834), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U931 ( .A(G96), .B(KEYINPUT103), .ZN(G221) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT104), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U938 ( .A(G286), .B(G301), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n840), .B(n941), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n938), .B(n841), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  NOR2_X1 U942 ( .A1(G37), .A2(n844), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT113), .B(n845), .Z(G397) );
  XNOR2_X1 U944 ( .A(G1976), .B(G2474), .ZN(n855) );
  XOR2_X1 U945 ( .A(G1971), .B(G1961), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1981), .B(G1956), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2096), .B(G2100), .Z(n857) );
  XNOR2_X1 U956 ( .A(KEYINPUT42), .B(G2678), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U962 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(G227) );
  XNOR2_X1 U964 ( .A(KEYINPUT105), .B(n864), .ZN(G319) );
  NAND2_X1 U965 ( .A1(G100), .A2(n680), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G112), .A2(n886), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n888), .A2(G124), .ZN(n867) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n867), .Z(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(KEYINPUT107), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G136), .A2(n610), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U974 ( .A(G160), .B(G162), .Z(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n902) );
  XOR2_X1 U976 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n885) );
  NAND2_X1 U979 ( .A1(n886), .A2(G115), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G127), .A2(n888), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n879), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G139), .A2(n610), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n881), .A2(n880), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n680), .A2(G103), .ZN(n882) );
  XOR2_X1 U986 ( .A(KEYINPUT110), .B(n882), .Z(n883) );
  NOR2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n985) );
  XOR2_X1 U988 ( .A(n885), .B(n985), .Z(n900) );
  NAND2_X1 U989 ( .A1(n886), .A2(G118), .ZN(n887) );
  XNOR2_X1 U990 ( .A(n887), .B(KEYINPUT108), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G130), .A2(n888), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n891), .B(KEYINPUT109), .ZN(n896) );
  NAND2_X1 U994 ( .A1(G142), .A2(n610), .ZN(n893) );
  NAND2_X1 U995 ( .A1(G106), .A2(n680), .ZN(n892) );
  NAND2_X1 U996 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U997 ( .A(KEYINPUT45), .B(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n897), .B(n978), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(G164), .B(n898), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G395) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G397), .A2(n909), .ZN(n913) );
  INV_X1 U1009 ( .A(G319), .ZN(n910) );
  NOR2_X1 U1010 ( .A1(n910), .A2(G401), .ZN(n911) );
  XNOR2_X1 U1011 ( .A(n911), .B(KEYINPUT114), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n914), .A2(G395), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(KEYINPUT115), .ZN(G225) );
  XOR2_X1 U1015 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1017 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n924) );
  XOR2_X1 U1020 ( .A(G2067), .B(G26), .Z(n918) );
  NAND2_X1 U1021 ( .A1(n918), .A2(G28), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G27), .B(n919), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(n920), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G25), .B(G1991), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1028 ( .A(KEYINPUT53), .B(n927), .Z(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(G34), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(n928), .B(KEYINPUT119), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(G2084), .B(n929), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G35), .B(G2090), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(n934), .B(KEYINPUT120), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(G29), .A2(n935), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(KEYINPUT55), .B(n936), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n937), .A2(G11), .ZN(n969) );
  XNOR2_X1 U1039 ( .A(G301), .B(G1961), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(n938), .B(G1341), .ZN(n939) );
  NOR2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(G1348), .A2(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(G1956), .B(G299), .ZN(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n950), .B(KEYINPUT122), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1051 ( .A(KEYINPUT57), .B(n953), .Z(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n963) );
  XNOR2_X1 U1053 ( .A(G1971), .B(G303), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(n956), .B(KEYINPUT123), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT124), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1059 ( .A(G16), .B(KEYINPUT121), .Z(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT56), .B(n964), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(KEYINPUT125), .B(n967), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n996) );
  INV_X1 U1064 ( .A(n970), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n992) );
  XOR2_X1 U1066 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT117), .B(n975), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n976), .B(KEYINPUT51), .ZN(n984) );
  XOR2_X1 U1070 ( .A(G2084), .B(G160), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n990) );
  XOR2_X1 U1075 ( .A(G2072), .B(n985), .Z(n987) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT50), .B(n988), .Z(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n993), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n994), .A2(G29), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XOR2_X1 U1084 ( .A(G1966), .B(G21), .Z(n1008) );
  XOR2_X1 U1085 ( .A(G4), .B(KEYINPUT126), .Z(n998) );
  XNOR2_X1 U1086 ( .A(G1348), .B(KEYINPUT59), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n998), .B(n997), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(G19), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G1956), .B(G20), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(n1006), .B(KEYINPUT60), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(KEYINPUT127), .B(n1009), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(n1010), .B(G5), .Z(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1020), .Z(n1021) );
  NOR2_X1 U1107 ( .A1(G16), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

