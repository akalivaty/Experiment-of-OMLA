//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n464), .B1(new_n461), .B2(KEYINPUT71), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G125), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT70), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(new_n475), .B1(G113), .B2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(KEYINPUT70), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n472), .B1(new_n478), .B2(G2105), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(new_n470), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n469), .B1(new_n465), .B2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n465), .B2(new_n467), .ZN(new_n490));
  AND2_X1   g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n469), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n465), .B2(new_n467), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n473), .A2(G138), .A3(new_n469), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n507), .A2(G62), .ZN(new_n515));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT74), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n514), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n513), .A2(new_n518), .ZN(G166));
  AND2_X1   g094(.A1(new_n507), .A2(new_n508), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(G89), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT75), .B(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(new_n526), .A3(G543), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT76), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT76), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G168));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n507), .B2(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n532), .B1(new_n535), .B2(new_n514), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n504), .B2(new_n506), .ZN(new_n538));
  OAI211_X1 g113(.A(KEYINPUT77), .B(G651), .C1(new_n538), .C2(new_n534), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n507), .A2(G90), .A3(new_n508), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n508), .A2(G52), .A3(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT78), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n546), .B(new_n543), .C1(new_n536), .C2(new_n539), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(G543), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n514), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n508), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT80), .B(G43), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n520), .A2(G81), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n553), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n508), .A2(new_n575), .A3(G53), .A4(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n520), .A2(G91), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(G299));
  NAND2_X1  g154(.A1(new_n530), .A2(KEYINPUT81), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n524), .B(new_n581), .C1(new_n528), .C2(new_n529), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  NAND2_X1  g160(.A1(new_n520), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n559), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n520), .A2(G86), .B1(new_n559), .B2(G48), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n507), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT82), .ZN(G305));
  AOI22_X1  g171(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT83), .ZN(new_n598));
  INV_X1    g173(.A(G72), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI221_X1 g175(.A(KEYINPUT83), .B1(new_n599), .B2(new_n502), .C1(new_n553), .C2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(G651), .A3(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n520), .A2(G85), .B1(new_n559), .B2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n553), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n559), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n520), .A2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(KEYINPUT10), .B1(new_n520), .B2(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n605), .B1(new_n615), .B2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(new_n605), .B(new_n616), .S(new_n617), .Z(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT85), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(new_n583), .B2(G868), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(new_n583), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n473), .A2(new_n462), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n469), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G135), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n633), .B1(new_n634), .B2(new_n635), .C1(new_n636), .C2(new_n470), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n632), .A2(G2100), .B1(G2096), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n638), .B(new_n639), .C1(G2100), .C2(new_n632), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT88), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT87), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND4_X1  g231(.A1(new_n646), .A2(new_n647), .A3(KEYINPUT14), .A4(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n656), .B1(new_n653), .B2(new_n657), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT89), .ZN(G401));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT90), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  XOR2_X1   g245(.A(new_n664), .B(KEYINPUT17), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n665), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n667), .B1(new_n664), .B2(new_n665), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(KEYINPUT91), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n666), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(KEYINPUT91), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n670), .B(new_n673), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT19), .Z(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(KEYINPUT20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n689), .B(KEYINPUT92), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n686), .A2(new_n687), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n684), .B(KEYINPUT19), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n688), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT93), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n692), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n692), .A2(new_n695), .A3(new_n700), .A4(new_n702), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n706), .B1(new_n704), .B2(new_n707), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n683), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n710), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n712), .A2(new_n682), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G229));
  NAND2_X1  g290(.A1(new_n483), .A2(G141), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n485), .A2(G129), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(new_n721), .B1(G105), .B2(new_n462), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n725), .B2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT27), .B(G1996), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT99), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT94), .B(G16), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G19), .ZN(new_n732));
  INV_X1    g307(.A(new_n731), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n562), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(G1341), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(G1341), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n730), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n731), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT101), .ZN(new_n742));
  INV_X1    g317(.A(G1956), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G16), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G5), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G171), .B2(new_n745), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n738), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT30), .B(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n751), .A2(new_n725), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n637), .B2(new_n725), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(new_n469), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n483), .A2(G139), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n725), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n725), .B2(G33), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n755), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n766), .B1(new_n765), .B2(new_n764), .C1(new_n727), .C2(new_n728), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n725), .A2(G35), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT100), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n487), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT29), .ZN(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n725), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(G116), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n483), .B2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n485), .A2(G128), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(KEYINPUT97), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(KEYINPUT97), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(G29), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n767), .A2(new_n773), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n745), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n745), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(G1966), .Z(new_n791));
  NOR2_X1   g366(.A1(G27), .A2(G29), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2078), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n725), .B1(new_n796), .B2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n796), .B2(G34), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G160), .B2(G29), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(G2084), .ZN(new_n800));
  NOR2_X1   g375(.A1(G4), .A2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT96), .Z(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n614), .B2(new_n745), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n803), .A2(new_n804), .B1(new_n799), .B2(G2084), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n800), .B(new_n805), .C1(new_n804), .C2(new_n803), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n788), .A2(new_n791), .A3(new_n795), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n750), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(new_n733), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n483), .A2(G131), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(G107), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(G2105), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n485), .B2(G119), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G25), .B(new_n818), .S(G29), .Z(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XOR2_X1   g395(.A(new_n819), .B(new_n820), .Z(new_n821));
  NOR2_X1   g396(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G6), .A2(G16), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT82), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n595), .B(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n824), .B1(new_n826), .B2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT95), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT32), .B(G1981), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n745), .A2(G23), .ZN(new_n833));
  INV_X1    g408(.A(G288), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n745), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT33), .B(G1976), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n733), .A2(G22), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G166), .B2(new_n733), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1971), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n831), .A2(new_n832), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n823), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n831), .A2(new_n832), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n810), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n810), .A3(new_n845), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n809), .B1(new_n847), .B2(new_n848), .ZN(G311));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n808), .B1(new_n850), .B2(new_n846), .ZN(G150));
  AOI22_X1  g426(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n514), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT102), .B(G55), .Z(new_n854));
  AOI22_X1  g429(.A1(new_n520), .A2(G93), .B1(new_n559), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n562), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n623), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g437(.A(G860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n856), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT106), .B1(new_n761), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(KEYINPUT106), .B2(new_n761), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n724), .A2(new_n500), .ZN(new_n873));
  NAND2_X1  g448(.A1(G164), .A2(new_n723), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n784), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n784), .B1(new_n873), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n879), .A2(new_n871), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT108), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n818), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n813), .A2(KEYINPUT108), .A3(new_n817), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n630), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n483), .A2(G142), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n485), .A2(G130), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n469), .A2(KEYINPUT107), .A3(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT107), .B1(new_n469), .B2(G118), .ZN(new_n890));
  OR2_X1    g465(.A1(G106), .A2(G2105), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n889), .A2(G2104), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n630), .B1(new_n883), .B2(new_n884), .ZN(new_n894));
  OR3_X1    g469(.A1(new_n886), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n886), .B2(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n881), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n880), .A3(new_n878), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G160), .B(new_n637), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G162), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  INV_X1    g479(.A(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n897), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g483(.A(new_n857), .B(new_n625), .ZN(new_n909));
  INV_X1    g484(.A(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n614), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(G299), .B(new_n609), .C1(new_n613), .C2(new_n612), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n909), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n914), .B(new_n921), .C1(new_n909), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n826), .A2(G166), .ZN(new_n923));
  NAND2_X1  g498(.A1(G305), .A2(G303), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n602), .A2(new_n834), .A3(new_n603), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n834), .B1(new_n602), .B2(new_n603), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n929), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n926), .A3(new_n927), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT110), .B1(new_n928), .B2(new_n929), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n923), .A4(new_n924), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n920), .A2(new_n922), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n920), .B2(new_n922), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n856), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n939), .B1(G868), .B2(new_n940), .ZN(G295));
  OAI21_X1  g516(.A(new_n939), .B1(G868), .B2(new_n940), .ZN(G331));
  OAI211_X1 g517(.A(new_n580), .B(new_n582), .C1(new_n545), .C2(new_n547), .ZN(new_n943));
  OAI21_X1  g518(.A(G64), .B1(new_n551), .B2(new_n552), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n533), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT77), .B1(new_n945), .B2(G651), .ZN(new_n946));
  INV_X1    g521(.A(new_n539), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n544), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n546), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n540), .A2(KEYINPUT78), .A3(new_n544), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(G168), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(KEYINPUT111), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND3_X1  g528(.A1(G301), .A2(new_n953), .A3(G168), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n952), .A2(new_n857), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n857), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n913), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n954), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n858), .ZN(new_n959));
  INV_X1    g534(.A(new_n918), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n952), .A2(new_n857), .A3(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n962), .A3(new_n936), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n904), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n936), .B1(new_n957), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT43), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n913), .A2(KEYINPUT41), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n913), .B2(new_n915), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n957), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n936), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n904), .A4(new_n963), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n955), .A2(new_n956), .A3(new_n918), .ZN(new_n979));
  INV_X1    g554(.A(new_n913), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n959), .B2(new_n961), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n971), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(new_n973), .A3(new_n904), .A4(new_n963), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n936), .B1(new_n957), .B2(new_n969), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n964), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n978), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n978), .A2(new_n986), .A3(KEYINPUT44), .A4(new_n983), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(G397));
  NAND2_X1  g564(.A1(new_n478), .A2(G2105), .ZN(new_n990));
  INV_X1    g565(.A(new_n472), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(G40), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n500), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1996), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n723), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n997), .B(KEYINPUT113), .Z(new_n1001));
  XNOR2_X1  g576(.A(new_n784), .B(G2067), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n724), .A2(new_n998), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1000), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n818), .B(new_n820), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1001), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(G290), .B(G1986), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n997), .B2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(G160), .A2(G40), .A3(new_n993), .A4(new_n500), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n590), .A2(new_n594), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G86), .ZN(new_n1016));
  INV_X1    g591(.A(G48), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n509), .A2(new_n1016), .B1(new_n511), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n514), .B1(new_n591), .B2(new_n592), .ZN(new_n1019));
  OAI21_X1  g594(.A(G1981), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1011), .B(G8), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n834), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1015), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1012), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n834), .A2(G1976), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1011), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1011), .A2(G8), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1032), .B(new_n1034), .C1(new_n1024), .C2(new_n1023), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1025), .A2(KEYINPUT116), .A3(new_n1034), .A4(new_n1032), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n990), .A2(G40), .A3(new_n991), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n993), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n996), .ZN(new_n1042));
  INV_X1    g617(.A(G1971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n500), .B2(new_n993), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n992), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n500), .A2(new_n1045), .A3(new_n993), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n772), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(KEYINPUT114), .A3(new_n1049), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G303), .A2(G8), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT55), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1052), .A2(new_n1053), .A3(G8), .A4(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1029), .B1(new_n1039), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1044), .A2(new_n1059), .A3(new_n1049), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1055), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1035), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1057), .A3(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1040), .A2(new_n794), .A3(new_n1041), .A4(new_n996), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT126), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT53), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1046), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1040), .A2(new_n1048), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n748), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(KEYINPUT126), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1065), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT62), .ZN(new_n1077));
  INV_X1    g652(.A(G2084), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1047), .A2(new_n1078), .A3(new_n1048), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1040), .A2(new_n1041), .A3(new_n996), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1079), .B(G168), .C1(new_n1080), .C2(G1966), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(G8), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(new_n1080), .B2(G1966), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(G8), .A3(new_n530), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1081), .B2(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1077), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1081), .A2(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT51), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT62), .A3(new_n1085), .A4(new_n1083), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1058), .B1(new_n1076), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1348), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1011), .A2(G2067), .ZN(new_n1095));
  NOR4_X1   g670(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT60), .A4(new_n614), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1011), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1042), .A2(G1996), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n563), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT123), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1099), .B(new_n563), .C1(KEYINPUT123), .C2(new_n1101), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1096), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n615), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1070), .A2(new_n804), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1095), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n614), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n577), .A2(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n574), .A2(new_n1113), .A3(new_n576), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1112), .A2(new_n572), .A3(new_n578), .A4(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT121), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT121), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1111), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1070), .A2(new_n743), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1040), .A2(new_n1041), .A3(new_n996), .A4(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1120), .A2(KEYINPUT124), .A3(new_n1121), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1110), .A2(KEYINPUT60), .B1(new_n1124), .B2(KEYINPUT61), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1119), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1127), .A2(new_n1117), .B1(KEYINPUT57), .B2(new_n910), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1132), .A2(KEYINPUT61), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1105), .A2(new_n1125), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1106), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT122), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1130), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1065), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1068), .A2(G301), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1075), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n1145), .B2(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1147), .B(new_n1148), .C1(new_n1075), .C2(new_n1144), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1093), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1084), .A2(G8), .A3(new_n583), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1063), .A2(new_n1057), .A3(new_n1064), .A4(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1153), .A2(KEYINPUT118), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT118), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1152), .A2(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1052), .A2(G8), .A3(new_n1053), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1055), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1160));
  AND4_X1   g735(.A1(new_n1057), .A2(new_n1157), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1155), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1010), .B1(new_n1151), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1002), .A2(new_n723), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1007), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT47), .Z(new_n1167));
  NAND4_X1  g742(.A1(new_n1005), .A2(new_n820), .A3(new_n813), .A4(new_n817), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n784), .A2(G2067), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1007), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n997), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT48), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1008), .A2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1167), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1163), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g751(.A(new_n680), .B(G319), .C1(new_n659), .C2(new_n660), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n711), .B2(new_n713), .ZN(new_n1179));
  AND2_X1   g753(.A1(new_n907), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g754(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(KEYINPUT127), .B1(new_n975), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n1181), .A2(new_n1182), .ZN(G308));
  NAND2_X1  g757(.A1(new_n975), .A2(new_n1180), .ZN(G225));
endmodule


