

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U545 ( .A(KEYINPUT17), .B(n512), .Z(n960) );
  NAND2_X1 U546 ( .A1(n691), .A2(n844), .ZN(n692) );
  XOR2_X1 U547 ( .A(n740), .B(KEYINPUT97), .Z(n509) );
  XNOR2_X1 U548 ( .A(n716), .B(KEYINPUT94), .ZN(n510) );
  AND2_X1 U549 ( .A1(n753), .A2(n752), .ZN(n511) );
  XNOR2_X1 U550 ( .A(n693), .B(KEYINPUT90), .ZN(n691) );
  INV_X1 U551 ( .A(n717), .ZN(n693) );
  INV_X1 U552 ( .A(KEYINPUT28), .ZN(n671) );
  INV_X1 U553 ( .A(KEYINPUT92), .ZN(n696) );
  INV_X1 U554 ( .A(KEYINPUT29), .ZN(n689) );
  XNOR2_X1 U555 ( .A(n690), .B(n689), .ZN(n699) );
  INV_X1 U556 ( .A(n710), .ZN(n711) );
  XNOR2_X1 U557 ( .A(n712), .B(KEYINPUT95), .ZN(n713) );
  NAND2_X1 U558 ( .A1(n755), .A2(n665), .ZN(n717) );
  NOR2_X1 U559 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n755) );
  INV_X1 U561 ( .A(G2105), .ZN(n516) );
  NOR2_X1 U562 ( .A1(G651), .A2(n606), .ZN(n630) );
  AND2_X1 U563 ( .A1(n516), .A2(G2104), .ZN(n959) );
  XNOR2_X1 U564 ( .A(n517), .B(KEYINPUT64), .ZN(n967) );
  NOR2_X1 U565 ( .A1(n521), .A2(n520), .ZN(G160) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n512) );
  NAND2_X1 U567 ( .A1(n960), .A2(G137), .ZN(n515) );
  NAND2_X1 U568 ( .A1(G101), .A2(n959), .ZN(n513) );
  XOR2_X1 U569 ( .A(KEYINPUT23), .B(n513), .Z(n514) );
  NAND2_X1 U570 ( .A1(n515), .A2(n514), .ZN(n521) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n966) );
  NAND2_X1 U572 ( .A1(G113), .A2(n966), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n516), .A2(G2104), .ZN(n517) );
  NAND2_X1 U574 ( .A1(G125), .A2(n967), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n519), .A2(n518), .ZN(n520) );
  INV_X1 U576 ( .A(G651), .ZN(n524) );
  NOR2_X1 U577 ( .A1(G543), .A2(n524), .ZN(n522) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n522), .Z(n629) );
  NAND2_X1 U579 ( .A1(n629), .A2(G64), .ZN(n523) );
  XNOR2_X1 U580 ( .A(KEYINPUT65), .B(n523), .ZN(n532) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U582 ( .A1(G90), .A2(n633), .ZN(n526) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n606) );
  NOR2_X1 U584 ( .A1(n606), .A2(n524), .ZN(n634) );
  NAND2_X1 U585 ( .A1(G77), .A2(n634), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U587 ( .A(n527), .B(KEYINPUT9), .ZN(n528) );
  XNOR2_X1 U588 ( .A(n528), .B(KEYINPUT66), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n630), .A2(G52), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n532), .A2(n531), .ZN(G171) );
  NAND2_X1 U592 ( .A1(G138), .A2(n960), .ZN(n534) );
  NAND2_X1 U593 ( .A1(G102), .A2(n959), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U595 ( .A1(G114), .A2(n966), .ZN(n536) );
  NAND2_X1 U596 ( .A1(G126), .A2(n967), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U599 ( .A1(G85), .A2(n633), .ZN(n540) );
  NAND2_X1 U600 ( .A1(G72), .A2(n634), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G60), .A2(n629), .ZN(n542) );
  NAND2_X1 U603 ( .A1(G47), .A2(n630), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  OR2_X1 U605 ( .A1(n544), .A2(n543), .ZN(G290) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G132), .ZN(G219) );
  INV_X1 U608 ( .A(G82), .ZN(G220) );
  INV_X1 U609 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U610 ( .A(KEYINPUT72), .B(KEYINPUT6), .ZN(n548) );
  NAND2_X1 U611 ( .A1(G63), .A2(n629), .ZN(n546) );
  NAND2_X1 U612 ( .A1(G51), .A2(n630), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n633), .A2(G89), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G76), .A2(n634), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(KEYINPUT5), .B(n552), .Z(n553) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n556) );
  XNOR2_X1 U621 ( .A(KEYINPUT73), .B(KEYINPUT7), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(n557), .ZN(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT68), .ZN(n559) );
  XNOR2_X1 U627 ( .A(KEYINPUT10), .B(n559), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n804) );
  NAND2_X1 U629 ( .A1(n804), .A2(G567), .ZN(n560) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U631 ( .A1(n633), .A2(G81), .ZN(n561) );
  XNOR2_X1 U632 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U633 ( .A1(G68), .A2(n634), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n564), .Z(n568) );
  NAND2_X1 U636 ( .A1(G56), .A2(n629), .ZN(n565) );
  XNOR2_X1 U637 ( .A(n565), .B(KEYINPUT69), .ZN(n566) );
  XNOR2_X1 U638 ( .A(n566), .B(KEYINPUT14), .ZN(n567) );
  NOR2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n630), .A2(G43), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n990) );
  INV_X1 U642 ( .A(G860), .ZN(n935) );
  OR2_X1 U643 ( .A1(n990), .A2(n935), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G79), .A2(n634), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n571), .B(KEYINPUT70), .ZN(n578) );
  NAND2_X1 U647 ( .A1(G92), .A2(n633), .ZN(n573) );
  NAND2_X1 U648 ( .A1(G66), .A2(n629), .ZN(n572) );
  NAND2_X1 U649 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G54), .A2(n630), .ZN(n574) );
  XNOR2_X1 U651 ( .A(KEYINPUT71), .B(n574), .ZN(n575) );
  NOR2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U654 ( .A(KEYINPUT15), .B(n579), .ZN(n989) );
  INV_X1 U655 ( .A(n989), .ZN(n875) );
  INV_X1 U656 ( .A(G868), .ZN(n648) );
  NAND2_X1 U657 ( .A1(n875), .A2(n648), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G65), .A2(n629), .ZN(n583) );
  NAND2_X1 U660 ( .A1(G53), .A2(n630), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U662 ( .A1(G91), .A2(n633), .ZN(n585) );
  NAND2_X1 U663 ( .A1(G78), .A2(n634), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n886) );
  INV_X1 U666 ( .A(n886), .ZN(G299) );
  NAND2_X1 U667 ( .A1(G868), .A2(G286), .ZN(n589) );
  NAND2_X1 U668 ( .A1(G299), .A2(n648), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n935), .A2(G559), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n590), .A2(n989), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n591), .B(KEYINPUT16), .ZN(n592) );
  XOR2_X1 U673 ( .A(KEYINPUT75), .B(n592), .Z(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n990), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n989), .A2(G868), .ZN(n593) );
  NOR2_X1 U676 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U677 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U678 ( .A1(G99), .A2(n959), .ZN(n597) );
  NAND2_X1 U679 ( .A1(G135), .A2(n960), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n967), .A2(G123), .ZN(n598) );
  XNOR2_X1 U682 ( .A(n598), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U683 ( .A1(G111), .A2(n966), .ZN(n599) );
  XNOR2_X1 U684 ( .A(n599), .B(KEYINPUT76), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(n974) );
  XNOR2_X1 U687 ( .A(G2096), .B(n974), .ZN(n605) );
  INV_X1 U688 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G87), .A2(n606), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G49), .A2(n630), .ZN(n608) );
  NAND2_X1 U692 ( .A1(G74), .A2(G651), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n629), .A2(n609), .ZN(n610) );
  XOR2_X1 U695 ( .A(KEYINPUT79), .B(n610), .Z(n611) );
  NAND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U698 ( .A1(G88), .A2(n633), .ZN(n615) );
  NAND2_X1 U699 ( .A1(G75), .A2(n634), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G62), .A2(n629), .ZN(n617) );
  NAND2_X1 U702 ( .A1(G50), .A2(n630), .ZN(n616) );
  NAND2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U704 ( .A1(n619), .A2(n618), .ZN(G166) );
  INV_X1 U705 ( .A(G166), .ZN(G303) );
  NAND2_X1 U706 ( .A1(G73), .A2(n634), .ZN(n620) );
  XNOR2_X1 U707 ( .A(n620), .B(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G86), .A2(n633), .ZN(n622) );
  NAND2_X1 U709 ( .A1(G61), .A2(n629), .ZN(n621) );
  NAND2_X1 U710 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U711 ( .A1(G48), .A2(n630), .ZN(n623) );
  XNOR2_X1 U712 ( .A(KEYINPUT81), .B(n623), .ZN(n624) );
  NOR2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G559), .A2(n989), .ZN(n628) );
  XOR2_X1 U716 ( .A(n990), .B(n628), .Z(n934) );
  NAND2_X1 U717 ( .A1(G67), .A2(n629), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G55), .A2(n630), .ZN(n631) );
  NAND2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n639) );
  NAND2_X1 U720 ( .A1(G93), .A2(n633), .ZN(n636) );
  NAND2_X1 U721 ( .A1(G80), .A2(n634), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U723 ( .A(KEYINPUT77), .B(n637), .Z(n638) );
  NOR2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U725 ( .A(KEYINPUT78), .B(n640), .Z(n936) );
  XNOR2_X1 U726 ( .A(KEYINPUT19), .B(G303), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n641), .B(G305), .ZN(n642) );
  XNOR2_X1 U728 ( .A(n936), .B(n642), .ZN(n644) );
  XNOR2_X1 U729 ( .A(G290), .B(n886), .ZN(n643) );
  XNOR2_X1 U730 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U731 ( .A(G288), .B(n645), .ZN(n991) );
  XOR2_X1 U732 ( .A(n934), .B(n991), .Z(n646) );
  XNOR2_X1 U733 ( .A(KEYINPUT82), .B(n646), .ZN(n647) );
  NOR2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n650) );
  NOR2_X1 U735 ( .A1(n936), .A2(G868), .ZN(n649) );
  NOR2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n651) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n651), .Z(n652) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n652), .ZN(n653) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n653), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n654), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G120), .A2(G108), .ZN(n655) );
  NOR2_X1 U745 ( .A1(G237), .A2(n655), .ZN(n656) );
  NAND2_X1 U746 ( .A1(G69), .A2(n656), .ZN(n810) );
  NAND2_X1 U747 ( .A1(n810), .A2(G567), .ZN(n661) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n657) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n657), .Z(n658) );
  NOR2_X1 U750 ( .A1(G218), .A2(n658), .ZN(n659) );
  NAND2_X1 U751 ( .A1(G96), .A2(n659), .ZN(n811) );
  NAND2_X1 U752 ( .A1(n811), .A2(G2106), .ZN(n660) );
  NAND2_X1 U753 ( .A1(n661), .A2(n660), .ZN(n958) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n662) );
  XOR2_X1 U755 ( .A(KEYINPUT83), .B(n662), .Z(n663) );
  NOR2_X1 U756 ( .A1(n958), .A2(n663), .ZN(n809) );
  NAND2_X1 U757 ( .A1(G36), .A2(n809), .ZN(n664) );
  XNOR2_X1 U758 ( .A(n664), .B(KEYINPUT84), .ZN(G176) );
  AND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n665) );
  NOR2_X1 U760 ( .A1(G2084), .A2(n717), .ZN(n700) );
  NAND2_X1 U761 ( .A1(G8), .A2(n700), .ZN(n714) );
  INV_X1 U762 ( .A(n691), .ZN(n666) );
  NAND2_X1 U763 ( .A1(n666), .A2(G1956), .ZN(n667) );
  XNOR2_X1 U764 ( .A(KEYINPUT93), .B(n667), .ZN(n670) );
  NAND2_X1 U765 ( .A1(G2072), .A2(n691), .ZN(n668) );
  XNOR2_X1 U766 ( .A(KEYINPUT27), .B(n668), .ZN(n669) );
  NOR2_X1 U767 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U768 ( .A1(n886), .A2(n673), .ZN(n672) );
  XNOR2_X1 U769 ( .A(n672), .B(n671), .ZN(n688) );
  NAND2_X1 U770 ( .A1(n886), .A2(n673), .ZN(n686) );
  INV_X1 U771 ( .A(G1996), .ZN(n845) );
  NOR2_X1 U772 ( .A1(n717), .A2(n845), .ZN(n674) );
  XOR2_X1 U773 ( .A(n674), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U774 ( .A1(n717), .A2(G1341), .ZN(n675) );
  NAND2_X1 U775 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U776 ( .A1(n990), .A2(n677), .ZN(n678) );
  OR2_X1 U777 ( .A1(n989), .A2(n678), .ZN(n684) );
  NAND2_X1 U778 ( .A1(n989), .A2(n678), .ZN(n682) );
  NAND2_X1 U779 ( .A1(G2067), .A2(n691), .ZN(n680) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n717), .ZN(n679) );
  NAND2_X1 U781 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U782 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U783 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U784 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U785 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .ZN(n844) );
  XNOR2_X1 U787 ( .A(n692), .B(KEYINPUT91), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n693), .A2(G1961), .ZN(n694) );
  NOR2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U790 ( .A(n697), .B(n696), .ZN(n704) );
  NAND2_X1 U791 ( .A1(G171), .A2(n704), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n709) );
  NAND2_X1 U793 ( .A1(G8), .A2(n717), .ZN(n751) );
  NOR2_X1 U794 ( .A1(G1966), .A2(n751), .ZN(n710) );
  NOR2_X1 U795 ( .A1(n700), .A2(n710), .ZN(n701) );
  NAND2_X1 U796 ( .A1(G8), .A2(n701), .ZN(n702) );
  XNOR2_X1 U797 ( .A(KEYINPUT30), .B(n702), .ZN(n703) );
  NOR2_X1 U798 ( .A1(G168), .A2(n703), .ZN(n706) );
  NOR2_X1 U799 ( .A1(n704), .A2(G171), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U801 ( .A(KEYINPUT31), .B(n707), .Z(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n716) );
  NAND2_X1 U803 ( .A1(n510), .A2(n711), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n746) );
  AND2_X1 U805 ( .A1(G286), .A2(G8), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n725) );
  INV_X1 U807 ( .A(G8), .ZN(n723) );
  NOR2_X1 U808 ( .A1(G1971), .A2(n751), .ZN(n719) );
  NOR2_X1 U809 ( .A1(G2090), .A2(n717), .ZN(n718) );
  NOR2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n720), .A2(G303), .ZN(n721) );
  XNOR2_X1 U812 ( .A(n721), .B(KEYINPUT96), .ZN(n722) );
  OR2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  AND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U815 ( .A(n726), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U816 ( .A1(G1976), .A2(G288), .ZN(n870) );
  AND2_X1 U817 ( .A1(n745), .A2(n870), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n746), .A2(n727), .ZN(n734) );
  INV_X1 U819 ( .A(n870), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n735) );
  NOR2_X1 U821 ( .A1(G1971), .A2(G303), .ZN(n728) );
  NOR2_X1 U822 ( .A1(n735), .A2(n728), .ZN(n871) );
  OR2_X1 U823 ( .A1(n729), .A2(n871), .ZN(n730) );
  OR2_X1 U824 ( .A1(n751), .A2(n730), .ZN(n732) );
  INV_X1 U825 ( .A(KEYINPUT33), .ZN(n731) );
  AND2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U827 ( .A1(n734), .A2(n733), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n735), .A2(KEYINPUT33), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n736), .A2(n751), .ZN(n737) );
  XOR2_X1 U830 ( .A(G1981), .B(G305), .Z(n882) );
  NAND2_X1 U831 ( .A1(n739), .A2(n882), .ZN(n740) );
  NOR2_X1 U832 ( .A1(G1981), .A2(G305), .ZN(n741) );
  XOR2_X1 U833 ( .A(n741), .B(KEYINPUT24), .Z(n742) );
  XNOR2_X1 U834 ( .A(KEYINPUT88), .B(n742), .ZN(n743) );
  NOR2_X1 U835 ( .A1(n751), .A2(n743), .ZN(n744) );
  XNOR2_X1 U836 ( .A(n744), .B(KEYINPUT89), .ZN(n753) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n749) );
  NOR2_X1 U838 ( .A1(G2090), .A2(G303), .ZN(n747) );
  NAND2_X1 U839 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n509), .A2(n511), .ZN(n788) );
  NAND2_X1 U843 ( .A1(G160), .A2(G40), .ZN(n754) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n799) );
  NAND2_X1 U845 ( .A1(G104), .A2(n959), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G140), .A2(n960), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U848 ( .A(KEYINPUT34), .B(n758), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G116), .A2(n966), .ZN(n760) );
  NAND2_X1 U850 ( .A1(G128), .A2(n967), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U852 ( .A(KEYINPUT86), .B(n761), .Z(n762) );
  XNOR2_X1 U853 ( .A(KEYINPUT35), .B(n762), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U855 ( .A(KEYINPUT36), .B(n765), .ZN(n981) );
  XNOR2_X1 U856 ( .A(G2067), .B(KEYINPUT37), .ZN(n797) );
  NOR2_X1 U857 ( .A1(n981), .A2(n797), .ZN(n917) );
  NAND2_X1 U858 ( .A1(n799), .A2(n917), .ZN(n795) );
  INV_X1 U859 ( .A(n795), .ZN(n786) );
  NAND2_X1 U860 ( .A1(G141), .A2(n960), .ZN(n767) );
  NAND2_X1 U861 ( .A1(G117), .A2(n966), .ZN(n766) );
  NAND2_X1 U862 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U863 ( .A1(n959), .A2(G105), .ZN(n768) );
  XOR2_X1 U864 ( .A(KEYINPUT38), .B(n768), .Z(n769) );
  NOR2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U866 ( .A1(G129), .A2(n967), .ZN(n771) );
  NAND2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n978) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n978), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G95), .A2(n959), .ZN(n774) );
  NAND2_X1 U870 ( .A1(G131), .A2(n960), .ZN(n773) );
  NAND2_X1 U871 ( .A1(n774), .A2(n773), .ZN(n778) );
  NAND2_X1 U872 ( .A1(G107), .A2(n966), .ZN(n776) );
  NAND2_X1 U873 ( .A1(G119), .A2(n967), .ZN(n775) );
  NAND2_X1 U874 ( .A1(n776), .A2(n775), .ZN(n777) );
  OR2_X1 U875 ( .A1(n778), .A2(n777), .ZN(n984) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n984), .ZN(n779) );
  NAND2_X1 U877 ( .A1(n780), .A2(n779), .ZN(n913) );
  NAND2_X1 U878 ( .A1(n913), .A2(n799), .ZN(n781) );
  XNOR2_X1 U879 ( .A(n781), .B(KEYINPUT87), .ZN(n792) );
  INV_X1 U880 ( .A(n792), .ZN(n784) );
  XNOR2_X1 U881 ( .A(G1986), .B(G290), .ZN(n890) );
  NAND2_X1 U882 ( .A1(n890), .A2(n799), .ZN(n782) );
  XOR2_X1 U883 ( .A(KEYINPUT85), .B(n782), .Z(n783) );
  NAND2_X1 U884 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n788), .A2(n787), .ZN(n802) );
  NOR2_X1 U887 ( .A1(n978), .A2(G1996), .ZN(n789) );
  XNOR2_X1 U888 ( .A(n789), .B(KEYINPUT98), .ZN(n921) );
  NOR2_X1 U889 ( .A1(G1991), .A2(n984), .ZN(n910) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n790) );
  NOR2_X1 U891 ( .A1(n910), .A2(n790), .ZN(n791) );
  NOR2_X1 U892 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U893 ( .A1(n921), .A2(n793), .ZN(n794) );
  XNOR2_X1 U894 ( .A(KEYINPUT39), .B(n794), .ZN(n796) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n981), .A2(n797), .ZN(n924) );
  NAND2_X1 U897 ( .A1(n798), .A2(n924), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n804), .ZN(G217) );
  NAND2_X1 U902 ( .A1(G15), .A2(G2), .ZN(n805) );
  XOR2_X1 U903 ( .A(KEYINPUT100), .B(n805), .Z(n806) );
  NAND2_X1 U904 ( .A1(n806), .A2(G661), .ZN(n807) );
  XOR2_X1 U905 ( .A(KEYINPUT101), .B(n807), .Z(G259) );
  NAND2_X1 U906 ( .A1(G3), .A2(G1), .ZN(n808) );
  NAND2_X1 U907 ( .A1(n809), .A2(n808), .ZN(G188) );
  XOR2_X1 U908 ( .A(G96), .B(KEYINPUT102), .Z(G221) );
  NOR2_X1 U909 ( .A1(n811), .A2(n810), .ZN(G325) );
  XNOR2_X1 U910 ( .A(KEYINPUT103), .B(G325), .ZN(G261) );
  XNOR2_X1 U911 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  NAND2_X1 U913 ( .A1(G100), .A2(n959), .ZN(n813) );
  NAND2_X1 U914 ( .A1(G112), .A2(n966), .ZN(n812) );
  NAND2_X1 U915 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U916 ( .A(n814), .B(KEYINPUT107), .ZN(n816) );
  NAND2_X1 U917 ( .A1(G136), .A2(n960), .ZN(n815) );
  NAND2_X1 U918 ( .A1(n816), .A2(n815), .ZN(n819) );
  NAND2_X1 U919 ( .A1(n967), .A2(G124), .ZN(n817) );
  XOR2_X1 U920 ( .A(KEYINPUT44), .B(n817), .Z(n818) );
  NOR2_X1 U921 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U922 ( .A(KEYINPUT108), .B(n820), .ZN(G162) );
  XNOR2_X1 U923 ( .A(G1966), .B(G21), .ZN(n822) );
  XNOR2_X1 U924 ( .A(G5), .B(G1961), .ZN(n821) );
  NOR2_X1 U925 ( .A1(n822), .A2(n821), .ZN(n832) );
  XOR2_X1 U926 ( .A(G1348), .B(KEYINPUT59), .Z(n823) );
  XNOR2_X1 U927 ( .A(G4), .B(n823), .ZN(n825) );
  XNOR2_X1 U928 ( .A(G20), .B(G1956), .ZN(n824) );
  NOR2_X1 U929 ( .A1(n825), .A2(n824), .ZN(n829) );
  XNOR2_X1 U930 ( .A(G1341), .B(G19), .ZN(n827) );
  XNOR2_X1 U931 ( .A(G6), .B(G1981), .ZN(n826) );
  NOR2_X1 U932 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U933 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U934 ( .A(KEYINPUT60), .B(n830), .Z(n831) );
  NAND2_X1 U935 ( .A1(n832), .A2(n831), .ZN(n840) );
  XNOR2_X1 U936 ( .A(G1986), .B(G24), .ZN(n834) );
  XNOR2_X1 U937 ( .A(G23), .B(G1976), .ZN(n833) );
  NOR2_X1 U938 ( .A1(n834), .A2(n833), .ZN(n837) );
  XNOR2_X1 U939 ( .A(G1971), .B(KEYINPUT125), .ZN(n835) );
  XNOR2_X1 U940 ( .A(n835), .B(G22), .ZN(n836) );
  NAND2_X1 U941 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U942 ( .A(KEYINPUT58), .B(n838), .ZN(n839) );
  NOR2_X1 U943 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U944 ( .A(KEYINPUT61), .B(n841), .Z(n843) );
  XNOR2_X1 U945 ( .A(KEYINPUT124), .B(G16), .ZN(n842) );
  NOR2_X1 U946 ( .A1(n843), .A2(n842), .ZN(n868) );
  XOR2_X1 U947 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n865) );
  XNOR2_X1 U948 ( .A(G2090), .B(G35), .ZN(n859) );
  XNOR2_X1 U949 ( .A(G27), .B(n844), .ZN(n851) );
  XNOR2_X1 U950 ( .A(G32), .B(n845), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n846), .A2(G28), .ZN(n849) );
  XNOR2_X1 U952 ( .A(G25), .B(G1991), .ZN(n847) );
  XNOR2_X1 U953 ( .A(KEYINPUT116), .B(n847), .ZN(n848) );
  NOR2_X1 U954 ( .A1(n849), .A2(n848), .ZN(n850) );
  NAND2_X1 U955 ( .A1(n851), .A2(n850), .ZN(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G26), .ZN(n853) );
  XNOR2_X1 U957 ( .A(G2072), .B(G33), .ZN(n852) );
  NOR2_X1 U958 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n854), .B(KEYINPUT117), .ZN(n855) );
  NOR2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U961 ( .A(KEYINPUT53), .B(n857), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n863) );
  XOR2_X1 U963 ( .A(G34), .B(KEYINPUT118), .Z(n861) );
  XNOR2_X1 U964 ( .A(G2084), .B(KEYINPUT54), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n861), .B(n860), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  NOR2_X1 U968 ( .A1(G29), .A2(n866), .ZN(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G11), .A2(n869), .ZN(n898) );
  XOR2_X1 U971 ( .A(G16), .B(KEYINPUT56), .Z(n896) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n873) );
  AND2_X1 U973 ( .A1(G303), .A2(G1971), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(KEYINPUT123), .B(n874), .Z(n880) );
  XNOR2_X1 U976 ( .A(G301), .B(G1961), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n875), .B(G1348), .ZN(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U979 ( .A(KEYINPUT122), .B(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n894) );
  XNOR2_X1 U981 ( .A(G1966), .B(G168), .ZN(n881) );
  XNOR2_X1 U982 ( .A(n881), .B(KEYINPUT120), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n885) );
  XOR2_X1 U984 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n892) );
  XOR2_X1 U986 ( .A(n990), .B(G1341), .Z(n888) );
  XNOR2_X1 U987 ( .A(n886), .B(G1956), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U989 ( .A1(n890), .A2(n889), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  NOR2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(KEYINPUT126), .ZN(n932) );
  NAND2_X1 U995 ( .A1(G103), .A2(n959), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G139), .A2(n960), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n906) );
  NAND2_X1 U998 ( .A1(G115), .A2(n966), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G127), .A2(n967), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n983) );
  XOR2_X1 U1003 ( .A(G2072), .B(n983), .Z(n908) );
  XOR2_X1 U1004 ( .A(G164), .B(G2078), .Z(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT50), .B(n909), .ZN(n919) );
  NOR2_X1 U1007 ( .A1(n910), .A2(n974), .ZN(n915) );
  XOR2_X1 U1008 ( .A(G160), .B(G2084), .Z(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT114), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n922), .Z(n923) );
  NAND2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1019 ( .A(KEYINPUT52), .B(n927), .Z(n928) );
  NOR2_X1 U1020 ( .A1(KEYINPUT55), .A2(n928), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(n929), .ZN(n930) );
  NAND2_X1 U1022 ( .A1(n930), .A2(G29), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1024 ( .A(KEYINPUT62), .B(n933), .Z(G311) );
  XNOR2_X1 U1025 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NAND2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(n937), .B(n936), .ZN(G145) );
  INV_X1 U1028 ( .A(G120), .ZN(G236) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1030 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n939) );
  XNOR2_X1 U1031 ( .A(G2678), .B(KEYINPUT105), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n939), .B(n938), .ZN(n940) );
  XOR2_X1 U1033 ( .A(n940), .B(G2100), .Z(n942) );
  XNOR2_X1 U1034 ( .A(G2084), .B(G2072), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n942), .B(n941), .ZN(n946) );
  XOR2_X1 U1036 ( .A(KEYINPUT43), .B(G2096), .Z(n944) );
  XNOR2_X1 U1037 ( .A(G2090), .B(KEYINPUT106), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n944), .B(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(n946), .B(n945), .Z(n948) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G2078), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n948), .B(n947), .ZN(G227) );
  XOR2_X1 U1042 ( .A(G1971), .B(G1956), .Z(n950) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G1961), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n950), .B(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(n951), .B(KEYINPUT41), .Z(n953) );
  XNOR2_X1 U1046 ( .A(G1986), .B(G1976), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G2474), .B(G1981), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G1991), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(n955), .B(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n957), .B(n956), .ZN(G229) );
  INV_X1 U1052 ( .A(n958), .ZN(G319) );
  XNOR2_X1 U1053 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(G106), .A2(n959), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(G142), .A2(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(KEYINPUT45), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n965), .B(n964), .ZN(n971) );
  NAND2_X1 U1059 ( .A1(G118), .A2(n966), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(G130), .A2(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G160), .B(n974), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G162), .B(n975), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(n980) );
  XNOR2_X1 U1068 ( .A(n978), .B(KEYINPUT46), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n980), .B(n979), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n982), .B(n981), .ZN(n987) );
  XNOR2_X1 U1071 ( .A(G164), .B(n983), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(n985), .B(n984), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(n987), .B(n986), .ZN(n988) );
  NOR2_X1 U1074 ( .A1(G37), .A2(n988), .ZN(G395) );
  XNOR2_X1 U1075 ( .A(n989), .B(G286), .ZN(n994) );
  XNOR2_X1 U1076 ( .A(G301), .B(n990), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(n994), .B(n993), .ZN(n995) );
  NOR2_X1 U1079 ( .A1(G37), .A2(n995), .ZN(G397) );
  NOR2_X1 U1080 ( .A1(G227), .A2(G229), .ZN(n997) );
  XNOR2_X1 U1081 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(n997), .B(n996), .ZN(n1009) );
  XOR2_X1 U1083 ( .A(G2443), .B(G2430), .Z(n999) );
  XNOR2_X1 U1084 ( .A(G1348), .B(G2451), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n999), .B(n998), .ZN(n1006) );
  XOR2_X1 U1086 ( .A(G2438), .B(KEYINPUT99), .Z(n1001) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G2454), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(n1002), .B(G2435), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(G2446), .B(G2427), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1004), .B(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1007), .A2(G14), .ZN(n1012) );
  NAND2_X1 U1094 ( .A1(G319), .A2(n1012), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NOR2_X1 U1096 ( .A1(G395), .A2(G397), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(G225) );
  INV_X1 U1098 ( .A(G225), .ZN(G308) );
  INV_X1 U1099 ( .A(n1012), .ZN(G401) );
endmodule

