

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741;

  BUF_X1 U375 ( .A(n645), .Z(n353) );
  NOR2_X1 U376 ( .A1(n434), .A2(n631), .ZN(n433) );
  XNOR2_X1 U377 ( .A(n598), .B(n597), .ZN(n645) );
  NOR2_X1 U378 ( .A1(G902), .A2(n696), .ZN(n524) );
  NAND2_X2 U379 ( .A1(n410), .A2(n409), .ZN(n606) );
  NAND2_X1 U380 ( .A1(n352), .A2(n592), .ZN(n391) );
  NAND2_X1 U381 ( .A1(n394), .A2(n393), .ZN(n352) );
  XNOR2_X1 U382 ( .A(n464), .B(n443), .ZN(n712) );
  INV_X2 U383 ( .A(G953), .ZN(n691) );
  XNOR2_X2 U384 ( .A(G119), .B(KEYINPUT72), .ZN(n390) );
  XNOR2_X2 U385 ( .A(n373), .B(n396), .ZN(n405) );
  XNOR2_X2 U386 ( .A(n541), .B(n525), .ZN(n663) );
  AND2_X1 U387 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U388 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U389 ( .A1(n653), .A2(n440), .ZN(n654) );
  NAND2_X1 U390 ( .A1(n365), .A2(n581), .ZN(n373) );
  XNOR2_X1 U391 ( .A(n537), .B(n424), .ZN(n738) );
  NOR2_X1 U392 ( .A1(n534), .A2(n594), .ZN(n633) );
  XNOR2_X1 U393 ( .A(n554), .B(n553), .ZN(n577) );
  XNOR2_X1 U394 ( .A(n422), .B(n359), .ZN(n586) );
  XOR2_X1 U395 ( .A(n625), .B(KEYINPUT62), .Z(n626) );
  XNOR2_X1 U396 ( .A(n725), .B(n521), .ZN(n696) );
  NAND2_X2 U397 ( .A1(n379), .A2(n378), .ZN(n688) );
  XNOR2_X1 U398 ( .A(n402), .B(n545), .ZN(n570) );
  NOR2_X1 U399 ( .A1(n738), .A2(n737), .ZN(n402) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n468) );
  XNOR2_X1 U401 ( .A(n414), .B(G125), .ZN(n475) );
  INV_X1 U402 ( .A(G146), .ZN(n414) );
  NOR2_X1 U403 ( .A1(n586), .A2(n529), .ZN(n512) );
  INV_X1 U404 ( .A(G137), .ZN(n452) );
  INV_X1 U405 ( .A(KEYINPUT45), .ZN(n415) );
  XNOR2_X1 U406 ( .A(n475), .B(n413), .ZN(n726) );
  XNOR2_X1 U407 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n413) );
  NAND2_X1 U408 ( .A1(G234), .A2(G237), .ZN(n506) );
  AND2_X1 U409 ( .A1(n371), .A2(n370), .ZN(n367) );
  NAND2_X1 U410 ( .A1(n382), .A2(n372), .ZN(n370) );
  NAND2_X1 U411 ( .A1(n688), .A2(n372), .ZN(n371) );
  XNOR2_X1 U412 ( .A(n411), .B(n481), .ZN(n562) );
  OR2_X1 U413 ( .A1(n609), .A2(G902), .ZN(n411) );
  XNOR2_X1 U414 ( .A(n391), .B(KEYINPUT107), .ZN(n434) );
  INV_X1 U415 ( .A(n633), .ZN(n393) );
  NOR2_X1 U416 ( .A1(n570), .A2(n647), .ZN(n376) );
  XNOR2_X1 U417 ( .A(n428), .B(n427), .ZN(n496) );
  INV_X1 U418 ( .A(KEYINPUT8), .ZN(n427) );
  NAND2_X1 U419 ( .A1(n691), .A2(G234), .ZN(n428) );
  XOR2_X1 U420 ( .A(G146), .B(KEYINPUT83), .Z(n518) );
  XNOR2_X1 U421 ( .A(n420), .B(n713), .ZN(n520) );
  XNOR2_X1 U422 ( .A(n457), .B(n442), .ZN(n420) );
  XOR2_X1 U423 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n442) );
  INV_X1 U424 ( .A(KEYINPUT33), .ZN(n385) );
  NAND2_X1 U425 ( .A1(n599), .A2(n385), .ZN(n383) );
  INV_X1 U426 ( .A(KEYINPUT1), .ZN(n525) );
  XNOR2_X1 U427 ( .A(n583), .B(n363), .ZN(n587) );
  XNOR2_X1 U428 ( .A(n439), .B(n437), .ZN(n464) );
  XNOR2_X1 U429 ( .A(n438), .B(G116), .ZN(n437) );
  XNOR2_X1 U430 ( .A(n390), .B(n389), .ZN(n439) );
  INV_X1 U431 ( .A(KEYINPUT3), .ZN(n438) );
  XNOR2_X1 U432 ( .A(n419), .B(G107), .ZN(n713) );
  XNOR2_X1 U433 ( .A(G110), .B(G104), .ZN(n419) );
  XOR2_X1 U434 ( .A(G140), .B(KEYINPUT69), .Z(n516) );
  XOR2_X1 U435 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n493) );
  XNOR2_X1 U436 ( .A(G119), .B(G128), .ZN(n491) );
  INV_X1 U437 ( .A(G134), .ZN(n454) );
  XNOR2_X1 U438 ( .A(n478), .B(n726), .ZN(n479) );
  NOR2_X1 U439 ( .A1(n604), .A2(n652), .ZN(n409) );
  XNOR2_X1 U440 ( .A(n604), .B(KEYINPUT90), .ZN(n730) );
  XNOR2_X1 U441 ( .A(n401), .B(KEYINPUT39), .ZN(n572) );
  NAND2_X1 U442 ( .A1(n356), .A2(n406), .ZN(n401) );
  NAND2_X1 U443 ( .A1(n369), .A2(n368), .ZN(n366) );
  NOR2_X1 U444 ( .A1(n382), .A2(n372), .ZN(n368) );
  INV_X1 U445 ( .A(n688), .ZN(n369) );
  NOR2_X1 U446 ( .A1(n562), .A2(n561), .ZN(n581) );
  OR2_X1 U447 ( .A1(n707), .A2(G902), .ZN(n422) );
  INV_X1 U448 ( .A(n562), .ZN(n556) );
  NOR2_X2 U449 ( .A1(n577), .A2(n576), .ZN(n418) );
  XOR2_X1 U450 ( .A(KEYINPUT68), .B(G131), .Z(n476) );
  INV_X1 U451 ( .A(G113), .ZN(n389) );
  XOR2_X1 U452 ( .A(G140), .B(KEYINPUT12), .Z(n470) );
  XOR2_X1 U453 ( .A(KEYINPUT105), .B(KEYINPUT11), .Z(n472) );
  XOR2_X1 U454 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n446) );
  XNOR2_X1 U455 ( .A(KEYINPUT4), .B(KEYINPUT98), .ZN(n445) );
  XNOR2_X1 U456 ( .A(n475), .B(n361), .ZN(n421) );
  NAND2_X1 U457 ( .A1(n374), .A2(n408), .ZN(n604) );
  AND2_X1 U458 ( .A1(n430), .A2(n649), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n375), .B(n571), .ZN(n374) );
  INV_X1 U460 ( .A(n596), .ZN(n382) );
  INV_X1 U461 ( .A(KEYINPUT34), .ZN(n372) );
  XNOR2_X1 U462 ( .A(G116), .B(G107), .ZN(n483) );
  XNOR2_X1 U463 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U464 ( .A1(n381), .A2(n380), .ZN(n378) );
  AND2_X1 U465 ( .A1(n384), .A2(n383), .ZN(n379) );
  NOR2_X1 U466 ( .A1(n599), .A2(n385), .ZN(n380) );
  XNOR2_X1 U467 ( .A(n514), .B(n399), .ZN(n546) );
  INV_X1 U468 ( .A(KEYINPUT111), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n377), .B(KEYINPUT41), .ZN(n687) );
  NOR2_X1 U470 ( .A1(n676), .A2(n675), .ZN(n377) );
  INV_X1 U471 ( .A(n662), .ZN(n425) );
  NOR2_X1 U472 ( .A1(n530), .A2(n529), .ZN(n426) );
  INV_X1 U473 ( .A(KEYINPUT30), .ZN(n407) );
  OR2_X1 U474 ( .A1(n538), .A2(n583), .ZN(n539) );
  NAND2_X1 U475 ( .A1(n586), .A2(n658), .ZN(n662) );
  XNOR2_X1 U476 ( .A(n466), .B(n465), .ZN(n625) );
  XNOR2_X1 U477 ( .A(n423), .B(n498), .ZN(n707) );
  XNOR2_X1 U478 ( .A(n497), .B(n354), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U480 ( .A1(n397), .A2(n652), .ZN(n608) );
  XOR2_X1 U481 ( .A(KEYINPUT97), .B(n614), .Z(n711) );
  XNOR2_X1 U482 ( .A(n619), .B(KEYINPUT55), .ZN(n620) );
  XNOR2_X1 U483 ( .A(KEYINPUT114), .B(KEYINPUT40), .ZN(n424) );
  INV_X1 U484 ( .A(KEYINPUT35), .ZN(n396) );
  NAND2_X1 U485 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U486 ( .A(n388), .B(KEYINPUT32), .ZN(n741) );
  XNOR2_X1 U487 ( .A(KEYINPUT31), .B(KEYINPUT104), .ZN(n597) );
  XNOR2_X1 U488 ( .A(n387), .B(KEYINPUT110), .ZN(n404) );
  AND2_X1 U489 ( .A1(n412), .A2(n562), .ZN(n644) );
  INV_X1 U490 ( .A(n561), .ZN(n412) );
  AND2_X1 U491 ( .A1(n601), .A2(n358), .ZN(n631) );
  XNOR2_X1 U492 ( .A(KEYINPUT92), .B(n600), .ZN(n601) );
  AND2_X1 U493 ( .A1(n429), .A2(n599), .ZN(n600) );
  XNOR2_X1 U494 ( .A(n516), .B(KEYINPUT100), .ZN(n354) );
  XNOR2_X1 U495 ( .A(n559), .B(KEYINPUT38), .ZN(n355) );
  AND2_X1 U496 ( .A1(n357), .A2(n355), .ZN(n356) );
  AND2_X1 U497 ( .A1(n425), .A2(n426), .ZN(n357) );
  AND2_X1 U498 ( .A1(n659), .A2(n435), .ZN(n358) );
  XOR2_X1 U499 ( .A(n503), .B(n502), .Z(n359) );
  AND2_X1 U500 ( .A1(n582), .A2(n658), .ZN(n360) );
  AND2_X1 U501 ( .A1(G224), .A2(n691), .ZN(n361) );
  INV_X1 U502 ( .A(n430), .ZN(n650) );
  XOR2_X1 U503 ( .A(KEYINPUT76), .B(KEYINPUT22), .Z(n362) );
  XNOR2_X1 U504 ( .A(KEYINPUT6), .B(KEYINPUT108), .ZN(n363) );
  XNOR2_X2 U505 ( .A(n364), .B(n415), .ZN(n720) );
  NAND2_X1 U506 ( .A1(n417), .A2(n416), .ZN(n364) );
  AND2_X1 U507 ( .A1(n741), .A2(n404), .ZN(n386) );
  NAND2_X1 U508 ( .A1(n441), .A2(n376), .ZN(n375) );
  NOR2_X1 U509 ( .A1(n687), .A2(n555), .ZN(n543) );
  NAND2_X1 U510 ( .A1(n355), .A2(n673), .ZN(n676) );
  INV_X1 U511 ( .A(n595), .ZN(n381) );
  XNOR2_X2 U512 ( .A(n418), .B(n579), .ZN(n596) );
  NAND2_X1 U513 ( .A1(n595), .A2(n385), .ZN(n384) );
  NAND2_X1 U514 ( .A1(n405), .A2(n386), .ZN(n395) );
  NAND2_X1 U515 ( .A1(n429), .A2(n585), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n429), .A2(n590), .ZN(n388) );
  XNOR2_X1 U517 ( .A(n404), .B(G110), .ZN(G12) );
  INV_X1 U518 ( .A(n645), .ZN(n394) );
  NAND2_X1 U519 ( .A1(n395), .A2(KEYINPUT44), .ZN(n436) );
  NOR2_X1 U520 ( .A1(n395), .A2(KEYINPUT44), .ZN(n591) );
  INV_X1 U521 ( .A(n405), .ZN(n740) );
  INV_X1 U522 ( .A(n603), .ZN(n397) );
  NAND2_X1 U523 ( .A1(n705), .A2(G472), .ZN(n627) );
  AND2_X4 U524 ( .A1(n607), .A2(n608), .ZN(n705) );
  NAND2_X1 U525 ( .A1(n705), .A2(G210), .ZN(n621) );
  NAND2_X1 U526 ( .A1(n398), .A2(n639), .ZN(n564) );
  NAND2_X1 U527 ( .A1(n557), .A2(KEYINPUT47), .ZN(n398) );
  XNOR2_X2 U528 ( .A(n467), .B(G472), .ZN(n583) );
  AND2_X2 U529 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X2 U530 ( .A1(n663), .A2(n662), .ZN(n580) );
  XNOR2_X2 U531 ( .A(n580), .B(KEYINPUT79), .ZN(n595) );
  BUF_X1 U532 ( .A(n577), .Z(n400) );
  XNOR2_X2 U533 ( .A(n403), .B(n362), .ZN(n429) );
  NAND2_X1 U534 ( .A1(n596), .A2(n360), .ZN(n403) );
  XNOR2_X1 U535 ( .A(n535), .B(n407), .ZN(n406) );
  NAND2_X1 U536 ( .A1(n406), .A2(n357), .ZN(n558) );
  XNOR2_X2 U537 ( .A(n482), .B(n456), .ZN(n460) );
  XNOR2_X2 U538 ( .A(n455), .B(n454), .ZN(n482) );
  XNOR2_X2 U539 ( .A(n444), .B(G143), .ZN(n455) );
  XNOR2_X2 U540 ( .A(n460), .B(n516), .ZN(n725) );
  INV_X1 U541 ( .A(n606), .ZN(n653) );
  INV_X1 U542 ( .A(n720), .ZN(n410) );
  XNOR2_X1 U543 ( .A(n432), .B(KEYINPUT93), .ZN(n416) );
  XNOR2_X1 U544 ( .A(n591), .B(KEYINPUT75), .ZN(n417) );
  XNOR2_X1 U545 ( .A(n455), .B(n421), .ZN(n448) );
  XNOR2_X1 U546 ( .A(n460), .B(n459), .ZN(n466) );
  NOR2_X1 U547 ( .A1(n530), .A2(n662), .ZN(n593) );
  NAND2_X1 U548 ( .A1(n431), .A2(n673), .ZN(n554) );
  OR2_X1 U549 ( .A1(n528), .A2(n431), .ZN(n430) );
  XNOR2_X1 U550 ( .A(n533), .B(n531), .ZN(n431) );
  NAND2_X1 U551 ( .A1(n436), .A2(n433), .ZN(n432) );
  INV_X1 U552 ( .A(n602), .ZN(n435) );
  XNOR2_X2 U553 ( .A(G128), .B(KEYINPUT85), .ZN(n444) );
  AND2_X1 U554 ( .A1(n652), .A2(n720), .ZN(n440) );
  AND2_X1 U555 ( .A1(n569), .A2(n568), .ZN(n441) );
  XNOR2_X1 U556 ( .A(n544), .B(KEYINPUT46), .ZN(n545) );
  INV_X1 U557 ( .A(KEYINPUT48), .ZN(n571) );
  XNOR2_X1 U558 ( .A(n452), .B(KEYINPUT4), .ZN(n453) );
  XNOR2_X1 U559 ( .A(n458), .B(G146), .ZN(n459) );
  XNOR2_X1 U560 ( .A(n476), .B(n453), .ZN(n456) );
  XNOR2_X1 U561 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U562 ( .A(KEYINPUT95), .ZN(n578) );
  XNOR2_X1 U563 ( .A(KEYINPUT16), .B(G122), .ZN(n443) );
  INV_X1 U564 ( .A(n531), .ZN(n532) );
  XNOR2_X1 U565 ( .A(n578), .B(KEYINPUT0), .ZN(n579) );
  XNOR2_X1 U566 ( .A(n549), .B(KEYINPUT94), .ZN(n550) );
  XNOR2_X1 U567 ( .A(n707), .B(n706), .ZN(n708) );
  AND2_X1 U568 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X2 U569 ( .A1(n555), .A2(n400), .ZN(n640) );
  XNOR2_X1 U570 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U571 ( .A(KEYINPUT15), .B(G902), .ZN(n499) );
  INV_X1 U572 ( .A(n499), .ZN(n605) );
  XOR2_X1 U573 ( .A(KEYINPUT66), .B(G101), .Z(n457) );
  XNOR2_X1 U574 ( .A(n712), .B(n520), .ZN(n450) );
  XNOR2_X1 U575 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U576 ( .A(n448), .B(n447), .Z(n449) );
  XNOR2_X1 U577 ( .A(n450), .B(n449), .ZN(n618) );
  NOR2_X2 U578 ( .A1(n605), .A2(n618), .ZN(n533) );
  NOR2_X1 U579 ( .A1(G237), .A2(G902), .ZN(n451) );
  XOR2_X1 U580 ( .A(KEYINPUT80), .B(n451), .Z(n515) );
  NAND2_X1 U581 ( .A1(n515), .A2(G210), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT5), .B(n457), .Z(n458) );
  XOR2_X1 U583 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n462) );
  NAND2_X1 U584 ( .A1(n468), .A2(G210), .ZN(n461) );
  XNOR2_X1 U585 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U586 ( .A1(n625), .A2(G902), .ZN(n467) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(G475), .ZN(n481) );
  NAND2_X1 U588 ( .A1(G214), .A2(n468), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(n469), .ZN(n474) );
  XNOR2_X1 U590 ( .A(G113), .B(G122), .ZN(n471) );
  XNOR2_X1 U591 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U592 ( .A(n474), .B(n473), .Z(n480) );
  XNOR2_X1 U593 ( .A(n476), .B(G143), .ZN(n477) );
  XNOR2_X1 U594 ( .A(n477), .B(G104), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n480), .B(n479), .ZN(n609) );
  XOR2_X1 U596 ( .A(KEYINPUT106), .B(G122), .Z(n484) );
  XNOR2_X1 U597 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n482), .B(n485), .ZN(n489) );
  XOR2_X1 U599 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n487) );
  NAND2_X1 U600 ( .A1(G217), .A2(n496), .ZN(n486) );
  XNOR2_X1 U601 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U602 ( .A(n489), .B(n488), .ZN(n703) );
  NOR2_X1 U603 ( .A1(G902), .A2(n703), .ZN(n490) );
  XNOR2_X1 U604 ( .A(G478), .B(n490), .ZN(n561) );
  NAND2_X1 U605 ( .A1(n556), .A2(n561), .ZN(n536) );
  XOR2_X1 U606 ( .A(G110), .B(G137), .Z(n492) );
  XNOR2_X1 U607 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U608 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n726), .B(n495), .ZN(n498) );
  NAND2_X1 U610 ( .A1(G221), .A2(n496), .ZN(n497) );
  XOR2_X1 U611 ( .A(KEYINPUT20), .B(KEYINPUT101), .Z(n501) );
  NAND2_X1 U612 ( .A1(G234), .A2(n499), .ZN(n500) );
  XNOR2_X1 U613 ( .A(n501), .B(n500), .ZN(n510) );
  NAND2_X1 U614 ( .A1(n510), .A2(G217), .ZN(n503) );
  XNOR2_X1 U615 ( .A(KEYINPUT82), .B(KEYINPUT25), .ZN(n502) );
  NOR2_X1 U616 ( .A1(G900), .A2(n691), .ZN(n504) );
  NAND2_X1 U617 ( .A1(n504), .A2(G902), .ZN(n505) );
  NAND2_X1 U618 ( .A1(G952), .A2(n691), .ZN(n573) );
  NAND2_X1 U619 ( .A1(n505), .A2(n573), .ZN(n509) );
  XOR2_X1 U620 ( .A(KEYINPUT99), .B(KEYINPUT14), .Z(n507) );
  XNOR2_X1 U621 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U622 ( .A(KEYINPUT78), .B(n508), .ZN(n657) );
  NAND2_X1 U623 ( .A1(n509), .A2(n657), .ZN(n529) );
  NAND2_X1 U624 ( .A1(G221), .A2(n510), .ZN(n511) );
  XOR2_X1 U625 ( .A(KEYINPUT21), .B(n511), .Z(n658) );
  NAND2_X1 U626 ( .A1(n512), .A2(n658), .ZN(n538) );
  NOR2_X1 U627 ( .A1(n536), .A2(n538), .ZN(n513) );
  NAND2_X1 U628 ( .A1(n587), .A2(n513), .ZN(n514) );
  NAND2_X1 U629 ( .A1(n515), .A2(G214), .ZN(n673) );
  NAND2_X1 U630 ( .A1(G227), .A2(n691), .ZN(n517) );
  XNOR2_X1 U631 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U632 ( .A(G469), .B(KEYINPUT71), .ZN(n522) );
  XNOR2_X1 U633 ( .A(n522), .B(KEYINPUT70), .ZN(n523) );
  XNOR2_X2 U634 ( .A(n524), .B(n523), .ZN(n541) );
  NAND2_X1 U635 ( .A1(n673), .A2(n435), .ZN(n526) );
  NOR2_X1 U636 ( .A1(n546), .A2(n526), .ZN(n527) );
  XNOR2_X1 U637 ( .A(n527), .B(KEYINPUT43), .ZN(n528) );
  INV_X1 U638 ( .A(n541), .ZN(n530) );
  XNOR2_X1 U639 ( .A(n533), .B(n532), .ZN(n559) );
  INV_X1 U640 ( .A(n583), .ZN(n534) );
  NAND2_X1 U641 ( .A1(n534), .A2(n673), .ZN(n535) );
  INV_X1 U642 ( .A(n536), .ZN(n642) );
  AND2_X1 U643 ( .A1(n572), .A2(n642), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n539), .B(KEYINPUT28), .ZN(n540) );
  XNOR2_X1 U645 ( .A(n540), .B(KEYINPUT113), .ZN(n542) );
  NAND2_X1 U646 ( .A1(n542), .A2(n541), .ZN(n555) );
  NAND2_X1 U647 ( .A1(n562), .A2(n561), .ZN(n675) );
  XNOR2_X1 U648 ( .A(n543), .B(KEYINPUT42), .ZN(n737) );
  XNOR2_X1 U649 ( .A(KEYINPUT91), .B(KEYINPUT64), .ZN(n544) );
  INV_X1 U650 ( .A(KEYINPUT115), .ZN(n547) );
  XNOR2_X1 U651 ( .A(n547), .B(n546), .ZN(n548) );
  NOR2_X1 U652 ( .A1(n548), .A2(n554), .ZN(n551) );
  INV_X1 U653 ( .A(KEYINPUT36), .ZN(n549) );
  XNOR2_X1 U654 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U655 ( .A1(n552), .A2(n435), .ZN(n647) );
  XNOR2_X1 U656 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n553) );
  NOR2_X1 U657 ( .A1(n642), .A2(n644), .ZN(n677) );
  INV_X1 U658 ( .A(n677), .ZN(n565) );
  NAND2_X1 U659 ( .A1(n640), .A2(n565), .ZN(n557) );
  NOR2_X1 U660 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U661 ( .A(KEYINPUT112), .B(n560), .ZN(n563) );
  NAND2_X1 U662 ( .A1(n563), .A2(n581), .ZN(n639) );
  XOR2_X1 U663 ( .A(KEYINPUT86), .B(n564), .Z(n569) );
  XOR2_X1 U664 ( .A(n565), .B(KEYINPUT87), .Z(n592) );
  NAND2_X1 U665 ( .A1(n640), .A2(n592), .ZN(n566) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(n566), .ZN(n567) );
  XNOR2_X1 U667 ( .A(n567), .B(KEYINPUT77), .ZN(n568) );
  NAND2_X1 U668 ( .A1(n572), .A2(n644), .ZN(n649) );
  NOR2_X1 U669 ( .A1(G898), .A2(n691), .ZN(n716) );
  NAND2_X1 U670 ( .A1(G902), .A2(n716), .ZN(n574) );
  NAND2_X1 U671 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U672 ( .A1(n575), .A2(n657), .ZN(n576) );
  INV_X1 U673 ( .A(n587), .ZN(n599) );
  INV_X1 U674 ( .A(n675), .ZN(n582) );
  OR2_X1 U675 ( .A1(n534), .A2(n586), .ZN(n584) );
  INV_X1 U676 ( .A(n663), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n584), .A2(n602), .ZN(n585) );
  XOR2_X1 U678 ( .A(n586), .B(KEYINPUT109), .Z(n659) );
  OR2_X1 U679 ( .A1(n587), .A2(n659), .ZN(n588) );
  NOR2_X1 U680 ( .A1(n435), .A2(n588), .ZN(n589) );
  XNOR2_X1 U681 ( .A(KEYINPUT84), .B(n589), .ZN(n590) );
  NAND2_X1 U682 ( .A1(n593), .A2(n596), .ZN(n594) );
  NOR2_X1 U683 ( .A1(n595), .A2(n583), .ZN(n669) );
  NAND2_X1 U684 ( .A1(n596), .A2(n669), .ZN(n598) );
  NOR2_X1 U685 ( .A1(n730), .A2(n720), .ZN(n603) );
  NAND2_X1 U686 ( .A1(n705), .A2(G475), .ZN(n613) );
  XOR2_X1 U687 ( .A(n609), .B(KEYINPUT96), .Z(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n610) );
  XNOR2_X1 U689 ( .A(n613), .B(n612), .ZN(n615) );
  NOR2_X1 U690 ( .A1(G952), .A2(n691), .ZN(n614) );
  INV_X1 U691 ( .A(n711), .ZN(n628) );
  NAND2_X1 U692 ( .A1(n615), .A2(n628), .ZN(n617) );
  XNOR2_X1 U693 ( .A(KEYINPUT65), .B(KEYINPUT60), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(G60) );
  XNOR2_X1 U695 ( .A(n618), .B(KEYINPUT54), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n622), .A2(n628), .ZN(n624) );
  INV_X1 U698 ( .A(KEYINPUT56), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(G51) );
  XNOR2_X1 U700 ( .A(n627), .B(n626), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U703 ( .A(n631), .B(G101), .Z(G3) );
  NAND2_X1 U704 ( .A1(n633), .A2(n642), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(G104), .ZN(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n635) );
  NAND2_X1 U707 ( .A1(n633), .A2(n644), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(G107), .B(n636), .ZN(G9) );
  XOR2_X1 U710 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U711 ( .A1(n640), .A2(n644), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U713 ( .A(G143), .B(n639), .ZN(G45) );
  NAND2_X1 U714 ( .A1(n640), .A2(n642), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(G146), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n642), .A2(n353), .ZN(n643) );
  XNOR2_X1 U717 ( .A(G113), .B(n643), .ZN(G15) );
  NAND2_X1 U718 ( .A1(n353), .A2(n644), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n646), .B(G116), .ZN(G18) );
  XNOR2_X1 U720 ( .A(G125), .B(n647), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U722 ( .A(G134), .B(n649), .ZN(G36) );
  XOR2_X1 U723 ( .A(G140), .B(n650), .Z(G42) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n730), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT88), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT89), .ZN(n694) );
  NAND2_X1 U728 ( .A1(G952), .A2(n657), .ZN(n686) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U730 ( .A(n660), .B(KEYINPUT49), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n583), .A2(n661), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n435), .A2(n662), .ZN(n664) );
  XOR2_X1 U733 ( .A(KEYINPUT50), .B(n664), .Z(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT116), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT117), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n687), .A2(n672), .ZN(n683) );
  NOR2_X1 U740 ( .A1(n355), .A2(n673), .ZN(n674) );
  NOR2_X1 U741 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(KEYINPUT118), .ZN(n679) );
  NOR2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U745 ( .A1(n681), .A2(n688), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U749 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n695), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n696), .B(KEYINPUT57), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U755 ( .A1(n705), .A2(G469), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n711), .A2(n701), .ZN(G54) );
  NAND2_X1 U758 ( .A1(G478), .A2(n705), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n711), .A2(n704), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n705), .A2(G217), .ZN(n709) );
  XOR2_X1 U762 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n706) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(G66) );
  XOR2_X1 U764 ( .A(KEYINPUT123), .B(n712), .Z(n715) );
  XNOR2_X1 U765 ( .A(G101), .B(n713), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n717) );
  NOR2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n724) );
  NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n718) );
  XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U770 ( .A1(n719), .A2(G898), .ZN(n722) );
  OR2_X1 U771 ( .A1(n720), .A2(G953), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(G69) );
  XOR2_X1 U774 ( .A(n725), .B(n726), .Z(n731) );
  XNOR2_X1 U775 ( .A(G227), .B(n731), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U777 ( .A1(G953), .A2(n728), .ZN(n729) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(n729), .Z(n735) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n732), .B(KEYINPUT124), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(n691), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n735), .A2(n734), .ZN(G72) );
  XOR2_X1 U783 ( .A(G137), .B(KEYINPUT126), .Z(n736) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(G39) );
  XNOR2_X1 U785 ( .A(n738), .B(G131), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n739), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U787 ( .A(n740), .B(G122), .Z(G24) );
  XNOR2_X1 U788 ( .A(G119), .B(n741), .ZN(G21) );
endmodule

