//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  AND2_X1   g0017(.A1(KEYINPUT65), .A2(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(KEYINPUT65), .A2(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n210), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n212), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT0), .Z(new_n234));
  NOR3_X1   g0034(.A1(new_n227), .A2(new_n231), .A3(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  INV_X1    g0038(.A(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G107), .ZN(new_n248));
  INV_X1    g0048(.A(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n251), .B(new_n255), .Z(G351));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT79), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n257), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(new_n210), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT7), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT7), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n262), .A2(new_n266), .A3(new_n210), .A4(new_n263), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G68), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G159), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT73), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(new_n210), .A3(new_n257), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT73), .B1(G20), .B2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n220), .A2(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n228), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n275), .B2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n268), .A2(KEYINPUT16), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT16), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n266), .A2(KEYINPUT80), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n258), .A2(new_n260), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n283), .A2(KEYINPUT80), .A3(new_n266), .A4(new_n210), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n282), .A2(new_n220), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n273), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n201), .B1(new_n220), .B2(G58), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n210), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n278), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n230), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n277), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT8), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n293), .B1(new_n294), .B2(G58), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT8), .B(G58), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT72), .B(new_n295), .C1(new_n296), .C2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(G58), .ZN(new_n298));
  OR4_X1    g0098(.A1(new_n293), .A2(new_n298), .A3(KEYINPUT72), .A4(KEYINPUT8), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n209), .B2(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n305), .B2(new_n300), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT70), .ZN(new_n308));
  OR2_X1    g0108(.A1(KEYINPUT69), .A2(G45), .ZN(new_n309));
  NAND2_X1  g0109(.A1(KEYINPUT69), .A2(G45), .ZN(new_n310));
  AOI21_X1  g0110(.A(G41), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(G1), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT69), .A2(G45), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT69), .A2(G45), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(KEYINPUT70), .B(new_n313), .C1(new_n318), .C2(G41), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G41), .ZN(new_n321));
  OAI211_X1 g0121(.A(G1), .B(G13), .C1(new_n257), .C2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G232), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n257), .A2(new_n216), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G223), .A2(G1698), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n262), .B2(new_n263), .ZN(new_n328));
  INV_X1    g0128(.A(G1698), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(G226), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n326), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n320), .B(new_n325), .C1(new_n332), .C2(new_n322), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G200), .ZN(new_n334));
  INV_X1    g0134(.A(new_n322), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n330), .B(new_n327), .C1(new_n262), .C2(new_n263), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n326), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(G190), .A3(new_n320), .A4(new_n325), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n292), .A2(new_n307), .A3(new_n334), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n292), .A2(new_n307), .ZN(new_n342));
  INV_X1    g0142(.A(G169), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT81), .ZN(new_n345));
  INV_X1    g0145(.A(G179), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n337), .A2(new_n346), .A3(new_n320), .A4(new_n325), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(new_n344), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n342), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g0152(.A(KEYINPUT18), .B(new_n342), .C1(new_n348), .C2(new_n349), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n341), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n203), .A2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n271), .A2(new_n272), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n257), .A2(G20), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n355), .B1(new_n356), .B2(new_n357), .C1(new_n300), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n291), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n302), .A2(new_n202), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n304), .A2(G50), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n324), .A2(G226), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n281), .A2(G222), .A3(new_n329), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n254), .B2(new_n281), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n283), .A2(new_n329), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(G223), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n320), .B(new_n367), .C1(new_n371), .C2(new_n322), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n361), .A2(KEYINPUT9), .A3(new_n362), .A4(new_n363), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n372), .B2(G200), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n366), .A2(new_n374), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT10), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n372), .A2(G179), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n372), .A2(new_n343), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n364), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n301), .B(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n254), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n304), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n210), .A2(new_n254), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n357), .A2(new_n296), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT15), .B(G87), .Z(new_n389));
  AOI211_X1 g0189(.A(new_n387), .B(new_n388), .C1(new_n358), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n291), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n384), .B1(new_n254), .B2(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n281), .A2(G232), .A3(new_n329), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n281), .A2(G1698), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n393), .B1(new_n206), .B2(new_n281), .C1(new_n394), .C2(new_n222), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n335), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n324), .A2(G244), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n320), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n398), .A2(G179), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n343), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AND4_X1   g0201(.A1(new_n354), .A2(new_n379), .A3(new_n382), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n271), .A2(new_n272), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(G50), .B1(G77), .B2(new_n358), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n221), .A2(G20), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n391), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT11), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n302), .A2(KEYINPUT12), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n383), .A2(KEYINPUT12), .A3(new_n221), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n386), .A2(KEYINPUT12), .ZN(new_n410));
  INV_X1    g0210(.A(G68), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n258), .A2(new_n260), .A3(G226), .A4(new_n329), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n258), .A2(new_n260), .A3(G232), .A4(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n335), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n324), .A2(G238), .ZN(new_n420));
  AND4_X1   g0220(.A1(new_n414), .A2(new_n320), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n315), .A2(new_n319), .B1(new_n324), .B2(G238), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n414), .B1(new_n422), .B2(new_n419), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G190), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n421), .B2(new_n423), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n413), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n392), .B1(G200), .B2(new_n398), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n398), .A2(new_n373), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n421), .B2(new_n423), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(G169), .C1(new_n421), .C2(new_n423), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(KEYINPUT14), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT77), .ZN(new_n437));
  INV_X1    g0237(.A(new_n432), .ZN(new_n438));
  XOR2_X1   g0238(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n439));
  AOI22_X1  g0239(.A1(new_n438), .A2(new_n439), .B1(G179), .B2(new_n424), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n433), .A2(new_n441), .A3(KEYINPUT14), .A4(new_n435), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n413), .ZN(new_n444));
  AOI211_X1 g0244(.A(new_n428), .B(new_n431), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n402), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n262), .A2(new_n263), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n329), .A2(G264), .ZN(new_n449));
  INV_X1    g0249(.A(G257), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n329), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n283), .A2(G303), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n335), .ZN(new_n455));
  INV_X1    g0255(.A(G45), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G1), .ZN(new_n457));
  AND2_X1   g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NOR2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n460), .A2(new_n312), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n322), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G270), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n249), .A2(G20), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n466), .A2(new_n291), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n291), .A4(new_n467), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n470), .A2(new_n471), .B1(new_n383), .B2(new_n249), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n301), .B(new_n385), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n257), .B2(G1), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n209), .A2(KEYINPUT82), .A3(G33), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n291), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(G116), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n343), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n464), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n455), .A2(new_n461), .A3(new_n463), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n472), .A2(new_n478), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(G179), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n464), .A2(KEYINPUT21), .A3(new_n479), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n484), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n464), .A2(new_n373), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(G200), .B2(new_n464), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n473), .A2(new_n389), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n477), .A2(new_n301), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n216), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n448), .A2(new_n210), .A3(G68), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT19), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n210), .B1(new_n417), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(G87), .B2(new_n207), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n499), .A2(KEYINPUT84), .A3(new_n496), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT84), .B1(new_n499), .B2(new_n496), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n495), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n492), .B(new_n494), .C1(new_n503), .C2(new_n291), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n322), .B(G250), .C1(G1), .C2(new_n456), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n457), .A2(G274), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n257), .A2(new_n249), .ZN(new_n507));
  INV_X1    g0307(.A(G244), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n262), .A2(new_n263), .B1(new_n508), .B2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n222), .A2(new_n329), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n505), .B(new_n506), .C1(new_n511), .C2(new_n322), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G200), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(G1698), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n448), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n335), .B1(new_n515), .B2(new_n507), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(G190), .A3(new_n505), .A4(new_n506), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n504), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n492), .B1(new_n503), .B2(new_n291), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n477), .A2(new_n301), .A3(new_n389), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n512), .A2(new_n343), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n516), .A2(new_n346), .A3(new_n505), .A4(new_n506), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n462), .A2(G257), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n370), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .A4(new_n329), .ZN(new_n529));
  AOI211_X1 g0329(.A(new_n508), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n529), .C1(new_n530), .C2(KEYINPUT4), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n335), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n346), .A3(new_n461), .ZN(new_n533));
  AOI21_X1  g0333(.A(G1698), .B1(new_n262), .B2(new_n263), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT4), .B1(new_n534), .B2(G244), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n529), .B(new_n465), .C1(new_n394), .C2(new_n217), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n335), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n461), .A3(new_n526), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n343), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n282), .A2(new_n284), .A3(G107), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n403), .A2(G77), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n542), .A2(new_n205), .A3(G107), .ZN(new_n543));
  XNOR2_X1  g0343(.A(G97), .B(G107), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n540), .B(new_n541), .C1(new_n210), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n291), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n302), .A2(new_n205), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n477), .A2(G97), .A3(new_n301), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n533), .A2(new_n539), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT83), .B1(new_n538), .B2(new_n373), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n532), .A2(new_n553), .A3(G190), .A4(new_n461), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n538), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n525), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n493), .A2(new_n206), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n281), .A2(new_n210), .A3(G87), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n210), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n560), .A2(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n448), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n358), .A2(G116), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .A4(new_n567), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n559), .B1(new_n572), .B2(new_n291), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n301), .A2(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT25), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n450), .A2(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n217), .A2(new_n329), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n448), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n257), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n322), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n460), .A2(G264), .A3(new_n322), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n461), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G169), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT85), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n460), .A2(KEYINPUT85), .A3(G264), .A4(new_n322), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n461), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n582), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G179), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n573), .A2(new_n575), .B1(new_n586), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n573), .A2(new_n575), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n585), .A2(G190), .B1(new_n592), .B2(G200), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n447), .A2(new_n491), .A3(new_n558), .A4(new_n598), .ZN(new_n599));
  XOR2_X1   g0399(.A(new_n599), .B(KEYINPUT86), .Z(G372));
  NAND3_X1  g0400(.A1(new_n573), .A2(new_n597), .A3(new_n575), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n594), .B2(new_n487), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n525), .A2(new_n557), .A3(new_n551), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n524), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n551), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT26), .B1(new_n525), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n518), .A2(new_n524), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n607), .A2(new_n551), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n447), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n382), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n352), .A2(new_n353), .ZN(new_n614));
  INV_X1    g0414(.A(new_n401), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n443), .B2(new_n444), .ZN(new_n616));
  XNOR2_X1  g0416(.A(new_n339), .B(KEYINPUT17), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n427), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n613), .B1(new_n619), .B2(new_n379), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n612), .A2(new_n620), .ZN(G369));
  INV_X1    g0421(.A(G330), .ZN(new_n622));
  INV_X1    g0422(.A(G13), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(G20), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT27), .B1(new_n625), .B2(G1), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT27), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n627), .A3(new_n209), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(G213), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT87), .ZN(new_n630));
  XNOR2_X1  g0430(.A(KEYINPUT88), .B(G343), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n632), .B(KEYINPUT89), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n484), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n491), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n484), .A3(new_n487), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n622), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n594), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(new_n601), .C1(new_n596), .C2(new_n633), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n487), .A2(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n634), .A2(new_n594), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n598), .A2(new_n487), .A3(new_n633), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n638), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  OR3_X1    g0445(.A1(new_n602), .A2(KEYINPUT90), .A3(new_n634), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n602), .B2(new_n634), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(G399));
  NAND2_X1  g0449(.A1(new_n232), .A2(new_n321), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G1), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n229), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT28), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n633), .B1(new_n604), .B2(new_n610), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT29), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g0457(.A(KEYINPUT29), .B(new_n633), .C1(new_n604), .C2(new_n610), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n558), .A2(new_n598), .A3(new_n491), .A4(new_n633), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT30), .ZN(new_n661));
  INV_X1    g0461(.A(new_n512), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n483), .A2(new_n662), .A3(G179), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n532), .A2(new_n592), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n464), .A2(new_n346), .A3(new_n512), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(KEYINPUT30), .A3(new_n532), .A4(new_n592), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n582), .A2(new_n590), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n668), .B(new_n461), .C1(new_n532), .C2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n464), .A3(new_n512), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n461), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n538), .A3(KEYINPUT91), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n346), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n665), .B(new_n667), .C1(new_n671), .C2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT31), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n675), .A2(new_n676), .A3(new_n634), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n675), .B2(new_n634), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n660), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n659), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n654), .B1(new_n681), .B2(G1), .ZN(G364));
  INV_X1    g0482(.A(new_n650), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n209), .B1(new_n624), .B2(G45), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n346), .A2(G200), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n210), .A2(G190), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n690), .A2(KEYINPUT94), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(KEYINPUT94), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n210), .A2(new_n373), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n688), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n694), .A2(G77), .B1(G58), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n210), .A2(new_n346), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G200), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n373), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n698), .B1(new_n202), .B2(new_n702), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT95), .Z(new_n704));
  NOR2_X1   g0504(.A1(G179), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n689), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n706), .A2(KEYINPUT32), .A3(new_n269), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT32), .B1(new_n706), .B2(new_n269), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n346), .A2(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n695), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n216), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n689), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n283), .B(new_n711), .C1(G107), .C2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n708), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n707), .B(new_n716), .C1(new_n715), .C2(new_n714), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n210), .B1(new_n705), .B2(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G97), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n700), .A2(G190), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n722), .B2(new_n411), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n704), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n718), .A2(new_n579), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n281), .B1(new_n701), .B2(G326), .ZN(new_n727));
  INV_X1    g0527(.A(G322), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(new_n696), .ZN(new_n729));
  XNOR2_X1  g0529(.A(KEYINPUT33), .B(G317), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n726), .B(new_n729), .C1(new_n721), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G283), .ZN(new_n732));
  INV_X1    g0532(.A(G329), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n712), .A2(new_n732), .B1(new_n706), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n694), .B2(G311), .ZN(new_n735));
  INV_X1    g0535(.A(G303), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n731), .B(new_n735), .C1(new_n736), .C2(new_n710), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT98), .Z(new_n739));
  OAI211_X1 g0539(.A(G1), .B(G13), .C1(new_n210), .C2(G169), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n687), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n448), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n232), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n229), .B2(new_n318), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n255), .A2(new_n456), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n751), .A2(new_n752), .B1(G116), .B2(new_n232), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n232), .A2(new_n281), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(G87), .B2(new_n207), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n747), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n636), .A2(new_n637), .ZN(new_n757));
  INV_X1    g0557(.A(new_n746), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n743), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n638), .A2(new_n686), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(G330), .B2(new_n757), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(G396));
  NOR2_X1   g0562(.A1(new_n742), .A2(new_n744), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n687), .B1(new_n763), .B2(new_n254), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G137), .A2(new_n701), .B1(new_n721), .B2(G150), .ZN(new_n766));
  INV_X1    g0566(.A(G143), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n766), .B1(new_n767), .B2(new_n696), .C1(new_n269), .C2(new_n693), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT102), .Z(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT34), .ZN(new_n770));
  INV_X1    g0570(.A(G132), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n710), .A2(new_n202), .B1(new_n706), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n748), .B(new_n772), .C1(G58), .C2(new_n719), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n770), .B(new_n773), .C1(new_n411), .C2(new_n712), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n696), .A2(new_n579), .B1(new_n706), .B2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n720), .B1(new_n702), .B2(new_n736), .C1(new_n732), .C2(new_n722), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(G116), .C2(new_n694), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n283), .B1(new_n710), .B2(new_n206), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT100), .Z(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(new_n216), .C2(new_n712), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT101), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n765), .B1(new_n783), .B2(new_n742), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT103), .Z(new_n785));
  OR2_X1    g0585(.A1(new_n401), .A2(KEYINPUT104), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n401), .A2(KEYINPUT104), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n431), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n634), .A2(new_n392), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n615), .A2(new_n634), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n785), .B1(new_n745), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(new_n611), .B2(new_n633), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n431), .B1(new_n787), .B2(new_n786), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n796), .B(new_n633), .C1(new_n604), .C2(new_n610), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OR3_X1    g0598(.A1(new_n795), .A2(new_n680), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n680), .B1(new_n795), .B2(new_n798), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n687), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n794), .A2(new_n801), .ZN(G384));
  INV_X1    g0602(.A(KEYINPUT109), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n443), .A2(new_n444), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n634), .A2(new_n444), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n427), .A3(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n444), .B(new_n634), .C1(new_n443), .C2(new_n428), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n808), .A2(KEYINPUT40), .A3(new_n679), .A4(new_n793), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT37), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n411), .B1(new_n264), .B2(KEYINPUT7), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n288), .B1(new_n267), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n391), .B1(new_n813), .B2(KEYINPUT16), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n306), .B1(new_n814), .B2(new_n289), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n344), .A2(new_n347), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT81), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT105), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND4_X1   g0621(.A1(new_n292), .A2(new_n307), .A3(new_n338), .A4(new_n334), .ZN(new_n822));
  INV_X1    g0622(.A(new_n630), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n292), .B2(new_n307), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n820), .B(new_n342), .C1(new_n348), .C2(new_n349), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT107), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n339), .B1(new_n815), .B2(new_n823), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT37), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n819), .B2(new_n820), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT37), .B1(new_n350), .B2(KEYINPUT105), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT107), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n828), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n614), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n824), .B1(new_n836), .B2(new_n341), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n268), .A2(new_n276), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n278), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n306), .B1(new_n814), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(new_n817), .B2(new_n818), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n339), .B1(new_n843), .B2(new_n823), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT37), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n821), .B2(new_n827), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n277), .A2(new_n291), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n813), .A2(KEYINPUT16), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n307), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n630), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n847), .B(KEYINPUT38), .C1(new_n354), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n803), .B1(new_n810), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n839), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n835), .B2(new_n837), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n851), .B1(new_n614), .B2(new_n617), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n850), .B1(new_n348), .B2(new_n349), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n339), .A3(new_n851), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n831), .A2(new_n832), .B1(new_n859), .B2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n857), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n863), .A2(new_n809), .A3(KEYINPUT109), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n861), .B1(new_n857), .B2(new_n860), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n852), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n808), .A2(new_n679), .A3(new_n793), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n447), .A2(new_n679), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n872), .B(new_n873), .Z(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G330), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n614), .A2(new_n630), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n786), .A2(new_n633), .A3(new_n787), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n797), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n808), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(new_n869), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n840), .A2(KEYINPUT108), .A3(new_n881), .A4(new_n852), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n862), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT108), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n443), .A2(new_n444), .A3(new_n633), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n876), .B(new_n880), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n657), .A2(new_n445), .A3(new_n402), .A4(new_n658), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n620), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n889), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n875), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n209), .B2(new_n624), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT35), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n210), .B(new_n230), .C1(new_n545), .C2(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(G116), .C1(new_n895), .C2(new_n545), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n274), .A2(G50), .A3(G77), .A4(new_n228), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(G50), .B2(new_n411), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n623), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n894), .A2(new_n898), .A3(new_n901), .ZN(G367));
  INV_X1    g0702(.A(new_n710), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(KEYINPUT46), .A3(G116), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT46), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n710), .B2(new_n249), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n904), .B(new_n906), .C1(new_n722), .C2(new_n579), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n748), .B1(new_n702), .B2(new_n775), .ZN(new_n908));
  INV_X1    g0708(.A(G317), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n696), .A2(new_n736), .B1(new_n706), .B2(new_n909), .ZN(new_n910));
  OR3_X1    g0710(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n694), .A2(G283), .B1(G107), .B2(new_n719), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(KEYINPUT111), .B2(new_n913), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n914), .B1(KEYINPUT111), .B2(new_n913), .C1(new_n205), .C2(new_n712), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n281), .B1(new_n722), .B2(new_n269), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n702), .A2(new_n767), .B1(new_n718), .B2(new_n411), .ZN(new_n917));
  INV_X1    g0717(.A(new_n706), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n916), .B(new_n917), .C1(G137), .C2(new_n918), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n712), .A2(new_n254), .B1(new_n696), .B2(new_n356), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n694), .B2(G50), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n919), .B(new_n921), .C1(new_n298), .C2(new_n710), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT47), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n687), .B1(new_n924), .B2(new_n742), .ZN(new_n925));
  INV_X1    g0725(.A(new_n389), .ZN(new_n926));
  INV_X1    g0726(.A(new_n750), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n747), .B1(new_n232), .B2(new_n926), .C1(new_n927), .C2(new_n245), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n633), .A2(new_n504), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n525), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n925), .B(new_n928), .C1(new_n758), .C2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n645), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n638), .B1(new_n643), .B2(new_n644), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n680), .A3(new_n659), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT110), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT45), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n557), .B(new_n551), .C1(new_n555), .C2(new_n633), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n634), .A2(new_n605), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n938), .B(new_n942), .C1(new_n646), .C2(new_n647), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT45), .B1(new_n648), .B2(new_n941), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n646), .A2(new_n647), .A3(new_n942), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT44), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n645), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n946), .A2(new_n947), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n950), .A2(new_n951), .B1(new_n943), .B2(new_n944), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n933), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n681), .B1(new_n937), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n650), .B(KEYINPUT41), .Z(new_n956));
  AOI21_X1  g0756(.A(new_n685), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n942), .A2(new_n644), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n939), .A2(new_n639), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n633), .B1(new_n960), .B2(new_n605), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n645), .A2(new_n942), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n962), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n966), .B2(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n932), .B1(new_n957), .B2(new_n972), .ZN(G387));
  NAND2_X1  g0773(.A1(new_n935), .A2(new_n685), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G311), .A2(new_n721), .B1(new_n701), .B2(G322), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n909), .B2(new_n696), .C1(new_n736), .C2(new_n693), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT48), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n732), .B2(new_n718), .C1(new_n579), .C2(new_n710), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT49), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n918), .A2(G326), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n448), .B1(G116), .B2(new_n713), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n903), .A2(G77), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n712), .B2(new_n205), .C1(new_n696), .C2(new_n202), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n448), .B1(new_n702), .B2(new_n269), .C1(new_n926), .C2(new_n718), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G68), .C2(new_n694), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n356), .B2(new_n706), .C1(new_n300), .C2(new_n722), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n687), .B1(new_n990), .B2(new_n742), .ZN(new_n991));
  INV_X1    g0791(.A(new_n651), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G68), .B2(G77), .ZN(new_n993));
  INV_X1    g0793(.A(new_n296), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n202), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n456), .C1(KEYINPUT50), .C2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(KEYINPUT50), .B2(new_n995), .ZN(new_n997));
  INV_X1    g0797(.A(new_n240), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n927), .B(new_n997), .C1(new_n998), .C2(new_n318), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n754), .A2(new_n651), .B1(G107), .B2(new_n232), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT112), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n747), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n640), .A2(new_n642), .A3(new_n746), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n683), .B1(new_n681), .B2(new_n935), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n936), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n974), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(G393));
  NAND2_X1  g0807(.A1(new_n954), .A2(new_n936), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n683), .C1(new_n937), .C2(new_n954), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n949), .A2(new_n953), .A3(new_n685), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT113), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n747), .B1(new_n205), .B2(new_n232), .C1(new_n927), .C2(new_n250), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n283), .B1(new_n712), .B2(new_n206), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n722), .A2(new_n736), .B1(new_n718), .B2(new_n249), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G322), .C2(new_n918), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n701), .A2(G317), .B1(new_n697), .B2(G311), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT52), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n694), .A2(G294), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n903), .A2(G283), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n701), .A2(G150), .B1(new_n697), .B2(G159), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT51), .Z(new_n1022));
  NOR2_X1   g0822(.A1(new_n718), .A2(new_n254), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1023), .B(new_n748), .C1(G50), .C2(new_n721), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n221), .A2(new_n710), .B1(new_n712), .B2(new_n216), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n694), .B2(new_n994), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n706), .A2(new_n767), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n687), .B1(new_n1029), .B2(new_n742), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1012), .B(new_n1030), .C1(new_n941), .C2(new_n758), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1010), .A2(new_n1011), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1010), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1009), .B1(new_n1032), .B2(new_n1033), .ZN(G390));
  NAND4_X1  g0834(.A1(new_n402), .A2(new_n445), .A3(G330), .A4(new_n679), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n890), .A2(new_n620), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n679), .A2(new_n793), .A3(G330), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n806), .A2(new_n807), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n878), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n808), .A2(G330), .A3(new_n679), .A4(new_n793), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1041), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1037), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n879), .A2(new_n887), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n882), .B(new_n1046), .C1(new_n883), .C2(new_n885), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n853), .A2(new_n887), .A3(new_n879), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n1042), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  OAI211_X1 g0850(.A(KEYINPUT114), .B(new_n1045), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1042), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1047), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1051), .A2(new_n1057), .A3(new_n683), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n685), .A3(new_n1056), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n722), .A2(new_n206), .B1(new_n702), .B2(new_n732), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1060), .A2(new_n281), .A3(new_n711), .A4(new_n1023), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n712), .A2(new_n411), .B1(new_n706), .B2(new_n579), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n694), .B2(G97), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n249), .C2(new_n696), .ZN(new_n1064));
  INV_X1    g0864(.A(G137), .ZN(new_n1065));
  INV_X1    g0865(.A(G128), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n722), .A2(new_n1065), .B1(new_n702), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G159), .B2(new_n719), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n694), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n710), .A2(new_n356), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT53), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n281), .B1(new_n712), .B2(new_n202), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G132), .B2(new_n697), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(G125), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n706), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1064), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(new_n742), .B1(new_n300), .B2(new_n763), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n686), .B(new_n1079), .C1(new_n886), .C2(new_n745), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1058), .A2(new_n1059), .A3(new_n1080), .ZN(G378));
  AOI22_X1  g0881(.A1(new_n701), .A2(G125), .B1(G150), .B2(new_n719), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT119), .Z(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G128), .B2(new_n697), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n903), .A2(new_n1069), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT118), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n693), .A2(new_n1065), .B1(new_n771), .B2(new_n722), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT117), .Z(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT59), .Z(new_n1090));
  AOI21_X1  g0890(.A(G41), .B1(new_n918), .B2(G124), .ZN(new_n1091));
  AOI21_X1  g0891(.A(G33), .B1(new_n713), .B2(G159), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n693), .A2(new_n926), .B1(new_n205), .B2(new_n722), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT115), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G107), .A2(new_n697), .B1(new_n918), .B2(G283), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n748), .C1(new_n298), .C2(new_n712), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n985), .B1(new_n411), .B2(new_n718), .C1(new_n702), .C2(new_n249), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1095), .A2(G41), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(G41), .B1(new_n448), .B2(G33), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1099), .A2(KEYINPUT58), .B1(G50), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT116), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(KEYINPUT58), .B2(new_n1099), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1093), .B(new_n1103), .C1(new_n1102), .C2(new_n1101), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1104), .A2(new_n742), .B1(new_n202), .B2(new_n763), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT56), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n379), .A2(new_n382), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n364), .A2(new_n630), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT55), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n379), .A2(new_n382), .A3(new_n1108), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1111), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1106), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1117), .A2(new_n1113), .A3(KEYINPUT56), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n686), .B(new_n1105), .C1(new_n1119), .C2(new_n745), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(KEYINPUT120), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n880), .B1(new_n886), .B2(new_n888), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n614), .B2(new_n630), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n810), .A2(new_n853), .A3(new_n803), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT109), .B1(new_n863), .B2(new_n809), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(G330), .A4(new_n871), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1125), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n865), .A2(G330), .A3(new_n871), .A4(new_n1119), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n889), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1121), .B(new_n1123), .C1(new_n1136), .C2(new_n685), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1054), .A2(new_n1056), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1037), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(KEYINPUT57), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n683), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1132), .A2(new_n1135), .B1(new_n1140), .B2(new_n1037), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(KEYINPUT57), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1137), .B1(new_n1143), .B2(new_n1145), .ZN(G375));
  NAND2_X1  g0946(.A1(new_n1039), .A2(new_n744), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G159), .A2(new_n903), .B1(new_n713), .B2(G58), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n1066), .B2(new_n706), .C1(new_n1065), .C2(new_n696), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n721), .A2(new_n1069), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n448), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n694), .A2(G150), .B1(G50), .B2(new_n719), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1149), .B(new_n1151), .C1(new_n1153), .C2(KEYINPUT122), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(KEYINPUT122), .B2(new_n1153), .C1(new_n771), .C2(new_n702), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n283), .B1(new_n712), .B2(new_n254), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n722), .A2(new_n249), .B1(new_n702), .B2(new_n579), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n389), .C2(new_n719), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n710), .A2(new_n205), .B1(new_n696), .B2(new_n732), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n694), .B2(G107), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1158), .B(new_n1160), .C1(new_n736), .C2(new_n706), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n741), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n411), .B2(new_n763), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1147), .A2(new_n686), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n1138), .B2(new_n684), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n878), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1040), .A2(new_n1042), .A3(new_n1041), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1036), .A3(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n956), .B(KEYINPUT121), .Z(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1045), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT123), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(G381));
  AND3_X1   g0976(.A1(new_n1133), .A2(new_n889), .A3(new_n1134), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n889), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n685), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1121), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n1122), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(G378), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n650), .B1(new_n1144), .B2(KEYINPUT57), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1188), .A2(G387), .A3(G390), .ZN(new_n1189));
  INV_X1    g0989(.A(G384), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1175), .A4(new_n1191), .ZN(G407));
  INV_X1    g0992(.A(G213), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n631), .A2(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT124), .Z(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(G407), .B(G213), .C1(new_n1188), .C2(new_n1196), .ZN(G409));
  NAND2_X1  g0997(.A1(G375), .A2(G378), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1136), .A2(new_n1141), .A3(new_n1172), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1195), .B1(new_n1182), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n650), .B1(new_n1170), .B2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1168), .A2(new_n1036), .A3(KEYINPUT60), .A4(new_n1169), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(new_n1045), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT125), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1203), .A2(new_n1045), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT125), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1202), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G384), .B1(new_n1209), .B2(new_n1166), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1190), .B(new_n1165), .C1(new_n1205), .C2(new_n1208), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1198), .A2(new_n1200), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT62), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n1058), .A2(new_n1059), .A3(new_n1080), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1123), .B1(new_n1136), .B2(new_n685), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1180), .A4(new_n1199), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1181), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1196), .B(new_n1217), .C1(new_n1218), .C2(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1195), .A2(G2897), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1208), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1207), .B1(new_n1206), .B2(new_n1202), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1166), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1190), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1209), .A2(G384), .A3(new_n1166), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1220), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT61), .B1(new_n1219), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1198), .A2(new_n1200), .A3(new_n1231), .A4(new_n1212), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1214), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G390), .B(new_n932), .C1(new_n957), .C2(new_n972), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1191), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G387), .B(new_n1009), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1234), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT127), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1191), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1244), .A2(new_n1234), .A3(new_n1240), .A4(new_n1238), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1243), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1233), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(new_n1228), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1213), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1215), .B1(new_n1187), .B2(new_n1137), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1217), .A2(new_n1196), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1212), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1253), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1249), .A2(new_n1261), .ZN(G405));
  NAND2_X1  g1062(.A1(new_n1198), .A2(new_n1188), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1212), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1198), .A2(new_n1188), .A3(new_n1257), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1254), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(G402));
endmodule


