

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587;

  XNOR2_X1 U321 ( .A(n367), .B(KEYINPUT115), .ZN(n368) );
  INV_X1 U322 ( .A(KEYINPUT47), .ZN(n367) );
  XNOR2_X1 U323 ( .A(n392), .B(G169GAT), .ZN(n447) );
  XNOR2_X1 U324 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n377) );
  INV_X1 U325 ( .A(G113GAT), .ZN(n446) );
  XOR2_X1 U326 ( .A(KEYINPUT38), .B(n479), .Z(n508) );
  XOR2_X1 U327 ( .A(G29GAT), .B(G43GAT), .Z(n289) );
  XOR2_X1 U328 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n290) );
  XOR2_X1 U329 ( .A(n361), .B(KEYINPUT73), .Z(n291) );
  XOR2_X1 U330 ( .A(KEYINPUT103), .B(n475), .Z(n292) );
  XNOR2_X1 U331 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n471) );
  XNOR2_X1 U332 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U333 ( .A(KEYINPUT9), .ZN(n354) );
  INV_X1 U334 ( .A(KEYINPUT75), .ZN(n314) );
  XNOR2_X1 U335 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U336 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U337 ( .A(n369), .B(n368), .ZN(n376) );
  XNOR2_X1 U338 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U339 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U340 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U341 ( .A(n324), .B(n323), .ZN(n325) );
  NOR2_X1 U342 ( .A1(n420), .A2(n547), .ZN(n572) );
  XNOR2_X1 U343 ( .A(n326), .B(n325), .ZN(n370) );
  XNOR2_X1 U344 ( .A(n455), .B(n454), .ZN(n534) );
  XOR2_X1 U345 ( .A(n419), .B(n418), .Z(n547) );
  XNOR2_X1 U346 ( .A(n483), .B(G190GAT), .ZN(n484) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U348 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(G22GAT), .B(G197GAT), .Z(n294) );
  XNOR2_X1 U351 ( .A(G36GAT), .B(G50GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U353 ( .A(n295), .B(G141GAT), .Z(n297) );
  XOR2_X1 U354 ( .A(G113GAT), .B(G1GAT), .Z(n411) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(n411), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n302) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n289), .B(n298), .ZN(n357) );
  XOR2_X1 U359 ( .A(n357), .B(KEYINPUT66), .Z(n300) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U361 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U362 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U363 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n304) );
  XNOR2_X1 U364 ( .A(G15GAT), .B(KEYINPUT70), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U366 ( .A(G8GAT), .B(KEYINPUT68), .Z(n306) );
  XNOR2_X1 U367 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n305) );
  XNOR2_X1 U368 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(n310), .B(n309), .Z(n552) );
  INV_X1 U371 ( .A(n552), .ZN(n573) );
  XOR2_X1 U372 ( .A(G92GAT), .B(KEYINPUT72), .Z(n312) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G85GAT), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n361) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n291), .B(n313), .ZN(n317) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .Z(n339) );
  XNOR2_X1 U378 ( .A(G204GAT), .B(n339), .ZN(n315) );
  XOR2_X1 U379 ( .A(G176GAT), .B(G64GAT), .Z(n382) );
  XOR2_X1 U380 ( .A(n318), .B(n382), .Z(n326) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G71GAT), .Z(n450) );
  XOR2_X1 U382 ( .A(G78GAT), .B(G148GAT), .Z(n320) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n429) );
  XNOR2_X1 U385 ( .A(n450), .B(n429), .ZN(n324) );
  XOR2_X1 U386 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n322) );
  XNOR2_X1 U387 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n321) );
  XNOR2_X1 U388 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n370), .B(KEYINPUT41), .ZN(n565) );
  NOR2_X1 U390 ( .A1(n565), .A2(n573), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n327), .B(KEYINPUT46), .ZN(n346) );
  XOR2_X1 U392 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U393 ( .A(n428), .B(KEYINPUT83), .Z(n329) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U396 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n331) );
  XNOR2_X1 U397 ( .A(KEYINPUT14), .B(KEYINPUT82), .ZN(n330) );
  XNOR2_X1 U398 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U399 ( .A(n333), .B(n332), .Z(n338) );
  XOR2_X1 U400 ( .A(G15GAT), .B(G127GAT), .Z(n452) );
  XOR2_X1 U401 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n335) );
  XNOR2_X1 U402 ( .A(G1GAT), .B(G64GAT), .ZN(n334) );
  XNOR2_X1 U403 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n452), .B(n336), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U406 ( .A(G8GAT), .B(KEYINPUT80), .Z(n379) );
  XOR2_X1 U407 ( .A(n379), .B(n339), .Z(n341) );
  XNOR2_X1 U408 ( .A(G78GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U410 ( .A(n343), .B(n342), .Z(n345) );
  XNOR2_X1 U411 ( .A(G183GAT), .B(G71GAT), .ZN(n344) );
  XOR2_X1 U412 ( .A(n345), .B(n344), .Z(n559) );
  INV_X1 U413 ( .A(n559), .ZN(n581) );
  NOR2_X1 U414 ( .A1(n346), .A2(n559), .ZN(n366) );
  XOR2_X1 U415 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n348) );
  XNOR2_X1 U416 ( .A(KEYINPUT79), .B(KEYINPUT77), .ZN(n347) );
  XNOR2_X1 U417 ( .A(n348), .B(n347), .ZN(n365) );
  XOR2_X1 U418 ( .A(KEYINPUT65), .B(KEYINPUT78), .Z(n350) );
  XNOR2_X1 U419 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n349) );
  XNOR2_X1 U420 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U421 ( .A(G36GAT), .B(G190GAT), .Z(n388) );
  XOR2_X1 U422 ( .A(n351), .B(n388), .Z(n353) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(G106GAT), .ZN(n352) );
  XNOR2_X1 U424 ( .A(n353), .B(n352), .ZN(n359) );
  NAND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XOR2_X1 U426 ( .A(n359), .B(n358), .Z(n363) );
  XNOR2_X1 U427 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n360), .B(G162GAT), .ZN(n425) );
  XNOR2_X1 U429 ( .A(n425), .B(n361), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n543) );
  INV_X1 U432 ( .A(n543), .ZN(n562) );
  NAND2_X1 U433 ( .A1(n366), .A2(n543), .ZN(n369) );
  XOR2_X1 U434 ( .A(n543), .B(KEYINPUT109), .Z(n371) );
  XNOR2_X1 U435 ( .A(n371), .B(KEYINPUT36), .ZN(n585) );
  NOR2_X1 U436 ( .A1(n581), .A2(n585), .ZN(n372) );
  XNOR2_X1 U437 ( .A(KEYINPUT45), .B(n372), .ZN(n373) );
  NAND2_X1 U438 ( .A1(n373), .A2(n573), .ZN(n374) );
  NOR2_X1 U439 ( .A1(n370), .A2(n374), .ZN(n375) );
  NOR2_X1 U440 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n549) );
  XOR2_X1 U442 ( .A(n379), .B(G92GAT), .Z(n381) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U445 ( .A(n383), .B(n382), .Z(n390) );
  XNOR2_X1 U446 ( .A(G211GAT), .B(G218GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(KEYINPUT21), .ZN(n385) );
  XOR2_X1 U448 ( .A(n385), .B(KEYINPUT90), .Z(n387) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G204GAT), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n423) );
  XNOR2_X1 U451 ( .A(n423), .B(n388), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n394) );
  XNOR2_X1 U453 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n290), .B(n391), .ZN(n392) );
  INV_X1 U455 ( .A(n447), .ZN(n393) );
  XOR2_X1 U456 ( .A(n394), .B(n393), .Z(n462) );
  NOR2_X1 U457 ( .A1(n549), .A2(n462), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT54), .B(n395), .Z(n420) );
  XOR2_X1 U459 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n397) );
  XNOR2_X1 U460 ( .A(KEYINPUT2), .B(KEYINPUT91), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U462 ( .A(G141GAT), .B(n398), .Z(n436) );
  INV_X1 U463 ( .A(n436), .ZN(n419) );
  XOR2_X1 U464 ( .A(KEYINPUT98), .B(KEYINPUT1), .Z(n400) );
  XNOR2_X1 U465 ( .A(G120GAT), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n402) );
  XNOR2_X1 U468 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U470 ( .A(n404), .B(n403), .Z(n417) );
  XNOR2_X1 U471 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n405), .B(KEYINPUT87), .ZN(n453) );
  XOR2_X1 U473 ( .A(KEYINPUT4), .B(n453), .Z(n407) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n415) );
  XOR2_X1 U476 ( .A(G155GAT), .B(G148GAT), .Z(n409) );
  XNOR2_X1 U477 ( .A(G127GAT), .B(G162GAT), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U479 ( .A(n410), .B(G85GAT), .Z(n413) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U484 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n422) );
  XNOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT94), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n435) );
  XOR2_X1 U488 ( .A(n425), .B(KEYINPUT24), .Z(n427) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U491 ( .A(n428), .B(KEYINPUT93), .Z(n431) );
  XNOR2_X1 U492 ( .A(n429), .B(KEYINPUT95), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U496 ( .A(n437), .B(n436), .Z(n469) );
  NAND2_X1 U497 ( .A1(n572), .A2(n469), .ZN(n439) );
  XOR2_X1 U498 ( .A(KEYINPUT55), .B(KEYINPUT123), .Z(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n456) );
  XOR2_X1 U500 ( .A(KEYINPUT88), .B(G176GAT), .Z(n441) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U503 ( .A(KEYINPUT20), .B(G99GAT), .Z(n443) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G190GAT), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U506 ( .A(n445), .B(n444), .Z(n449) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U508 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U510 ( .A1(n456), .A2(n534), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT124), .ZN(n482) );
  NOR2_X1 U512 ( .A1(n573), .A2(n482), .ZN(n459) );
  INV_X1 U513 ( .A(G169GAT), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(G1348GAT) );
  NOR2_X1 U515 ( .A1(n581), .A2(n482), .ZN(n461) );
  INV_X1 U516 ( .A(G183GAT), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(G1350GAT) );
  XOR2_X1 U518 ( .A(n469), .B(KEYINPUT28), .Z(n528) );
  INV_X1 U519 ( .A(n462), .ZN(n525) );
  XNOR2_X1 U520 ( .A(n525), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT27), .B(n463), .ZN(n467) );
  NOR2_X1 U522 ( .A1(n528), .A2(n467), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n547), .ZN(n532) );
  XNOR2_X1 U524 ( .A(KEYINPUT100), .B(n532), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n534), .A2(n465), .ZN(n476) );
  NOR2_X1 U526 ( .A1(n534), .A2(n469), .ZN(n466) );
  XOR2_X1 U527 ( .A(KEYINPUT26), .B(n466), .Z(n570) );
  NOR2_X1 U528 ( .A1(n570), .A2(n467), .ZN(n548) );
  AND2_X1 U529 ( .A1(n525), .A2(n534), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT101), .B(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n470), .A2(n469), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n548), .A2(n473), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n474), .A2(n547), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n476), .A2(n292), .ZN(n490) );
  NOR2_X1 U535 ( .A1(n585), .A2(n490), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n581), .A2(n477), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT37), .B(n478), .ZN(n522) );
  NOR2_X1 U538 ( .A1(n573), .A2(n370), .ZN(n491) );
  NAND2_X1 U539 ( .A1(n522), .A2(n491), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n508), .A2(n534), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n482), .A2(n543), .ZN(n485) );
  INV_X1 U542 ( .A(KEYINPUT58), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n493) );
  XOR2_X1 U544 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n487) );
  NAND2_X1 U545 ( .A1(n559), .A2(n543), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT16), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n511) );
  AND2_X1 U549 ( .A1(n491), .A2(n511), .ZN(n500) );
  NAND2_X1 U550 ( .A1(n500), .A2(n547), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U552 ( .A(G1GAT), .B(n494), .Z(G1324GAT) );
  XOR2_X1 U553 ( .A(G8GAT), .B(KEYINPUT105), .Z(n496) );
  NAND2_X1 U554 ( .A1(n500), .A2(n525), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U557 ( .A1(n500), .A2(n534), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n502) );
  NAND2_X1 U561 ( .A1(n500), .A2(n528), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .Z(n505) );
  NAND2_X1 U565 ( .A1(n508), .A2(n547), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT110), .ZN(n507) );
  NAND2_X1 U568 ( .A1(n525), .A2(n508), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n528), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U572 ( .A1(n552), .A2(n565), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(KEYINPUT112), .ZN(n521) );
  AND2_X1 U574 ( .A1(n511), .A2(n521), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n547), .A2(n518), .ZN(n514) );
  XOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT111), .Z(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT42), .B(n512), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT113), .Z(n516) );
  NAND2_X1 U580 ( .A1(n518), .A2(n525), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n534), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n528), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT114), .ZN(n524) );
  AND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n529), .A2(n547), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n525), .A2(n529), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n534), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n549), .A2(n532), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n573), .A2(n542), .ZN(n535) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n535), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n542), .A2(n565), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n537) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n581), .A2(n542), .ZN(n540) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n540), .Z(n541) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT121), .Z(n554) );
  NAND2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(KEYINPUT120), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n563), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  INV_X1 U621 ( .A(n565), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n563), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT122), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U630 ( .A1(n482), .A2(n565), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT57), .Z(n567) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  INV_X1 U635 ( .A(n570), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n584) );
  NOR2_X1 U637 ( .A1(n573), .A2(n584), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U642 ( .A(n584), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n577), .A2(n370), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

