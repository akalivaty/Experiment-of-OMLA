//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n208), .A2(KEYINPUT23), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n205), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT23), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n213), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n212), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n229), .A2(new_n205), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT67), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(new_n209), .A3(new_n207), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT23), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n219), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT27), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT27), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G183gat), .ZN(new_n242));
  INV_X1    g041(.A(G190gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT28), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n249), .A3(new_n234), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n251), .A2(new_n212), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AND4_X1   g052(.A1(KEYINPUT68), .A2(new_n248), .A3(new_n217), .A4(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n217), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n255), .B1(new_n246), .B2(new_n247), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT68), .B1(new_n256), .B2(new_n253), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n238), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G134gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G127gat), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G134gat), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT70), .B(G113gat), .Z(new_n267));
  OAI211_X1 g066(.A(new_n263), .B(new_n266), .C1(new_n267), .C2(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n264), .A2(new_n265), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NAND2_X1  g069(.A1(G113gat), .A2(G120gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n260), .A2(new_n262), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n272), .B2(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n268), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n268), .B(KEYINPUT71), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n258), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT27), .B(G183gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT28), .B1(new_n283), .B2(new_n243), .ZN(new_n284));
  INV_X1    g083(.A(new_n247), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n253), .B(new_n217), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n256), .A2(KEYINPUT68), .A3(new_n253), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(new_n238), .B1(new_n279), .B2(new_n280), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n204), .B1(new_n282), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G71gat), .B(G99gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n293), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n258), .A2(new_n281), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n290), .A2(new_n279), .A3(new_n280), .A4(new_n238), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n300), .B1(new_n303), .B2(new_n204), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(KEYINPUT33), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT72), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n204), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(new_n301), .B2(new_n302), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n309));
  INV_X1    g108(.A(new_n305), .ZN(new_n310));
  NOR4_X1   g109(.A1(new_n308), .A2(new_n309), .A3(new_n300), .A4(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n299), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(new_n302), .A3(new_n307), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n313), .B(KEYINPUT34), .Z(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n314), .B(new_n299), .C1(new_n306), .C2(new_n311), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT36), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G141gat), .B(G148gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(G155gat), .B2(G162gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G148gat), .ZN(new_n330));
  INV_X1    g129(.A(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n339), .B(new_n268), .C1(new_n276), .C2(new_n275), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n338), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n277), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n341), .B1(new_n281), .B2(new_n345), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n279), .A2(KEYINPUT4), .A3(new_n339), .A4(new_n280), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n340), .A2(new_n341), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n351), .A4(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n277), .A2(new_n345), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n351), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n350), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n356), .B1(new_n355), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G57gat), .B(G85gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT6), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n352), .B(new_n368), .C1(new_n361), .C2(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n375), .B(KEYINPUT74), .Z(new_n376));
  NAND2_X1  g175(.A1(new_n238), .A2(new_n286), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n380), .B1(new_n290), .B2(new_n238), .ZN(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n379), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n377), .A2(new_n391), .A3(new_n376), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n224), .A2(new_n237), .B1(new_n253), .B2(new_n256), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT75), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n290), .B2(new_n238), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n392), .B(new_n394), .C1(new_n395), .C2(new_n376), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n390), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  AOI21_X1  g199(.A(KEYINPUT30), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n389), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n379), .A2(new_n381), .ZN(new_n403));
  INV_X1    g202(.A(new_n389), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n405), .A3(new_n400), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n400), .B(KEYINPUT76), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n406), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n401), .B1(new_n408), .B2(KEYINPUT30), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n374), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n343), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n345), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n344), .A2(new_n378), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n389), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n414), .A3(G22gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(G22gat), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  OAI211_X1 g216(.A(G228gat), .B(G233gat), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT31), .B(G50gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  AND2_X1   g220(.A1(new_n421), .A2(KEYINPUT79), .ZN(new_n422));
  INV_X1    g221(.A(new_n417), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n415), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n418), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n421), .A2(KEYINPUT79), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(new_n418), .B2(new_n425), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n320), .A2(KEYINPUT73), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n318), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n321), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n348), .A2(new_n349), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n359), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n358), .A2(new_n359), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n359), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n368), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n363), .A2(new_n369), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n443), .A2(KEYINPUT40), .A3(new_n368), .A4(new_n444), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n431), .B1(new_n450), .B2(new_n409), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n452));
  NAND2_X1  g251(.A1(new_n397), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n400), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n397), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT38), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n396), .B2(new_n389), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n404), .B2(new_n403), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n396), .A2(new_n458), .A3(new_n389), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT37), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n407), .A2(KEYINPUT38), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n453), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n457), .A2(new_n464), .A3(new_n406), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n373), .A2(KEYINPUT82), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n374), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n451), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n437), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n316), .A2(new_n431), .A3(new_n317), .ZN(new_n473));
  INV_X1    g272(.A(new_n409), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n369), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n371), .B2(new_n370), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n466), .B1(new_n477), .B2(KEYINPUT82), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT35), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n316), .A2(new_n431), .A3(KEYINPUT83), .A4(new_n317), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n410), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n484), .B2(new_n479), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n472), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G29gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n488));
  INV_X1    g287(.A(G36gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n487), .B2(KEYINPUT14), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(G29gat), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(G43gat), .A2(G50gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(G43gat), .A2(G50gat), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT15), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n495), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT86), .B(G43gat), .ZN(new_n500));
  INV_X1    g299(.A(G50gat), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT15), .B(new_n496), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n493), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT88), .ZN(new_n505));
  INV_X1    g304(.A(G1gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G8gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT89), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT87), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n503), .A2(new_n512), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n510), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n503), .A2(new_n511), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(KEYINPUT18), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n511), .B(new_n503), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n518), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n531), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n520), .A2(new_n521), .A3(new_n524), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n486), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT90), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT91), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n538), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G71gat), .B2(G78gat), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n541));
  AND2_X1   g340(.A1(G57gat), .A2(G64gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G57gat), .A2(G64gat), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n540), .B(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT21), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n511), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT94), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT93), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT92), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n551), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n545), .A2(new_n546), .ZN(new_n556));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n555), .A2(new_n560), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT97), .B1(new_n564), .B2(KEYINPUT96), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n565), .B(new_n568), .C1(KEYINPUT97), .C2(new_n564), .ZN(new_n569));
  OAI221_X1 g368(.A(KEYINPUT97), .B1(new_n564), .B2(KEYINPUT96), .C1(new_n566), .C2(new_n567), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n566), .B2(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n514), .B(new_n575), .C1(new_n512), .C2(new_n503), .ZN(new_n576));
  INV_X1    g375(.A(new_n575), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n503), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT95), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n563), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G120gat), .B(G148gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT99), .ZN(new_n594));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n575), .B(new_n545), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n598), .A2(G230gat), .A3(G233gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n575), .A2(new_n545), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n598), .B2(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n601), .B(new_n606), .C1(new_n600), .C2(new_n599), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT100), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n596), .B(KEYINPUT101), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n599), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n592), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n537), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n477), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(G1gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(G1324gat));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n474), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n618), .A2(G8gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(KEYINPUT16), .B(G8gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT42), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(KEYINPUT42), .B2(new_n621), .ZN(G1325gat));
  INV_X1    g422(.A(G15gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n624), .A3(new_n319), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n321), .A2(new_n436), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n614), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n625), .B1(new_n629), .B2(new_n624), .ZN(G1326gat));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n432), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT43), .B(G22gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1327gat));
  NOR2_X1   g432(.A1(new_n563), .A2(new_n612), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n590), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT103), .Z(new_n636));
  AND2_X1   g435(.A1(new_n636), .A2(new_n537), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n487), .A3(new_n477), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT45), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n535), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n485), .A2(KEYINPUT104), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n480), .B(new_n644), .C1(new_n484), .C2(new_n479), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n646), .B2(new_n472), .ZN(new_n647));
  AOI211_X1 g446(.A(KEYINPUT105), .B(new_n471), .C1(new_n643), .C2(new_n645), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n590), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n649), .B1(new_n486), .B2(new_n590), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n641), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(G29gat), .B1(new_n653), .B2(new_n374), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n654), .ZN(G1328gat));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n489), .A3(new_n474), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT46), .Z(new_n657));
  OAI21_X1  g456(.A(G36gat), .B1(new_n653), .B2(new_n409), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(G1329gat));
  NOR3_X1   g458(.A1(new_n653), .A2(new_n626), .A3(new_n500), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n319), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n500), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT47), .Z(G1330gat));
  OAI211_X1 g462(.A(new_n432), .B(new_n641), .C1(new_n651), .C2(new_n652), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(G50gat), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n432), .A2(new_n501), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT107), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n636), .A2(new_n537), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(KEYINPUT48), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n665), .B2(KEYINPUT106), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n672), .A3(G50gat), .ZN(new_n673));
  AOI211_X1 g472(.A(KEYINPUT108), .B(KEYINPUT48), .C1(new_n671), .C2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n646), .A2(new_n472), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT105), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n646), .A2(new_n642), .A3(new_n472), .ZN(new_n678));
  INV_X1    g477(.A(new_n650), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n652), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n431), .B(new_n640), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT106), .B1(new_n682), .B2(new_n501), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n673), .A3(new_n668), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT48), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n675), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n669), .B1(new_n674), .B2(new_n686), .ZN(G1331gat));
  NOR2_X1   g486(.A1(new_n647), .A2(new_n648), .ZN(new_n688));
  INV_X1    g487(.A(new_n535), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n612), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n592), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n374), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT109), .B(G57gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1332gat));
  NOR2_X1   g494(.A1(new_n692), .A2(new_n409), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  AND2_X1   g496(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n696), .B2(new_n697), .ZN(G1333gat));
  OR3_X1    g499(.A1(new_n692), .A2(G71gat), .A3(new_n318), .ZN(new_n701));
  OAI21_X1  g500(.A(G71gat), .B1(new_n692), .B2(new_n626), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g503(.A1(new_n692), .A2(new_n431), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(G78gat), .Z(G1335gat));
  INV_X1    g505(.A(KEYINPUT51), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n563), .B1(KEYINPUT110), .B2(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n676), .A2(new_n689), .A3(new_n590), .A4(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n707), .A2(KEYINPUT110), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n612), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713), .B2(new_n477), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n563), .B(new_n690), .C1(new_n680), .C2(new_n681), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n374), .A2(new_n566), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(G1336gat));
  AND2_X1   g516(.A1(new_n715), .A2(new_n474), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n474), .A2(new_n567), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n718), .A2(new_n567), .B1(new_n712), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT52), .ZN(G1337gat));
  AND2_X1   g520(.A1(new_n715), .A2(new_n627), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(KEYINPUT111), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(KEYINPUT111), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(G99gat), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n318), .A2(G99gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n712), .B2(new_n726), .ZN(G1338gat));
  NOR2_X1   g526(.A1(new_n431), .A2(G106gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n612), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT113), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(KEYINPUT53), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(KEYINPUT113), .ZN(new_n732));
  INV_X1    g531(.A(G106gat), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n715), .A2(new_n432), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n731), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n729), .B(KEYINPUT112), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n734), .A2(new_n733), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT53), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(G1339gat));
  NOR3_X1   g538(.A1(new_n592), .A2(new_n535), .A3(new_n612), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n522), .A2(new_n523), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n517), .A2(new_n518), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n530), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT116), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(KEYINPUT116), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n534), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n591), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n597), .B1(new_n606), .B2(KEYINPUT54), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n604), .A2(new_n605), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(KEYINPUT54), .A3(new_n606), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n608), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n756), .B2(new_n757), .ZN(new_n761));
  INV_X1    g560(.A(new_n756), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n759), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n612), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n746), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n764), .B2(new_n535), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n590), .ZN(new_n769));
  INV_X1    g568(.A(new_n563), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n740), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n374), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n475), .ZN(new_n773));
  OAI21_X1  g572(.A(G113gat), .B1(new_n773), .B2(new_n689), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n482), .A2(new_n483), .ZN(new_n775));
  NOR4_X1   g574(.A1(new_n771), .A2(new_n374), .A3(new_n474), .A4(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n267), .A3(new_n535), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(G1340gat));
  NOR3_X1   g577(.A1(new_n773), .A2(new_n265), .A3(new_n766), .ZN(new_n779));
  AOI21_X1  g578(.A(G120gat), .B1(new_n776), .B2(new_n612), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(G1341gat));
  NOR3_X1   g580(.A1(new_n773), .A2(new_n261), .A3(new_n770), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n776), .A2(new_n563), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(KEYINPUT117), .ZN(new_n784));
  AOI21_X1  g583(.A(G127gat), .B1(new_n783), .B2(KEYINPUT117), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n782), .B1(new_n784), .B2(new_n785), .ZN(G1342gat));
  NAND3_X1  g585(.A1(new_n776), .A2(new_n259), .A3(new_n590), .ZN(new_n787));
  XNOR2_X1  g586(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G134gat), .B1(new_n773), .B2(new_n591), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(G1343gat));
  NOR3_X1   g591(.A1(new_n627), .A2(new_n374), .A3(new_n474), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n432), .A2(KEYINPUT57), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n746), .A2(new_n766), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n764), .A2(new_n535), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n590), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n765), .B1(new_n797), .B2(KEYINPUT119), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n768), .A2(new_n799), .A3(new_n590), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n770), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n740), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n794), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n765), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n770), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n802), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT57), .B1(new_n806), .B2(new_n432), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n535), .B(new_n793), .C1(new_n803), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G141gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n626), .A2(new_n432), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n409), .B1(new_n810), .B2(KEYINPUT120), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(KEYINPUT120), .B2(new_n810), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n772), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n329), .A3(new_n535), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT58), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(new_n771), .B2(new_n431), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n799), .B1(new_n768), .B2(new_n590), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n797), .A2(KEYINPUT119), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(new_n765), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n740), .B1(new_n823), .B2(new_n770), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n820), .B1(new_n824), .B2(new_n794), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n825), .A2(KEYINPUT121), .A3(new_n535), .A4(new_n793), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n818), .A2(G141gat), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n816), .B1(new_n827), .B2(new_n829), .ZN(G1344gat));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n331), .A3(new_n612), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n771), .A2(new_n819), .A3(new_n431), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(new_n807), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n612), .A3(new_n793), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n835), .B2(G148gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n832), .A2(G148gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n825), .A2(new_n793), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n837), .B1(new_n839), .B2(new_n612), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n831), .B1(new_n836), .B2(new_n840), .ZN(G1345gat));
  OAI21_X1  g640(.A(G155gat), .B1(new_n838), .B2(new_n770), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n813), .A2(new_n335), .A3(new_n563), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1346gat));
  OAI21_X1  g643(.A(G162gat), .B1(new_n838), .B2(new_n591), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n813), .A2(new_n336), .A3(new_n590), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n477), .A2(new_n409), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n319), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT123), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n432), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n806), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n209), .A3(new_n689), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n771), .B2(new_n477), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n806), .A2(KEYINPUT122), .A3(new_n374), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n775), .A2(new_n409), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n535), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n854), .B1(new_n861), .B2(new_n209), .ZN(G1348gat));
  AOI21_X1  g661(.A(G176gat), .B1(new_n860), .B2(new_n612), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n766), .B1(new_n208), .B2(new_n210), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n852), .B2(new_n864), .ZN(G1349gat));
  NAND4_X1  g664(.A1(new_n858), .A2(new_n283), .A3(new_n563), .A4(new_n859), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n852), .A2(new_n563), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G183gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(KEYINPUT124), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g668(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(G1350gat));
  AOI21_X1  g670(.A(new_n243), .B1(new_n852), .B2(new_n590), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT61), .Z(new_n873));
  NAND3_X1  g672(.A1(new_n860), .A2(new_n243), .A3(new_n590), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1351gat));
  AND2_X1   g674(.A1(new_n626), .A2(new_n848), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n834), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G197gat), .B1(new_n877), .B2(new_n689), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n810), .A2(new_n409), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n856), .B2(new_n857), .ZN(new_n881));
  INV_X1    g680(.A(G197gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n535), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n878), .B1(new_n885), .B2(new_n886), .ZN(G1352gat));
  NOR2_X1   g686(.A1(new_n766), .A2(G204gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n771), .A2(new_n855), .A3(new_n477), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT122), .B1(new_n806), .B2(new_n374), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n879), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT127), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n881), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT62), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n834), .A2(new_n612), .A3(new_n876), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G204gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(G1353gat));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n384), .A3(new_n563), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n834), .A2(new_n563), .A3(new_n876), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n903), .B2(G211gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(G1354gat));
  OAI21_X1  g705(.A(G218gat), .B1(new_n877), .B2(new_n591), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n385), .A3(new_n590), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1355gat));
endmodule


