//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n469), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n466), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n468), .A3(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR3_X1   g056(.A1(new_n472), .A2(new_n476), .A3(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(new_n467), .A2(new_n469), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G2105), .A3(new_n465), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n468), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n470), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n467), .A3(new_n492), .A4(new_n469), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n473), .A2(new_n469), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n493), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G114), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n468), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n496), .A2(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT69), .B1(new_n513), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n511), .A3(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n513), .A2(G651), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  AND3_X1   g095(.A1(new_n517), .A2(new_n518), .A3(new_n509), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n512), .A2(new_n520), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n521), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n525), .A2(KEYINPUT70), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT70), .B1(new_n525), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n519), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n509), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(G651), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(G43), .A2(new_n519), .B1(new_n521), .B2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AND2_X1   g130(.A1(new_n517), .A2(new_n518), .ZN(new_n556));
  AND2_X1   g131(.A1(G53), .A2(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT73), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n556), .A2(new_n563), .A3(new_n557), .A4(new_n558), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n541), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(G651), .A2(new_n568), .B1(new_n521), .B2(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n519), .A2(G49), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n521), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n507), .B2(new_n508), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n517), .A2(G48), .A3(G543), .A4(new_n518), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n517), .A2(G86), .A3(new_n518), .A4(new_n509), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(G72), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G60), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n541), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n511), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(new_n586), .B2(new_n585), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n521), .A2(G85), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT75), .B(G47), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n519), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n521), .A2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT76), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n511), .B1(new_n597), .B2(KEYINPUT76), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n598), .A2(new_n599), .B1(G54), .B2(new_n519), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n593), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  XOR2_X1   g183(.A(KEYINPUT77), .B(G559), .Z(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(G860), .B2(new_n609), .ZN(G148));
  NAND2_X1  g185(.A1(new_n602), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(G123), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n616), .A2(new_n468), .A3(G111), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n468), .B2(G111), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(G2104), .A3(new_n619), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n484), .A2(new_n615), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(G135), .B2(new_n489), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n478), .A2(new_n480), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n494), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT78), .B(G2100), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1956), .B(G2474), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n662), .C2(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT81), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  MUX2_X1   g252(.A(G6), .B(G305), .S(G16), .Z(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT85), .Z(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT32), .B(G1981), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n684), .ZN(new_n686));
  INV_X1    g261(.A(G1971), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(G23), .ZN(new_n689));
  INV_X1    g264(.A(G288), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n684), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n682), .A2(new_n683), .A3(new_n688), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT86), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n489), .A2(G131), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT82), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n484), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(G119), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n700), .B1(new_n709), .B2(new_n699), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  MUX2_X1   g291(.A(G24), .B(G290), .S(G16), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1986), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n697), .A2(new_n698), .A3(new_n715), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G4), .A2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n602), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT88), .B(G1348), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n684), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n550), .B2(new_n684), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1341), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n699), .A2(G26), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g306(.A(G128), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n468), .A2(G116), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n484), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n489), .A2(G140), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n699), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2067), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n726), .A2(new_n729), .A3(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT89), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT89), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G35), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G162), .B2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n746), .A2(G2090), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n684), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n684), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n684), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n684), .ZN(new_n753));
  OAI22_X1  g328(.A1(new_n750), .A2(new_n751), .B1(G1966), .B2(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n747), .B(new_n754), .C1(G1966), .C2(new_n753), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n741), .A2(new_n742), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n699), .A2(G32), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n489), .A2(G141), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT26), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n626), .A2(G105), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G129), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n758), .B(new_n763), .C1(new_n764), .C2(new_n484), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n757), .B1(new_n770), .B2(new_n699), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT27), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1996), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n684), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G33), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT90), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT25), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n489), .B2(G139), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(G2105), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n781), .B1(new_n789), .B2(new_n699), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT92), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2072), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n750), .A2(new_n751), .B1(G2090), .B2(new_n746), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G160), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n699), .B1(new_n796), .B2(G34), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(G34), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n797), .B2(KEYINPUT93), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n795), .A2(new_n699), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G2084), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT94), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n699), .A2(G27), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G164), .B2(new_n699), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G2078), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(G2078), .ZN(new_n809));
  INV_X1    g384(.A(G28), .ZN(new_n810));
  AOI21_X1  g385(.A(G29), .B1(new_n810), .B2(KEYINPUT30), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(KEYINPUT30), .B2(new_n810), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G11), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G11), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n622), .B2(G29), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n805), .A2(new_n808), .A3(new_n809), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n794), .A2(new_n804), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n773), .A2(new_n779), .A3(new_n792), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n756), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n722), .A2(new_n822), .ZN(G311));
  INV_X1    g398(.A(new_n721), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n720), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n821), .ZN(G150));
  NAND2_X1  g401(.A1(new_n602), .A2(G559), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT38), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n521), .A2(G93), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n519), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n829), .B(new_n830), .C1(new_n511), .C2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n549), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n549), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n828), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n832), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n708), .B(new_n628), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n489), .A2(G142), .ZN(new_n845));
  INV_X1    g420(.A(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n468), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI221_X1 g423(.A(new_n845), .B1(new_n484), .B2(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n789), .ZN(new_n853));
  INV_X1    g428(.A(new_n737), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n769), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n769), .A2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n500), .A2(new_n502), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n504), .B1(new_n860), .B2(G2105), .ZN(new_n861));
  AND4_X1   g436(.A1(new_n465), .A2(new_n467), .A3(new_n469), .A4(new_n497), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n504), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT68), .B(G114), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(new_n468), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(KEYINPUT99), .A3(new_n498), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n496), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n770), .A2(new_n737), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(new_n789), .A3(new_n855), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n858), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n868), .B1(new_n858), .B2(new_n870), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n852), .B(KEYINPUT101), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n850), .B(KEYINPUT100), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n622), .B(new_n795), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(KEYINPUT102), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n876), .B2(new_n850), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n883), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n883), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  OR2_X1    g464(.A1(new_n601), .A2(G299), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n601), .A2(G299), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n892), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n892), .B2(KEYINPUT41), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n836), .B(new_n611), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n892), .B(KEYINPUT103), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G303), .B(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(G290), .B(new_n690), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(KEYINPUT106), .A3(new_n903), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n605), .B1(new_n902), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n832), .B2(new_n605), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(G295));
  AOI21_X1  g494(.A(new_n916), .B1(new_n915), .B2(new_n918), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n835), .B(G301), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G168), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n836), .A2(G301), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n835), .A2(G171), .ZN(new_n925));
  OAI21_X1  g500(.A(G286), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n892), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n911), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(new_n934), .C1(new_n932), .C2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(new_n892), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n932), .B(new_n937), .C1(new_n898), .C2(new_n928), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n892), .A2(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n894), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n923), .A2(new_n926), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n911), .B(new_n941), .C1(new_n929), .C2(new_n901), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n921), .B1(new_n935), .B2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n933), .A2(KEYINPUT109), .A3(new_n942), .A4(new_n934), .ZN(new_n947));
  INV_X1    g522(.A(new_n934), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n938), .A2(new_n943), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n931), .A2(new_n932), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n938), .A2(new_n942), .A3(new_n943), .A4(new_n934), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n947), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n946), .B1(new_n955), .B2(new_n921), .ZN(G397));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n868), .B2(G1384), .ZN(new_n958));
  INV_X1    g533(.A(new_n476), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n483), .A2(G137), .A3(new_n468), .A4(new_n465), .ZN(new_n960));
  INV_X1    g535(.A(new_n481), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n959), .A2(new_n960), .A3(G40), .A4(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(G1996), .A3(new_n769), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT110), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n737), .B(G2067), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n769), .B2(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n963), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n708), .B(new_n712), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n963), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(G290), .B(G1986), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n963), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT124), .ZN(new_n976));
  INV_X1    g551(.A(new_n496), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n866), .A2(KEYINPUT99), .A3(new_n498), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT99), .B1(new_n866), .B2(new_n498), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2078), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n496), .B2(new_n505), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n957), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n472), .A2(new_n476), .A3(new_n481), .A4(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n982), .A2(new_n983), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n868), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n987), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n751), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT45), .B(new_n981), .C1(new_n496), .C2(new_n505), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n987), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n989), .A2(G2078), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n958), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(G171), .B1(new_n990), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G171), .B1(new_n988), .B2(new_n989), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n958), .A2(new_n982), .A3(new_n987), .A4(new_n997), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT123), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n863), .A2(new_n867), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n977), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n962), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(KEYINPUT123), .A3(new_n958), .A4(new_n997), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1001), .A2(new_n1004), .A3(new_n1008), .A4(new_n994), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1000), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n988), .A2(new_n989), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1004), .A2(new_n1008), .A3(new_n1012), .A4(new_n994), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G171), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n1015));
  INV_X1    g590(.A(new_n999), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n1001), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1010), .A2(new_n1011), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT113), .B(G8), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n980), .A2(new_n1021), .A3(new_n981), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n962), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(G2084), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1966), .B1(new_n958), .B2(new_n996), .ZN(new_n1026));
  OAI211_X1 g601(.A(G286), .B(new_n1020), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G168), .A2(new_n1019), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n980), .B2(new_n981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n987), .A2(new_n995), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1029), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1027), .B(KEYINPUT51), .C1(new_n1028), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1019), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1028), .A2(KEYINPUT51), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1018), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n868), .A2(G1384), .A3(new_n962), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G305), .A2(G1981), .ZN(new_n1046));
  INV_X1    g621(.A(G1981), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1045), .A2(new_n1049), .A3(new_n1019), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1046), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n1048), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1045), .A2(new_n1019), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n690), .A2(G1976), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n980), .A2(new_n981), .A3(new_n987), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1063), .A3(new_n1020), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1021), .B1(new_n980), .B2(new_n981), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n962), .ZN(new_n1069));
  INV_X1    g644(.A(G2090), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT115), .B(new_n987), .C1(new_n1006), .C2(new_n1021), .ZN(new_n1071));
  INV_X1    g646(.A(new_n984), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1021), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n982), .A2(new_n985), .A3(new_n987), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n687), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1020), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G303), .A2(G8), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT55), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1066), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1075), .A2(KEYINPUT111), .A3(new_n687), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1022), .A2(new_n1023), .A3(new_n1070), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1080), .ZN(new_n1089));
  AND4_X1   g664(.A1(new_n1082), .A2(new_n1088), .A3(G8), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1029), .B1(new_n1091), .B2(new_n1085), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1082), .B1(new_n1092), .B2(new_n1089), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1081), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n976), .B1(new_n1044), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT121), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1066), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1019), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1101), .B2(new_n1089), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1088), .A2(G8), .A3(new_n1089), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT112), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1092), .A2(new_n1082), .A3(new_n1089), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1099), .A2(new_n1106), .A3(KEYINPUT124), .A4(new_n1018), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n565), .A2(new_n1109), .A3(new_n569), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1073), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n980), .A2(new_n981), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n962), .B1(new_n1113), .B2(KEYINPUT50), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1114), .B2(KEYINPUT115), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1956), .B1(new_n1115), .B2(new_n1069), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT56), .B(G2072), .Z(new_n1117));
  NOR2_X1   g692(.A1(new_n1075), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1069), .A2(new_n1073), .A3(new_n1071), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1121), .B2(new_n778), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1111), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1348), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n991), .B2(new_n993), .ZN(new_n1126));
  INV_X1    g701(.A(G2067), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1045), .A2(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1129), .A2(new_n601), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1120), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1118), .B(new_n1111), .C1(new_n1121), .C2(new_n778), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1135), .B(new_n1111), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1119), .A2(KEYINPUT61), .A3(new_n1124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1063), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n982), .A2(new_n1145), .A3(new_n985), .A4(new_n987), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1063), .A2(new_n1147), .A3(new_n1142), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1150));
  AND3_X1   g725(.A1(new_n1149), .A2(new_n550), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n1128), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT60), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1153), .B2(new_n601), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1129), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1141), .A2(new_n1151), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n550), .A3(new_n1150), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1149), .A2(new_n550), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT59), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT119), .B(new_n1157), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1140), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1131), .B1(new_n1139), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1095), .A2(new_n1107), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1097), .A2(KEYINPUT62), .A3(new_n1098), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1000), .B(new_n1102), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1057), .A2(new_n1060), .A3(new_n690), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1045), .B(new_n1019), .C1(new_n1170), .C2(new_n1048), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1050), .A2(new_n1056), .B1(new_n1064), .B2(KEYINPUT52), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(G168), .A3(new_n1062), .A4(new_n1038), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1088), .A2(G8), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1175), .B2(new_n1080), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1172), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1038), .A2(G168), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(KEYINPUT63), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1093), .B2(new_n1090), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1178), .B1(new_n1100), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1169), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n975), .B1(new_n1163), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n969), .A2(new_n712), .A3(new_n708), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n854), .A2(G2067), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n963), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n1145), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT46), .ZN(new_n1192));
  INV_X1    g767(.A(new_n963), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n770), .A2(new_n966), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT47), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1193), .A2(G1986), .A3(G290), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT48), .Z(new_n1198));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1190), .A2(new_n1196), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1186), .A2(new_n1187), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1066), .A2(new_n1180), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1171), .B1(new_n1204), .B2(KEYINPUT63), .ZN(new_n1205));
  AOI22_X1  g780(.A1(new_n1104), .A2(new_n1105), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(new_n1066), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1095), .A2(new_n1162), .A3(new_n1107), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n974), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT125), .B1(new_n1210), .B2(new_n1200), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1202), .A2(new_n1211), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g787(.A1(new_n947), .A2(new_n951), .A3(new_n954), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n883), .A2(new_n886), .ZN(new_n1215));
  OR3_X1    g789(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1216));
  XNOR2_X1  g790(.A(new_n1216), .B(KEYINPUT126), .ZN(new_n1217));
  NOR2_X1   g791(.A1(G229), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n1214), .A2(new_n1215), .A3(new_n1218), .ZN(G225));
  INV_X1    g793(.A(G225), .ZN(G308));
endmodule


