

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788;

  NAND2_X1 U376 ( .A1(n656), .A2(G953), .ZN(n716) );
  XNOR2_X1 U377 ( .A(n653), .B(KEYINPUT59), .ZN(n654) );
  XNOR2_X1 U378 ( .A(n713), .B(n712), .ZN(n714) );
  OR2_X1 U379 ( .A1(n649), .A2(n394), .ZN(n374) );
  XNOR2_X1 U380 ( .A(G113), .B(KEYINPUT71), .ZN(n499) );
  AND2_X2 U381 ( .A1(n373), .A2(KEYINPUT64), .ZN(n370) );
  AND2_X2 U382 ( .A1(n470), .A2(n468), .ZN(n467) );
  NOR2_X2 U383 ( .A1(n758), .A2(n756), .ZN(n597) );
  XNOR2_X2 U384 ( .A(n597), .B(KEYINPUT41), .ZN(n738) );
  NAND2_X2 U385 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X2 U386 ( .A1(n458), .A2(n456), .ZN(n593) );
  XNOR2_X2 U387 ( .A(n354), .B(n537), .ZN(n563) );
  NAND2_X2 U388 ( .A1(n467), .A2(n465), .ZN(n354) );
  XNOR2_X1 U389 ( .A(KEYINPUT68), .B(G131), .ZN(n542) );
  XNOR2_X1 U390 ( .A(G110), .B(G107), .ZN(n476) );
  BUF_X1 U391 ( .A(n784), .Z(n357) );
  XNOR2_X1 U392 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n355) );
  NOR2_X1 U393 ( .A1(n641), .A2(n626), .ZN(n445) );
  AND2_X1 U394 ( .A1(n588), .A2(n666), .ZN(n589) );
  NAND2_X1 U395 ( .A1(n363), .A2(n587), .ZN(n666) );
  OR2_X1 U396 ( .A1(n729), .A2(n721), .ZN(n584) );
  XNOR2_X1 U397 ( .A(n445), .B(n355), .ZN(n367) );
  AND2_X1 U398 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U399 ( .A(n596), .B(KEYINPUT112), .ZN(n758) );
  NOR2_X1 U400 ( .A1(n368), .A2(n755), .ZN(n447) );
  XNOR2_X1 U401 ( .A(n553), .B(n552), .ZN(n580) );
  XNOR2_X1 U402 ( .A(n701), .B(n703), .ZN(n704) );
  XNOR2_X1 U403 ( .A(n507), .B(n480), .ZN(n701) );
  OR2_X1 U404 ( .A1(n472), .A2(n647), .ZN(n393) );
  INV_X1 U405 ( .A(G902), .ZN(n440) );
  INV_X1 U406 ( .A(KEYINPUT36), .ZN(n436) );
  AND2_X1 U407 ( .A1(n371), .A2(n374), .ZN(n364) );
  NAND2_X1 U408 ( .A1(n365), .A2(n405), .ZN(n403) );
  XNOR2_X1 U409 ( .A(n366), .B(n404), .ZN(n365) );
  NAND2_X1 U410 ( .A1(n589), .A2(KEYINPUT90), .ZN(n449) );
  OR2_X1 U411 ( .A1(n590), .A2(n666), .ZN(n420) );
  NAND2_X1 U412 ( .A1(n446), .A2(n367), .ZN(n366) );
  NAND2_X1 U413 ( .A1(n435), .A2(n434), .ZN(n682) );
  XNOR2_X1 U414 ( .A(n367), .B(G131), .ZN(G33) );
  NAND2_X2 U415 ( .A1(n380), .A2(n376), .ZN(n446) );
  XNOR2_X1 U416 ( .A(n437), .B(n436), .ZN(n435) );
  OR2_X1 U417 ( .A1(n664), .A2(KEYINPUT47), .ZN(n401) );
  NAND2_X1 U418 ( .A1(n379), .A2(n378), .ZN(n377) );
  XNOR2_X1 U419 ( .A(n757), .B(n426), .ZN(n583) );
  NAND2_X1 U420 ( .A1(n408), .A2(n407), .ZN(n615) );
  XNOR2_X1 U421 ( .A(n410), .B(n409), .ZN(n408) );
  NAND2_X1 U422 ( .A1(n368), .A2(n755), .ZN(n596) );
  NAND2_X1 U423 ( .A1(n573), .A2(n575), .ZN(n576) );
  XNOR2_X1 U424 ( .A(n383), .B(n498), .ZN(n422) );
  NAND2_X1 U425 ( .A1(n448), .A2(n384), .ZN(n383) );
  NAND2_X1 U426 ( .A1(n466), .A2(n530), .ZN(n465) );
  NAND2_X2 U427 ( .A1(n442), .A2(n438), .ZN(n745) );
  AND2_X1 U428 ( .A1(n444), .A2(n443), .ZN(n442) );
  XOR2_X1 U429 ( .A(KEYINPUT62), .B(n687), .Z(n688) );
  OR2_X1 U430 ( .A1(KEYINPUT88), .A2(n472), .ZN(n394) );
  NOR2_X1 U431 ( .A1(n647), .A2(n646), .ZN(n472) );
  XNOR2_X1 U432 ( .A(n413), .B(n440), .ZN(n644) );
  NAND2_X1 U433 ( .A1(n590), .A2(KEYINPUT44), .ZN(n455) );
  XNOR2_X1 U434 ( .A(n395), .B(G469), .ZN(n385) );
  XNOR2_X1 U435 ( .A(KEYINPUT16), .B(G122), .ZN(n521) );
  XNOR2_X2 U436 ( .A(G116), .B(KEYINPUT9), .ZN(n432) );
  XNOR2_X2 U437 ( .A(G107), .B(KEYINPUT99), .ZN(n427) );
  XNOR2_X1 U438 ( .A(G140), .B(KEYINPUT10), .ZN(n483) );
  XNOR2_X2 U439 ( .A(G122), .B(KEYINPUT100), .ZN(n428) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n531) );
  XNOR2_X2 U441 ( .A(G146), .B(G125), .ZN(n515) );
  XNOR2_X2 U442 ( .A(G116), .B(G101), .ZN(n500) );
  XNOR2_X1 U443 ( .A(KEYINPUT95), .B(KEYINPUT15), .ZN(n413) );
  INV_X2 U444 ( .A(G953), .ZN(n784) );
  XOR2_X1 U445 ( .A(G113), .B(G122), .Z(n541) );
  XNOR2_X1 U446 ( .A(G119), .B(G137), .ZN(n484) );
  XNOR2_X1 U447 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n488) );
  INV_X1 U448 ( .A(KEYINPUT42), .ZN(n378) );
  NAND2_X1 U449 ( .A1(n356), .A2(n623), .ZN(n624) );
  NAND2_X1 U450 ( .A1(n399), .A2(n401), .ZN(n356) );
  NOR2_X2 U451 ( .A1(n728), .A2(n581), .ZN(n582) );
  NAND2_X1 U452 ( .A1(n389), .A2(n390), .ZN(n392) );
  NOR2_X1 U453 ( .A1(n735), .A2(n372), .ZN(n371) );
  XNOR2_X2 U454 ( .A(n593), .B(KEYINPUT45), .ZN(n648) );
  XNOR2_X1 U455 ( .A(n571), .B(n570), .ZN(n683) );
  BUF_X1 U456 ( .A(n466), .Z(n358) );
  BUF_X2 U457 ( .A(n648), .Z(n777) );
  NAND2_X1 U458 ( .A1(n359), .A2(n455), .ZN(n362) );
  INV_X1 U459 ( .A(n369), .ZN(n359) );
  NAND2_X1 U460 ( .A1(n360), .A2(n450), .ZN(n458) );
  NAND2_X1 U461 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U462 ( .A1(n369), .A2(n449), .ZN(n361) );
  NOR2_X2 U463 ( .A1(n572), .A2(n576), .ZN(n667) );
  INV_X1 U464 ( .A(n572), .ZN(n363) );
  BUF_X2 U465 ( .A(n594), .Z(n617) );
  NAND2_X1 U466 ( .A1(n364), .A2(n373), .ZN(n389) );
  NAND2_X1 U467 ( .A1(n370), .A2(n364), .ZN(n391) );
  NAND2_X1 U468 ( .A1(n620), .A2(n368), .ZN(n612) );
  XNOR2_X2 U469 ( .A(n617), .B(n595), .ZN(n368) );
  NOR2_X2 U470 ( .A1(n591), .A2(n685), .ZN(n369) );
  XNOR2_X2 U471 ( .A(n375), .B(KEYINPUT80), .ZN(n373) );
  NAND2_X1 U472 ( .A1(n652), .A2(n393), .ZN(n372) );
  NAND2_X1 U473 ( .A1(n373), .A2(n652), .ZN(n736) );
  NOR2_X2 U474 ( .A1(n777), .A2(KEYINPUT2), .ZN(n735) );
  NAND2_X1 U475 ( .A1(n649), .A2(KEYINPUT2), .ZN(n375) );
  OR2_X1 U476 ( .A1(n738), .A2(n377), .ZN(n376) );
  INV_X1 U477 ( .A(n615), .ZN(n379) );
  NAND2_X1 U478 ( .A1(n615), .A2(KEYINPUT42), .ZN(n381) );
  NAND2_X1 U479 ( .A1(n738), .A2(KEYINPUT42), .ZN(n382) );
  XNOR2_X1 U480 ( .A(n418), .B(n385), .ZN(n384) );
  XNOR2_X1 U481 ( .A(n513), .B(G134), .ZN(n556) );
  XNOR2_X1 U482 ( .A(n387), .B(n395), .ZN(n386) );
  XNOR2_X2 U483 ( .A(n418), .B(G469), .ZN(n387) );
  XOR2_X1 U484 ( .A(n560), .B(KEYINPUT35), .Z(n388) );
  NAND2_X2 U485 ( .A1(n391), .A2(n392), .ZN(n708) );
  INV_X1 U486 ( .A(KEYINPUT64), .ZN(n390) );
  INV_X1 U487 ( .A(n573), .ZN(n434) );
  OR2_X1 U488 ( .A1(n762), .A2(n540), .ZN(n459) );
  INV_X1 U489 ( .A(n739), .ZN(n448) );
  NAND2_X1 U490 ( .A1(n627), .A2(n745), .ZN(n410) );
  NAND2_X1 U491 ( .A1(KEYINPUT90), .A2(n453), .ZN(n452) );
  INV_X1 U492 ( .A(KEYINPUT92), .ZN(n411) );
  XNOR2_X1 U493 ( .A(n481), .B(KEYINPUT20), .ZN(n495) );
  XNOR2_X1 U494 ( .A(n406), .B(KEYINPUT69), .ZN(n405) );
  NAND2_X1 U495 ( .A1(n633), .A2(n682), .ZN(n406) );
  XNOR2_X1 U496 ( .A(KEYINPUT4), .B(G137), .ZN(n474) );
  AND2_X1 U497 ( .A1(n632), .A2(n755), .ZN(n634) );
  NAND2_X1 U498 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U499 ( .A1(n495), .A2(G217), .ZN(n415) );
  INV_X1 U500 ( .A(G472), .ZN(n441) );
  NAND2_X1 U501 ( .A1(G902), .A2(G472), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n509), .B(KEYINPUT33), .ZN(n762) );
  INV_X1 U503 ( .A(KEYINPUT28), .ZN(n409) );
  INV_X1 U504 ( .A(KEYINPUT86), .ZN(n426) );
  INV_X1 U505 ( .A(KEYINPUT46), .ZN(n404) );
  AND2_X1 U506 ( .A1(n419), .A2(n420), .ZN(n454) );
  AND2_X1 U507 ( .A1(n471), .A2(n469), .ZN(n468) );
  OR2_X1 U508 ( .A1(n755), .A2(KEYINPUT19), .ZN(n469) );
  INV_X1 U509 ( .A(G237), .ZN(n524) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n544) );
  XNOR2_X1 U511 ( .A(G143), .B(G104), .ZN(n543) );
  XNOR2_X1 U512 ( .A(KEYINPUT3), .B(G119), .ZN(n501) );
  XNOR2_X1 U513 ( .A(n403), .B(n402), .ZN(n643) );
  INV_X1 U514 ( .A(KEYINPUT48), .ZN(n402) );
  INV_X1 U515 ( .A(KEYINPUT7), .ZN(n433) );
  AND2_X1 U516 ( .A1(n462), .A2(n559), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n463), .A2(KEYINPUT34), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n415), .B(n414), .ZN(n494) );
  XNOR2_X1 U519 ( .A(n482), .B(KEYINPUT25), .ZN(n414) );
  XNOR2_X1 U520 ( .A(n579), .B(KEYINPUT101), .ZN(n728) );
  NAND2_X1 U521 ( .A1(n424), .A2(n561), .ZN(n579) );
  OR2_X1 U522 ( .A1(n687), .A2(n439), .ZN(n438) );
  NAND2_X1 U523 ( .A1(n441), .A2(n440), .ZN(n439) );
  INV_X1 U524 ( .A(n416), .ZN(n572) );
  XNOR2_X1 U525 ( .A(G101), .B(G140), .ZN(n478) );
  NOR2_X2 U526 ( .A1(n615), .A2(n614), .ZN(n664) );
  BUF_X1 U527 ( .A(n728), .Z(n423) );
  INV_X1 U528 ( .A(KEYINPUT19), .ZN(n530) );
  XOR2_X1 U529 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n395) );
  AND2_X1 U530 ( .A1(n569), .A2(n568), .ZN(n396) );
  AND2_X1 U531 ( .A1(n539), .A2(n540), .ZN(n397) );
  AND2_X1 U532 ( .A1(n755), .A2(KEYINPUT19), .ZN(n398) );
  INV_X1 U533 ( .A(KEYINPUT44), .ZN(n453) );
  NAND2_X1 U534 ( .A1(n664), .A2(n400), .ZN(n399) );
  NAND2_X1 U535 ( .A1(n583), .A2(n616), .ZN(n400) );
  INV_X1 U536 ( .A(n387), .ZN(n407) );
  XNOR2_X2 U537 ( .A(n412), .B(n411), .ZN(n591) );
  NOR2_X2 U538 ( .A1(n683), .A2(n667), .ZN(n412) );
  XNOR2_X2 U539 ( .A(n566), .B(n417), .ZN(n416) );
  XOR2_X1 U540 ( .A(n565), .B(n564), .Z(n417) );
  NOR2_X2 U541 ( .A1(n701), .A2(G902), .ZN(n418) );
  NAND2_X1 U542 ( .A1(n584), .A2(n421), .ZN(n419) );
  AND2_X1 U543 ( .A1(n583), .A2(KEYINPUT90), .ZN(n421) );
  XNOR2_X1 U544 ( .A(n577), .B(KEYINPUT31), .ZN(n729) );
  NAND2_X1 U545 ( .A1(n422), .A2(n628), .ZN(n509) );
  AND2_X1 U546 ( .A1(n422), .A2(n745), .ZN(n751) );
  XNOR2_X2 U547 ( .A(n582), .B(KEYINPUT102), .ZN(n757) );
  XNOR2_X1 U548 ( .A(n548), .B(n670), .ZN(n549) );
  XNOR2_X1 U549 ( .A(n549), .B(n550), .ZN(n653) );
  NAND2_X1 U550 ( .A1(n762), .A2(n397), .ZN(n464) );
  AND2_X2 U551 ( .A1(n648), .A2(n673), .ZN(n649) );
  NAND2_X1 U552 ( .A1(n592), .A2(n457), .ZN(n456) );
  AND2_X2 U553 ( .A1(n464), .A2(n461), .ZN(n460) );
  INV_X1 U554 ( .A(n561), .ZN(n425) );
  XNOR2_X2 U555 ( .A(n558), .B(G478), .ZN(n561) );
  INV_X1 U556 ( .A(n580), .ZN(n424) );
  NAND2_X1 U557 ( .A1(n580), .A2(n425), .ZN(n626) );
  XNOR2_X1 U558 ( .A(n428), .B(n427), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n555), .B(n429), .ZN(n557) );
  XNOR2_X1 U560 ( .A(n431), .B(n430), .ZN(n429) );
  XNOR2_X1 U561 ( .A(n432), .B(n433), .ZN(n430) );
  NAND2_X1 U562 ( .A1(n634), .A2(n617), .ZN(n437) );
  NAND2_X1 U563 ( .A1(n687), .A2(G472), .ZN(n444) );
  XNOR2_X2 U564 ( .A(n745), .B(n508), .ZN(n628) );
  XNOR2_X1 U565 ( .A(n446), .B(G137), .ZN(G39) );
  INV_X1 U566 ( .A(n386), .ZN(n573) );
  NAND2_X1 U567 ( .A1(n454), .A2(n451), .ZN(n450) );
  NAND2_X1 U568 ( .A1(n589), .A2(n452), .ZN(n451) );
  XNOR2_X1 U569 ( .A(n591), .B(KEYINPUT91), .ZN(n457) );
  NAND2_X2 U570 ( .A1(n460), .A2(n459), .ZN(n560) );
  INV_X1 U571 ( .A(n539), .ZN(n463) );
  AND2_X1 U572 ( .A1(n617), .A2(n755), .ZN(n613) );
  INV_X1 U573 ( .A(n594), .ZN(n466) );
  NAND2_X1 U574 ( .A1(n594), .A2(n398), .ZN(n470) );
  XNOR2_X2 U575 ( .A(n528), .B(n527), .ZN(n594) );
  OR2_X1 U576 ( .A1(n536), .A2(n600), .ZN(n471) );
  XNOR2_X1 U577 ( .A(n567), .B(KEYINPUT105), .ZN(n569) );
  BUF_X1 U578 ( .A(n738), .Z(n770) );
  XNOR2_X1 U579 ( .A(n551), .B(G475), .ZN(n552) );
  INV_X1 U580 ( .A(KEYINPUT60), .ZN(n658) );
  XNOR2_X2 U581 ( .A(G143), .B(KEYINPUT83), .ZN(n473) );
  XNOR2_X2 U582 ( .A(n473), .B(G128), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n542), .B(n474), .ZN(n475) );
  XNOR2_X2 U584 ( .A(n556), .B(n475), .ZN(n671) );
  XNOR2_X2 U585 ( .A(n671), .B(G146), .ZN(n507) );
  XNOR2_X1 U586 ( .A(n476), .B(G104), .ZN(n783) );
  XNOR2_X1 U587 ( .A(n783), .B(KEYINPUT72), .ZN(n519) );
  NAND2_X1 U588 ( .A1(n357), .A2(G227), .ZN(n477) );
  XNOR2_X1 U589 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n519), .B(n479), .ZN(n480) );
  XOR2_X1 U591 ( .A(KEYINPUT97), .B(KEYINPUT81), .Z(n482) );
  NAND2_X1 U592 ( .A1(n644), .A2(G234), .ZN(n481) );
  XNOR2_X1 U593 ( .A(n483), .B(n515), .ZN(n670) );
  XOR2_X1 U594 ( .A(G110), .B(G128), .Z(n485) );
  XNOR2_X1 U595 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U596 ( .A(n670), .B(n486), .ZN(n492) );
  XOR2_X1 U597 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n490) );
  NAND2_X1 U598 ( .A1(n784), .A2(G234), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n554) );
  AND2_X1 U600 ( .A1(n554), .A2(G221), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n693) );
  AND2_X1 U603 ( .A1(n693), .A2(n440), .ZN(n493) );
  XNOR2_X1 U604 ( .A(n494), .B(n493), .ZN(n603) );
  AND2_X1 U605 ( .A1(n495), .A2(G221), .ZN(n497) );
  INV_X1 U606 ( .A(KEYINPUT21), .ZN(n496) );
  XNOR2_X1 U607 ( .A(n497), .B(n496), .ZN(n743) );
  OR2_X1 U608 ( .A1(n603), .A2(n743), .ZN(n739) );
  INV_X1 U609 ( .A(KEYINPUT78), .ZN(n498) );
  XNOR2_X1 U610 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n502), .B(n501), .ZN(n522) );
  NAND2_X1 U612 ( .A1(n784), .A2(n524), .ZN(n503) );
  XNOR2_X1 U613 ( .A(KEYINPUT79), .B(n503), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n547), .A2(G210), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n504), .B(KEYINPUT5), .ZN(n505) );
  XNOR2_X1 U616 ( .A(n522), .B(n505), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n507), .B(n506), .ZN(n687) );
  XNOR2_X1 U618 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n508) );
  XNOR2_X1 U619 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n511) );
  XNOR2_X1 U620 ( .A(KEYINPUT82), .B(KEYINPUT94), .ZN(n510) );
  XNOR2_X1 U621 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U622 ( .A(n513), .B(n512), .ZN(n518) );
  NAND2_X1 U623 ( .A1(n784), .A2(G224), .ZN(n514) );
  XNOR2_X1 U624 ( .A(n514), .B(KEYINPUT4), .ZN(n516) );
  XNOR2_X1 U625 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U626 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n782) );
  XNOR2_X1 U629 ( .A(n523), .B(n782), .ZN(n709) );
  INV_X1 U630 ( .A(n644), .ZN(n647) );
  OR2_X2 U631 ( .A1(n709), .A2(n647), .ZN(n528) );
  NAND2_X1 U632 ( .A1(n440), .A2(n524), .ZN(n529) );
  NAND2_X1 U633 ( .A1(n529), .A2(G210), .ZN(n526) );
  INV_X1 U634 ( .A(KEYINPUT84), .ZN(n525) );
  XNOR2_X1 U635 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U636 ( .A1(n529), .A2(G214), .ZN(n755) );
  XNOR2_X1 U637 ( .A(n531), .B(KEYINPUT14), .ZN(n532) );
  XNOR2_X1 U638 ( .A(KEYINPUT76), .B(n532), .ZN(n535) );
  AND2_X1 U639 ( .A1(n535), .A2(G953), .ZN(n533) );
  NAND2_X1 U640 ( .A1(G902), .A2(n533), .ZN(n598) );
  NOR2_X1 U641 ( .A1(G898), .A2(n598), .ZN(n534) );
  XNOR2_X1 U642 ( .A(n534), .B(KEYINPUT96), .ZN(n536) );
  NAND2_X1 U643 ( .A1(G952), .A2(n535), .ZN(n768) );
  NOR2_X1 U644 ( .A1(n768), .A2(G953), .ZN(n600) );
  INV_X1 U645 ( .A(KEYINPUT0), .ZN(n537) );
  BUF_X1 U646 ( .A(n563), .Z(n539) );
  INV_X1 U647 ( .A(KEYINPUT34), .ZN(n540) );
  XNOR2_X1 U648 ( .A(n542), .B(n541), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U650 ( .A(n546), .B(n545), .Z(n550) );
  NAND2_X1 U651 ( .A1(G214), .A2(n547), .ZN(n548) );
  NOR2_X1 U652 ( .A1(G902), .A2(n653), .ZN(n553) );
  XNOR2_X1 U653 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n551) );
  NAND2_X1 U654 ( .A1(n554), .A2(G217), .ZN(n555) );
  XNOR2_X1 U655 ( .A(n556), .B(n557), .ZN(n698) );
  NAND2_X1 U656 ( .A1(n698), .A2(n440), .ZN(n558) );
  NAND2_X1 U657 ( .A1(n580), .A2(n561), .ZN(n618) );
  INV_X1 U658 ( .A(n618), .ZN(n559) );
  XNOR2_X2 U659 ( .A(n560), .B(KEYINPUT35), .ZN(n685) );
  OR2_X1 U660 ( .A1(n580), .A2(n561), .ZN(n756) );
  NOR2_X1 U661 ( .A1(n756), .A2(n743), .ZN(n562) );
  NAND2_X1 U662 ( .A1(n563), .A2(n562), .ZN(n566) );
  XNOR2_X1 U663 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n565) );
  INV_X1 U664 ( .A(KEYINPUT73), .ZN(n564) );
  XNOR2_X1 U665 ( .A(n603), .B(KEYINPUT104), .ZN(n742) );
  NAND2_X1 U666 ( .A1(n386), .A2(n742), .ZN(n567) );
  INV_X1 U667 ( .A(n628), .ZN(n568) );
  NAND2_X1 U668 ( .A1(n416), .A2(n396), .ZN(n571) );
  XNOR2_X1 U669 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n570) );
  INV_X1 U670 ( .A(n603), .ZN(n574) );
  NOR2_X1 U671 ( .A1(n745), .A2(n574), .ZN(n575) );
  NAND2_X1 U672 ( .A1(n751), .A2(n539), .ZN(n577) );
  OR2_X1 U673 ( .A1(n739), .A2(n387), .ZN(n608) );
  NOR2_X1 U674 ( .A1(n608), .A2(n745), .ZN(n578) );
  AND2_X1 U675 ( .A1(n539), .A2(n578), .ZN(n721) );
  INV_X1 U676 ( .A(n626), .ZN(n581) );
  NAND2_X1 U677 ( .A1(n584), .A2(n583), .ZN(n588) );
  INV_X1 U678 ( .A(n742), .ZN(n585) );
  NAND2_X1 U679 ( .A1(n573), .A2(n585), .ZN(n586) );
  NOR2_X1 U680 ( .A1(n586), .A2(n628), .ZN(n587) );
  INV_X1 U681 ( .A(KEYINPUT90), .ZN(n590) );
  AND2_X1 U682 ( .A1(n388), .A2(n453), .ZN(n592) );
  XNOR2_X1 U683 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n595) );
  NOR2_X1 U684 ( .A1(G900), .A2(n598), .ZN(n599) );
  XOR2_X1 U685 ( .A(KEYINPUT107), .B(n599), .Z(n601) );
  NOR2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n743), .A2(n607), .ZN(n602) );
  XNOR2_X1 U688 ( .A(n602), .B(KEYINPUT70), .ZN(n604) );
  AND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n627) );
  NAND2_X1 U690 ( .A1(n745), .A2(n755), .ZN(n606) );
  INV_X1 U691 ( .A(KEYINPUT30), .ZN(n605) );
  XNOR2_X1 U692 ( .A(n606), .B(n605), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n620) );
  INV_X1 U695 ( .A(KEYINPUT39), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n612), .B(n611), .ZN(n641) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT19), .ZN(n614) );
  INV_X1 U698 ( .A(KEYINPUT47), .ZN(n616) );
  NAND2_X1 U699 ( .A1(n757), .A2(KEYINPUT47), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n618), .A2(n358), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n661) );
  NAND2_X1 U702 ( .A1(n621), .A2(n661), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n622), .B(KEYINPUT85), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT75), .ZN(n633) );
  INV_X1 U705 ( .A(KEYINPUT106), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n626), .B(n625), .ZN(n725) );
  AND2_X1 U707 ( .A1(n725), .A2(n627), .ZN(n629) );
  INV_X1 U708 ( .A(KEYINPUT108), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n631), .B(n630), .ZN(n632) );
  INV_X1 U710 ( .A(n634), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT109), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n636), .A2(n573), .ZN(n638) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n639), .A2(n358), .ZN(n669) );
  INV_X1 U716 ( .A(n423), .ZN(n640) );
  OR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n732) );
  AND2_X1 U718 ( .A1(n669), .A2(n732), .ZN(n642) );
  AND2_X2 U719 ( .A1(n643), .A2(n642), .ZN(n673) );
  INV_X1 U720 ( .A(KEYINPUT88), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  INV_X1 U722 ( .A(n673), .ZN(n651) );
  INV_X1 U723 ( .A(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n708), .A2(G475), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n657) );
  INV_X1 U726 ( .A(G952), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n716), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(G60) );
  XOR2_X1 U729 ( .A(G143), .B(KEYINPUT113), .Z(n660) );
  XNOR2_X1 U730 ( .A(n661), .B(n660), .ZN(G45) );
  NAND2_X1 U731 ( .A1(n664), .A2(n423), .ZN(n663) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(G30) );
  NAND2_X1 U734 ( .A1(n664), .A2(n725), .ZN(n665) );
  XNOR2_X1 U735 ( .A(n665), .B(G146), .ZN(G48) );
  XNOR2_X1 U736 ( .A(n666), .B(G101), .ZN(G3) );
  XOR2_X1 U737 ( .A(n667), .B(G110), .Z(G12) );
  XOR2_X1 U738 ( .A(G140), .B(KEYINPUT117), .Z(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(G42) );
  XNOR2_X1 U740 ( .A(n671), .B(n670), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(KEYINPUT125), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n674), .A2(n357), .ZN(n680) );
  XNOR2_X1 U744 ( .A(n675), .B(G227), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n676), .A2(G900), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT126), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n678), .A2(G953), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(G72) );
  XOR2_X1 U749 ( .A(G125), .B(KEYINPUT37), .Z(n681) );
  XNOR2_X1 U750 ( .A(n682), .B(n681), .ZN(G27) );
  BUF_X1 U751 ( .A(n683), .Z(n684) );
  XOR2_X1 U752 ( .A(n684), .B(G119), .Z(G21) );
  XOR2_X1 U753 ( .A(G122), .B(KEYINPUT127), .Z(n686) );
  XOR2_X1 U754 ( .A(n686), .B(n685), .Z(G24) );
  NAND2_X1 U755 ( .A1(n708), .A2(G472), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n690), .A2(n716), .ZN(n691) );
  XNOR2_X1 U758 ( .A(n691), .B(KEYINPUT63), .ZN(G57) );
  BUF_X1 U759 ( .A(n708), .Z(n692) );
  NAND2_X1 U760 ( .A1(n692), .A2(G217), .ZN(n695) );
  XOR2_X1 U761 ( .A(KEYINPUT124), .B(n693), .Z(n694) );
  XNOR2_X1 U762 ( .A(n695), .B(n694), .ZN(n696) );
  INV_X1 U763 ( .A(n716), .ZN(n699) );
  NOR2_X1 U764 ( .A1(n696), .A2(n699), .ZN(G66) );
  NAND2_X1 U765 ( .A1(n708), .A2(G478), .ZN(n697) );
  XOR2_X1 U766 ( .A(n698), .B(n697), .Z(n700) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(G63) );
  NAND2_X1 U768 ( .A1(n708), .A2(G469), .ZN(n705) );
  XNOR2_X1 U769 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT58), .ZN(n703) );
  XNOR2_X1 U771 ( .A(n705), .B(n704), .ZN(n706) );
  NAND2_X1 U772 ( .A1(n706), .A2(n716), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n707), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U774 ( .A1(n708), .A2(G210), .ZN(n715) );
  BUF_X1 U775 ( .A(n709), .Z(n713) );
  XOR2_X1 U776 ( .A(KEYINPUT55), .B(KEYINPUT93), .Z(n711) );
  XNOR2_X1 U777 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n710) );
  XOR2_X1 U778 ( .A(n711), .B(n710), .Z(n712) );
  XNOR2_X1 U779 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(KEYINPUT56), .ZN(n718) );
  XNOR2_X1 U782 ( .A(n719), .B(n718), .ZN(G51) );
  NAND2_X1 U783 ( .A1(n721), .A2(n725), .ZN(n720) );
  XNOR2_X1 U784 ( .A(n720), .B(G104), .ZN(G6) );
  XOR2_X1 U785 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n723) );
  NAND2_X1 U786 ( .A1(n721), .A2(n423), .ZN(n722) );
  XNOR2_X1 U787 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U788 ( .A(G107), .B(n724), .ZN(G9) );
  NAND2_X1 U789 ( .A1(n725), .A2(n729), .ZN(n726) );
  XNOR2_X1 U790 ( .A(n726), .B(KEYINPUT114), .ZN(n727) );
  XNOR2_X1 U791 ( .A(G113), .B(n727), .ZN(G15) );
  XOR2_X1 U792 ( .A(G116), .B(KEYINPUT115), .Z(n731) );
  NAND2_X1 U793 ( .A1(n729), .A2(n423), .ZN(n730) );
  XNOR2_X1 U794 ( .A(n731), .B(n730), .ZN(G18) );
  INV_X1 U795 ( .A(n732), .ZN(n733) );
  XOR2_X1 U796 ( .A(G134), .B(n733), .Z(n734) );
  XNOR2_X1 U797 ( .A(KEYINPUT116), .B(n734), .ZN(G36) );
  XOR2_X1 U798 ( .A(KEYINPUT87), .B(n735), .Z(n737) );
  NOR2_X1 U799 ( .A1(n737), .A2(n736), .ZN(n774) );
  NAND2_X1 U800 ( .A1(n573), .A2(n739), .ZN(n741) );
  XOR2_X1 U801 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n740) );
  XNOR2_X1 U802 ( .A(n741), .B(n740), .ZN(n749) );
  NAND2_X1 U803 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U804 ( .A(KEYINPUT49), .B(n744), .Z(n747) );
  INV_X1 U805 ( .A(n745), .ZN(n746) );
  NAND2_X1 U806 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U807 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U808 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U809 ( .A(n752), .B(KEYINPUT119), .ZN(n753) );
  XNOR2_X1 U810 ( .A(KEYINPUT51), .B(n753), .ZN(n754) );
  NOR2_X1 U811 ( .A1(n770), .A2(n754), .ZN(n765) );
  NOR2_X1 U812 ( .A1(n756), .A2(n447), .ZN(n760) );
  NOR2_X1 U813 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U814 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U815 ( .A(n761), .B(KEYINPUT120), .ZN(n763) );
  INV_X1 U816 ( .A(n762), .ZN(n769) );
  NOR2_X1 U817 ( .A1(n763), .A2(n769), .ZN(n764) );
  NOR2_X1 U818 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U819 ( .A(n766), .B(KEYINPUT52), .ZN(n767) );
  NOR2_X1 U820 ( .A1(n768), .A2(n767), .ZN(n772) );
  NOR2_X1 U821 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U822 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U824 ( .A1(n775), .A2(G953), .ZN(n776) );
  XNOR2_X1 U825 ( .A(n776), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U826 ( .A1(n777), .A2(n357), .ZN(n781) );
  NAND2_X1 U827 ( .A1(G953), .A2(G224), .ZN(n778) );
  XNOR2_X1 U828 ( .A(KEYINPUT61), .B(n778), .ZN(n779) );
  NAND2_X1 U829 ( .A1(n779), .A2(G898), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n788) );
  XOR2_X1 U831 ( .A(n783), .B(n782), .Z(n786) );
  NOR2_X1 U832 ( .A1(n357), .A2(G898), .ZN(n785) );
  NOR2_X1 U833 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U834 ( .A(n788), .B(n787), .ZN(G69) );
endmodule

