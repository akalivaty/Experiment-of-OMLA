

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U324 ( .A(n549), .B(n548), .ZN(n554) );
  NOR2_X1 U325 ( .A1(n560), .A2(n500), .ZN(n501) );
  XNOR2_X1 U326 ( .A(n503), .B(KEYINPUT47), .ZN(n504) );
  XNOR2_X1 U327 ( .A(n407), .B(n294), .ZN(n295) );
  XNOR2_X1 U328 ( .A(n296), .B(n295), .ZN(n298) );
  XNOR2_X1 U329 ( .A(n547), .B(KEYINPUT55), .ZN(n548) );
  NOR2_X1 U330 ( .A1(n545), .A2(n544), .ZN(n571) );
  XOR2_X1 U331 ( .A(n399), .B(n400), .Z(n553) );
  XNOR2_X1 U332 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n291), .B(KEYINPUT98), .ZN(n292) );
  XOR2_X1 U334 ( .A(KEYINPUT97), .B(n292), .Z(n450) );
  XOR2_X1 U335 ( .A(G57GAT), .B(KEYINPUT13), .Z(n348) );
  XNOR2_X1 U336 ( .A(G99GAT), .B(G71GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n293), .B(G120GAT), .ZN(n381) );
  XNOR2_X1 U338 ( .A(n348), .B(n381), .ZN(n296) );
  XOR2_X1 U339 ( .A(G204GAT), .B(G64GAT), .Z(n407) );
  AND2_X1 U340 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U341 ( .A(G176GAT), .B(KEYINPUT32), .Z(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n300) );
  XNOR2_X1 U344 ( .A(KEYINPUT33), .B(KEYINPUT75), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G148GAT), .Z(n304) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n417) );
  XNOR2_X1 U350 ( .A(G85GAT), .B(KEYINPUT74), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n305), .B(G92GAT), .ZN(n336) );
  XOR2_X1 U352 ( .A(n417), .B(n336), .Z(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n575) );
  XOR2_X1 U354 ( .A(G141GAT), .B(G22GAT), .Z(n426) );
  XOR2_X1 U355 ( .A(G197GAT), .B(G50GAT), .Z(n309) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G36GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(n426), .B(n310), .Z(n312) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n326) );
  XOR2_X1 U361 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U364 ( .A(KEYINPUT30), .B(G113GAT), .Z(n316) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U367 ( .A(n318), .B(n317), .Z(n324) );
  XOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT8), .Z(n320) );
  XNOR2_X1 U369 ( .A(KEYINPUT69), .B(KEYINPUT7), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n337) );
  XOR2_X1 U371 ( .A(G8GAT), .B(KEYINPUT71), .Z(n322) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n349) );
  XNOR2_X1 U374 ( .A(n337), .B(n349), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n326), .B(n325), .ZN(n550) );
  NAND2_X1 U377 ( .A1(n575), .A2(n550), .ZN(n461) );
  XOR2_X1 U378 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n328) );
  XNOR2_X1 U379 ( .A(G190GAT), .B(KEYINPUT10), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n335) );
  XOR2_X1 U381 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n330) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U384 ( .A(G50GAT), .B(G162GAT), .Z(n425) );
  XOR2_X1 U385 ( .A(n331), .B(n425), .Z(n333) );
  XNOR2_X1 U386 ( .A(G99GAT), .B(G106GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n344) );
  XOR2_X1 U389 ( .A(G36GAT), .B(KEYINPUT79), .Z(n409) );
  XOR2_X1 U390 ( .A(n336), .B(n409), .Z(n342) );
  XOR2_X1 U391 ( .A(G43GAT), .B(G134GAT), .Z(n389) );
  XOR2_X1 U392 ( .A(n337), .B(KEYINPUT9), .Z(n339) );
  NAND2_X1 U393 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n389), .B(n340), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n537) );
  INV_X1 U398 ( .A(n537), .ZN(n564) );
  XOR2_X1 U399 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n346) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(n348), .B(n347), .Z(n351) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XNOR2_X1 U404 ( .A(n349), .B(n388), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U406 ( .A(KEYINPUT14), .B(G64GAT), .Z(n353) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U409 ( .A(n355), .B(n354), .Z(n360) );
  XOR2_X1 U410 ( .A(G78GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n358), .B(KEYINPUT15), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n560) );
  INV_X1 U415 ( .A(n560), .ZN(n579) );
  NOR2_X1 U416 ( .A1(n564), .A2(n579), .ZN(n361) );
  XNOR2_X1 U417 ( .A(KEYINPUT16), .B(n361), .ZN(n448) );
  XOR2_X1 U418 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n363) );
  XNOR2_X1 U419 ( .A(G120GAT), .B(KEYINPUT5), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT90), .Z(n365) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n380) );
  XNOR2_X1 U425 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n368), .B(KEYINPUT2), .ZN(n418) );
  XOR2_X1 U427 ( .A(G113GAT), .B(KEYINPUT0), .Z(n384) );
  XOR2_X1 U428 ( .A(n418), .B(n384), .Z(n370) );
  NAND2_X1 U429 ( .A1(G225GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U431 ( .A(G85GAT), .B(G148GAT), .Z(n372) );
  XNOR2_X1 U432 ( .A(G141GAT), .B(G127GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U435 ( .A(KEYINPUT78), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U436 ( .A(G29GAT), .B(G134GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n545) );
  INV_X1 U440 ( .A(n545), .ZN(n440) );
  XOR2_X1 U441 ( .A(KEYINPUT82), .B(n381), .Z(n383) );
  NAND2_X1 U442 ( .A1(G227GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n387) );
  XNOR2_X1 U444 ( .A(KEYINPUT20), .B(KEYINPUT81), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n387), .B(n386), .Z(n391) );
  XNOR2_X1 U447 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n399) );
  XOR2_X1 U449 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n393) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U452 ( .A(n394), .B(KEYINPUT18), .Z(n396) );
  XNOR2_X1 U453 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U455 ( .A(G183GAT), .B(G176GAT), .Z(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n400) );
  INV_X1 U457 ( .A(n400), .ZN(n404) );
  XOR2_X1 U458 ( .A(KEYINPUT87), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U461 ( .A(G197GAT), .B(n403), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n404), .B(n429), .ZN(n413) );
  XOR2_X1 U463 ( .A(G92GAT), .B(KEYINPUT91), .Z(n406) );
  NAND2_X1 U464 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U466 ( .A(n408), .B(n407), .Z(n411) );
  XNOR2_X1 U467 ( .A(G8GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n540) );
  INV_X1 U470 ( .A(n540), .ZN(n487) );
  NAND2_X1 U471 ( .A1(n553), .A2(n487), .ZN(n431) );
  XOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n415) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U475 ( .A(n416), .B(KEYINPUT89), .Z(n420) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U478 ( .A(G204GAT), .B(KEYINPUT88), .Z(n422) );
  XNOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n428) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n546) );
  NAND2_X1 U485 ( .A1(n431), .A2(n546), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n432), .B(KEYINPUT95), .ZN(n433) );
  XNOR2_X1 U487 ( .A(KEYINPUT25), .B(n433), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(KEYINPUT94), .ZN(n438) );
  XOR2_X1 U489 ( .A(KEYINPUT27), .B(n540), .Z(n441) );
  NOR2_X1 U490 ( .A1(n546), .A2(n553), .ZN(n436) );
  XOR2_X1 U491 ( .A(KEYINPUT26), .B(KEYINPUT93), .Z(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n570) );
  NAND2_X1 U493 ( .A1(n441), .A2(n570), .ZN(n437) );
  NAND2_X1 U494 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND2_X1 U495 ( .A1(n440), .A2(n439), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n546), .B(KEYINPUT28), .ZN(n511) );
  INV_X1 U497 ( .A(n511), .ZN(n491) );
  NAND2_X1 U498 ( .A1(n545), .A2(n441), .ZN(n509) );
  NOR2_X1 U499 ( .A1(n491), .A2(n509), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n442), .B(KEYINPUT92), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n553), .B(KEYINPUT85), .ZN(n443) );
  NAND2_X1 U502 ( .A1(n444), .A2(n443), .ZN(n445) );
  NAND2_X1 U503 ( .A1(n446), .A2(n445), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n447), .B(KEYINPUT96), .ZN(n458) );
  NAND2_X1 U505 ( .A1(n448), .A2(n458), .ZN(n473) );
  NOR2_X1 U506 ( .A1(n461), .A2(n473), .ZN(n454) );
  NAND2_X1 U507 ( .A1(n454), .A2(n545), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(G1324GAT) );
  NAND2_X1 U509 ( .A1(n454), .A2(n487), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U511 ( .A(G15GAT), .B(KEYINPUT35), .Z(n453) );
  NAND2_X1 U512 ( .A1(n454), .A2(n553), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(G1326GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n456) );
  NAND2_X1 U515 ( .A1(n454), .A2(n491), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U517 ( .A(G22GAT), .B(n457), .ZN(G1327GAT) );
  NAND2_X1 U518 ( .A1(n458), .A2(n579), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n537), .B(KEYINPUT36), .ZN(n582) );
  NOR2_X1 U520 ( .A1(n459), .A2(n582), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT37), .ZN(n484) );
  NOR2_X1 U522 ( .A1(n461), .A2(n484), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(KEYINPUT38), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n545), .A2(n469), .ZN(n464) );
  XOR2_X1 U525 ( .A(G29GAT), .B(KEYINPUT39), .Z(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  XOR2_X1 U527 ( .A(G36GAT), .B(KEYINPUT101), .Z(n466) );
  NAND2_X1 U528 ( .A1(n487), .A2(n469), .ZN(n465) );
  XNOR2_X1 U529 ( .A(n466), .B(n465), .ZN(G1329GAT) );
  NAND2_X1 U530 ( .A1(n469), .A2(n553), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n467), .B(KEYINPUT40), .ZN(n468) );
  XNOR2_X1 U532 ( .A(G43GAT), .B(n468), .ZN(G1330GAT) );
  NAND2_X1 U533 ( .A1(n469), .A2(n491), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n470), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n471) );
  XNOR2_X1 U537 ( .A(n575), .B(n471), .ZN(n530) );
  INV_X1 U538 ( .A(n530), .ZN(n552) );
  INV_X1 U539 ( .A(n550), .ZN(n572) );
  NAND2_X1 U540 ( .A1(n552), .A2(n572), .ZN(n472) );
  XNOR2_X1 U541 ( .A(n472), .B(KEYINPUT102), .ZN(n485) );
  NOR2_X1 U542 ( .A1(n485), .A2(n473), .ZN(n480) );
  NAND2_X1 U543 ( .A1(n480), .A2(n545), .ZN(n474) );
  XNOR2_X1 U544 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U545 ( .A(G57GAT), .B(n476), .ZN(G1332GAT) );
  NAND2_X1 U546 ( .A1(n480), .A2(n487), .ZN(n477) );
  XNOR2_X1 U547 ( .A(n477), .B(KEYINPUT104), .ZN(n478) );
  XNOR2_X1 U548 ( .A(G64GAT), .B(n478), .ZN(G1333GAT) );
  NAND2_X1 U549 ( .A1(n553), .A2(n480), .ZN(n479) );
  XNOR2_X1 U550 ( .A(n479), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n482) );
  NAND2_X1 U552 ( .A1(n480), .A2(n491), .ZN(n481) );
  XNOR2_X1 U553 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U554 ( .A(G78GAT), .B(n483), .Z(G1335GAT) );
  NOR2_X1 U555 ( .A1(n485), .A2(n484), .ZN(n492) );
  NAND2_X1 U556 ( .A1(n545), .A2(n492), .ZN(n486) );
  XNOR2_X1 U557 ( .A(G85GAT), .B(n486), .ZN(G1336GAT) );
  NAND2_X1 U558 ( .A1(n492), .A2(n487), .ZN(n488) );
  XNOR2_X1 U559 ( .A(n488), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U560 ( .A1(n553), .A2(n492), .ZN(n489) );
  XNOR2_X1 U561 ( .A(n489), .B(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U562 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n494) );
  NAND2_X1 U564 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U565 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n495), .ZN(G1339GAT) );
  INV_X1 U567 ( .A(n553), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n579), .A2(n582), .ZN(n496) );
  XNOR2_X1 U569 ( .A(KEYINPUT45), .B(n496), .ZN(n497) );
  NAND2_X1 U570 ( .A1(n497), .A2(n575), .ZN(n498) );
  NOR2_X1 U571 ( .A1(n550), .A2(n498), .ZN(n507) );
  NOR2_X1 U572 ( .A1(n572), .A2(n530), .ZN(n499) );
  XNOR2_X1 U573 ( .A(n499), .B(KEYINPUT46), .ZN(n500) );
  XNOR2_X1 U574 ( .A(n501), .B(KEYINPUT108), .ZN(n502) );
  NAND2_X1 U575 ( .A1(n502), .A2(n537), .ZN(n505) );
  INV_X1 U576 ( .A(KEYINPUT109), .ZN(n503) );
  NOR2_X1 U577 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n508), .B(KEYINPUT48), .ZN(n541) );
  NOR2_X1 U579 ( .A1(n509), .A2(n541), .ZN(n510) );
  XNOR2_X1 U580 ( .A(n510), .B(KEYINPUT110), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n526), .A2(n511), .ZN(n512) );
  NOR2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n550), .A2(n522), .ZN(n514) );
  XNOR2_X1 U584 ( .A(n514), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U586 ( .A1(n522), .A2(n552), .ZN(n515) );
  XNOR2_X1 U587 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT111), .Z(n517) );
  XNOR2_X1 U589 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n520) );
  NAND2_X1 U591 ( .A1(n522), .A2(n560), .ZN(n519) );
  XNOR2_X1 U592 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U593 ( .A(G127GAT), .B(n521), .ZN(G1342GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U595 ( .A1(n522), .A2(n564), .ZN(n523) );
  XNOR2_X1 U596 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(n525), .ZN(G1343GAT) );
  NAND2_X1 U598 ( .A1(n570), .A2(n526), .ZN(n536) );
  NOR2_X1 U599 ( .A1(n572), .A2(n536), .ZN(n528) );
  XNOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n527) );
  XNOR2_X1 U601 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U602 ( .A(G141GAT), .B(n529), .ZN(G1344GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n530), .ZN(n534) );
  XOR2_X1 U604 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n532) );
  XNOR2_X1 U605 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n531) );
  XNOR2_X1 U606 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U607 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NOR2_X1 U608 ( .A1(n579), .A2(n536), .ZN(n535) );
  XOR2_X1 U609 ( .A(G155GAT), .B(n535), .Z(G1346GAT) );
  NOR2_X1 U610 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(n538), .Z(n539) );
  XNOR2_X1 U612 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  NOR2_X1 U613 ( .A1(n541), .A2(n540), .ZN(n543) );
  INV_X1 U614 ( .A(KEYINPUT54), .ZN(n542) );
  XNOR2_X1 U615 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U616 ( .A1(n571), .A2(n546), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n547) );
  AND2_X1 U618 ( .A1(n553), .A2(n554), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n565), .A2(n550), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n551), .B(G169GAT), .ZN(G1348GAT) );
  AND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n557) );
  XOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT121), .Z(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n565), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(n563), .Z(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n581) );
  NOR2_X1 U638 ( .A1(n572), .A2(n581), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(G218GAT), .B(n585), .Z(G1355GAT) );
endmodule

