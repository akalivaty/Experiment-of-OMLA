//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n253, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI21_X1  g0010(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n206), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI22_X1  g0027(.A1(new_n202), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI22_X1  g0031(.A1(new_n207), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n224), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT67), .B(G238), .Z(new_n234));
  OR2_X1    g0034(.A1(new_n234), .A2(new_n203), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n220), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(KEYINPUT1), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n218), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G13), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n220), .A2(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G257), .ZN(new_n241));
  AOI211_X1 g0041(.A(new_n223), .B(new_n240), .C1(new_n241), .C2(new_n231), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT0), .ZN(new_n244));
  AOI211_X1 g0044(.A(new_n238), .B(new_n244), .C1(new_n237), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0045(.A(G226), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G238), .B(G244), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G250), .B(G257), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G264), .B(G270), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G358));
  XNOR2_X1  g0054(.A(G68), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(new_n207), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(G58), .ZN(new_n257));
  XOR2_X1   g0057(.A(G87), .B(G97), .Z(new_n258));
  XNOR2_X1  g0058(.A(G107), .B(G116), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n257), .B(new_n260), .ZN(G351));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n212), .A2(new_n213), .A3(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n225), .A2(G1698), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n266), .B(new_n267), .C1(G226), .C2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G97), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n263), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(G238), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n274), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT13), .B1(new_n273), .B2(new_n280), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G179), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT74), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT74), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n283), .A2(new_n287), .A3(G179), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n283), .A2(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT14), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n293), .A3(G169), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n203), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n215), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n296), .B1(new_n297), .B2(new_n226), .C1(new_n299), .C2(new_n207), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n220), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n214), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n239), .A2(new_n215), .A3(G1), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT12), .ZN(new_n307));
  INV_X1    g0107(.A(new_n296), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n307), .A2(new_n239), .A3(G1), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n219), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n214), .A2(new_n301), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n203), .B1(new_n313), .B2(KEYINPUT12), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n295), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n290), .A2(G200), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n283), .A2(G190), .A3(new_n284), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n316), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G232), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n266), .B(new_n327), .C1(new_n234), .C2(new_n326), .ZN(new_n328));
  INV_X1    g0128(.A(new_n263), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(G107), .C2(new_n266), .ZN(new_n330));
  INV_X1    g0130(.A(new_n279), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n276), .A2(G274), .ZN(new_n332));
  AOI22_X1  g0132(.A1(G244), .A2(new_n331), .B1(new_n332), .B2(new_n275), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT15), .B(G87), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n297), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n339), .B1(G20), .B2(G77), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(new_n298), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n302), .B1(new_n226), .B2(new_n305), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n212), .A2(new_n213), .B1(new_n220), .B2(G33), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G77), .A3(new_n312), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n336), .B(new_n350), .C1(G179), .C2(new_n334), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n334), .A2(G200), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n330), .A2(G190), .A3(new_n333), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n349), .A3(new_n347), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n326), .A2(G222), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G223), .A2(G1698), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n266), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n329), .B(new_n358), .C1(G77), .C2(new_n266), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n331), .A2(G226), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n359), .A2(new_n277), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G179), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n361), .B2(G169), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n305), .A2(G50), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n313), .B2(G50), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n366), .A2(KEYINPUT70), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT70), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n368), .B(new_n365), .C1(new_n313), .C2(G50), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n341), .A2(new_n297), .B1(new_n371), .B2(new_n299), .ZN(new_n372));
  AOI22_X1  g0172(.A1(KEYINPUT69), .A2(new_n372), .B1(new_n208), .B2(G20), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n372), .A2(KEYINPUT69), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n348), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n355), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n318), .A2(new_n325), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n361), .A2(G190), .ZN(new_n380));
  INV_X1    g0180(.A(G200), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n361), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n366), .A2(KEYINPUT70), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n207), .B1(new_n348), .B2(new_n312), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n368), .B1(new_n385), .B2(new_n365), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n373), .A2(new_n374), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n302), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT72), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n387), .B2(new_n389), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT9), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT9), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT72), .B1(new_n370), .B2(new_n375), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n383), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT10), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT9), .B1(new_n392), .B2(new_n393), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n395), .A3(new_n391), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT10), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n383), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n379), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n341), .A2(new_n305), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n313), .B2(new_n341), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n229), .A2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n266), .B(new_n410), .C1(G223), .C2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n263), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n277), .B1(new_n225), .B2(new_n279), .ZN(new_n414));
  AND2_X1   g0214(.A1(KEYINPUT77), .A2(G190), .ZN(new_n415));
  NOR2_X1   g0215(.A1(KEYINPUT77), .A2(G190), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n413), .A2(new_n414), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(G200), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n264), .A2(new_n215), .A3(new_n265), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n265), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n203), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G58), .A2(G68), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n204), .A2(new_n205), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n298), .A2(G159), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n348), .B1(new_n432), .B2(KEYINPUT16), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT16), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n426), .B2(new_n431), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT75), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g0236(.A1(KEYINPUT3), .A2(G33), .ZN(new_n437));
  NOR2_X1   g0237(.A1(KEYINPUT3), .A2(G33), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT7), .B1(new_n439), .B2(new_n215), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n437), .A2(new_n438), .A3(new_n423), .A4(G20), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n428), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT16), .A3(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n435), .A2(new_n444), .A3(KEYINPUT75), .A4(new_n302), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n409), .B(new_n421), .C1(new_n436), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g0251(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n452));
  NAND3_X1  g0252(.A1(new_n435), .A2(new_n444), .A3(new_n302), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT75), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n408), .B1(new_n455), .B2(new_n445), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n452), .B1(new_n456), .B2(new_n421), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n409), .B1(new_n436), .B2(new_n446), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n420), .A2(G179), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n335), .B2(new_n420), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n462), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n456), .A2(KEYINPUT18), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT76), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n460), .A2(new_n459), .A3(new_n462), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT18), .B1(new_n456), .B2(new_n464), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT76), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n458), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n405), .A2(new_n406), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n295), .A2(new_n317), .B1(new_n323), .B2(new_n324), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n403), .B1(new_n402), .B2(new_n383), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT10), .B(new_n382), .C1(new_n400), .C2(new_n401), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n378), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n456), .B(new_n421), .C1(new_n448), .C2(new_n449), .ZN(new_n477));
  INV_X1    g0277(.A(new_n447), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(new_n452), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n469), .B1(new_n467), .B2(new_n468), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT79), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n219), .B(G45), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(new_n276), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT82), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n487), .B(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n276), .A2(G274), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n490), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n223), .B1(new_n264), .B2(new_n265), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g0300(.A(G1698), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n439), .B2(new_n227), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G283), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n500), .A2(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n266), .A2(G244), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n485), .B(new_n498), .C1(new_n506), .C2(new_n329), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n505), .A3(new_n503), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n266), .A2(G250), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n326), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n329), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n498), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT83), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n335), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n305), .A2(new_n270), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n515), .B(KEYINPUT81), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n305), .B1(new_n219), .B2(G33), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n517), .A2(new_n348), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(G97), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n298), .A2(G77), .ZN(new_n520));
  XNOR2_X1  g0320(.A(new_n520), .B(KEYINPUT80), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n522), .A2(new_n270), .A3(G107), .ZN(new_n523));
  XNOR2_X1  g0323(.A(G97), .B(G107), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n521), .B1(new_n215), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n230), .B1(new_n424), .B2(new_n425), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n302), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n498), .B1(new_n506), .B2(new_n329), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n519), .A2(new_n528), .B1(new_n529), .B2(new_n362), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n514), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  INV_X1    g0333(.A(G190), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n507), .A2(new_n513), .A3(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n519), .B(new_n528), .C1(new_n529), .C2(new_n381), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n513), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n529), .A2(KEYINPUT83), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(G190), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n536), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT84), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n532), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G116), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n305), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n517), .A2(G116), .A3(new_n348), .ZN(new_n546));
  AOI21_X1  g0346(.A(G20), .B1(new_n269), .B2(G97), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n503), .B1(G20), .B2(new_n544), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n302), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n302), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n545), .B(new_n546), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G264), .A2(G1698), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n266), .B(new_n552), .C1(new_n241), .C2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G303), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n439), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n329), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n487), .B(KEYINPUT82), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(new_n332), .A3(new_n494), .A4(new_n496), .ZN(new_n558));
  OAI211_X1 g0358(.A(G270), .B(new_n276), .C1(new_n488), .C2(new_n489), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n551), .A2(KEYINPUT21), .A3(G169), .A4(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n558), .A3(G179), .A4(new_n559), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n551), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(G169), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT21), .B1(new_n567), .B2(new_n551), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n417), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n560), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n551), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n560), .A2(G200), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(KEYINPUT88), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n572), .B2(new_n566), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(new_n574), .A3(new_n564), .A4(new_n561), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT88), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n495), .A2(G1), .A3(G274), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n223), .B1(new_n495), .B2(G1), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n276), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G238), .A2(G1698), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n227), .B2(G1698), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(new_n266), .B1(G33), .B2(G116), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n362), .B(new_n584), .C1(new_n587), .C2(new_n263), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n588), .A2(KEYINPUT85), .ZN(new_n589));
  AOI21_X1  g0389(.A(G20), .B1(new_n271), .B2(KEYINPUT19), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n222), .A2(new_n270), .A3(new_n230), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n222), .A2(new_n270), .A3(new_n230), .A4(KEYINPUT86), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n266), .A2(new_n215), .A3(G68), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n297), .B2(new_n270), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n302), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n337), .A2(new_n305), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n517), .A2(new_n348), .A3(new_n338), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n588), .A2(KEYINPUT85), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n586), .A2(new_n266), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G116), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n263), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n584), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n335), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n589), .A2(new_n603), .A3(new_n604), .A4(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n593), .A2(new_n594), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n596), .B(new_n598), .C1(new_n611), .C2(new_n590), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(new_n302), .B1(new_n305), .B2(new_n337), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n518), .A2(G87), .ZN(new_n614));
  OAI211_X1 g0414(.A(G190), .B(new_n584), .C1(new_n587), .C2(new_n263), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n584), .B1(new_n587), .B2(new_n263), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n610), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n241), .A2(new_n326), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n266), .A2(new_n621), .B1(G33), .B2(G294), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n499), .A2(new_n326), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n329), .ZN(new_n625));
  OAI211_X1 g0425(.A(G264), .B(new_n276), .C1(new_n488), .C2(new_n489), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n558), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G169), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(KEYINPUT90), .A3(G169), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n627), .A2(new_n362), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n266), .A2(new_n215), .A3(G87), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT22), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT22), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n266), .A2(new_n636), .A3(new_n215), .A4(G87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT24), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n215), .B2(G107), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT23), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT23), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(G116), .B2(new_n339), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n639), .B1(new_n638), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n302), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n305), .A2(new_n230), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT25), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(G107), .B2(new_n518), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n633), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n610), .A2(new_n618), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT87), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n627), .A2(new_n534), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n627), .A2(G200), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n655), .A2(new_n647), .A3(new_n650), .A4(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n620), .A2(new_n652), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  AND4_X1   g0458(.A1(new_n484), .A2(new_n543), .A3(new_n581), .A4(new_n658), .ZN(G372));
  AND3_X1   g0459(.A1(new_n614), .A2(new_n601), .A3(new_n600), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n617), .A2(new_n615), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n609), .A2(new_n588), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n660), .A2(new_n661), .B1(new_n662), .B2(new_n603), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n514), .A3(new_n664), .A4(new_n530), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n603), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n532), .A2(new_n654), .A3(new_n620), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n537), .A2(new_n542), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n652), .A2(new_n569), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n657), .A2(new_n663), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n671), .A3(new_n531), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n484), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n474), .B2(new_n475), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n399), .A2(KEYINPUT91), .A3(new_n404), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n463), .A2(new_n465), .ZN(new_n680));
  INV_X1    g0480(.A(new_n351), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n325), .A2(new_n681), .B1(new_n317), .B2(new_n295), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n682), .B2(new_n458), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n377), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n219), .A2(new_n215), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g0489(.A(KEYINPUT92), .B(G343), .Z(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n572), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n565), .B2(new_n568), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n581), .B(KEYINPUT93), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n652), .A2(new_n657), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n651), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n692), .ZN(new_n701));
  INV_X1    g0501(.A(new_n652), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n691), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n697), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n569), .A2(new_n691), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n652), .B2(new_n691), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(G399));
  NAND2_X1  g0511(.A1(new_n611), .A2(new_n544), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n240), .A2(G41), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n219), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n217), .B2(new_n713), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  AOI21_X1  g0516(.A(new_n691), .B1(new_n669), .B2(new_n673), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  OR3_X1    g0518(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT29), .ZN(new_n719));
  INV_X1    g0519(.A(new_n666), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n532), .A2(new_n663), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(KEYINPUT26), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n532), .A2(new_n654), .A3(new_n664), .A4(new_n620), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n691), .B1(new_n724), .B2(new_n673), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n718), .B1(new_n717), .B2(KEYINPUT29), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n719), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n658), .A2(new_n581), .A3(new_n543), .A4(new_n692), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n616), .A2(new_n362), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(new_n627), .A3(new_n560), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n529), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n625), .A2(new_n626), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n562), .A3(new_n616), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n538), .A3(new_n539), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n734), .A2(new_n538), .A3(KEYINPUT30), .A4(new_n539), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n691), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n692), .B1(new_n737), .B2(new_n738), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT31), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n729), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n728), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT95), .Z(new_n748));
  OAI21_X1  g0548(.A(new_n716), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n239), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n219), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n713), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n696), .B2(G330), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n696), .ZN(new_n755));
  INV_X1    g0555(.A(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n240), .A2(new_n266), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n217), .B2(new_n495), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(new_n257), .B2(new_n495), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n240), .A2(new_n439), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(G355), .B1(new_n544), .B2(new_n240), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n766));
  OR3_X1    g0566(.A1(KEYINPUT98), .A2(G13), .A3(G33), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT98), .B1(G13), .B2(G33), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n214), .B1(G20), .B2(new_n335), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n765), .A2(new_n766), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n215), .A2(G179), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n779), .A2(G329), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n215), .A2(new_n362), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n570), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n266), .B(new_n780), .C1(G326), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n781), .B(KEYINPUT99), .Z(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(new_n777), .ZN(new_n787));
  INV_X1    g0587(.A(G322), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n570), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n784), .B1(new_n785), .B2(new_n787), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n782), .A2(G190), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n776), .A2(new_n534), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n795), .B2(G283), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n534), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n215), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n796), .B1(new_n797), .B2(new_n799), .C1(new_n554), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n792), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n203), .B1(new_n799), .B2(new_n270), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n800), .A2(new_n222), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n439), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n783), .A2(G50), .B1(G107), .B2(new_n795), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n804), .A2(new_n805), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G159), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n778), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT32), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n787), .B2(new_n226), .C1(new_n202), .C2(new_n790), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n791), .A2(new_n801), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n756), .B(new_n775), .C1(new_n772), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n771), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n696), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n755), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n351), .A2(new_n691), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n350), .A2(new_n691), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n354), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n351), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n717), .B(new_n826), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(new_n746), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n753), .B1(new_n827), .B2(new_n746), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n772), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n770), .ZN(new_n832));
  INV_X1    g0632(.A(new_n800), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G107), .B1(new_n795), .B2(G87), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  INV_X1    g0635(.A(new_n783), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n802), .C1(new_n836), .C2(new_n554), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n266), .B1(new_n779), .B2(G311), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n270), .B2(new_n799), .C1(new_n787), .C2(new_n544), .ZN(new_n839));
  INV_X1    g0639(.A(new_n790), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n837), .B(new_n839), .C1(G294), .C2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n783), .A2(G137), .B1(G150), .B2(new_n792), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n787), .B2(new_n810), .C1(new_n843), .C2(new_n790), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n266), .B1(new_n778), .B2(new_n846), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n799), .A2(new_n202), .B1(new_n794), .B2(new_n203), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G50), .C2(new_n833), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n841), .B1(new_n845), .B2(new_n849), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n753), .B1(G77), .B2(new_n832), .C1(new_n850), .C2(new_n831), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n769), .B2(new_n825), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT101), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n830), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G384));
  INV_X1    g0655(.A(new_n525), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n216), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  NAND3_X1  g0660(.A1(new_n217), .A2(G77), .A3(new_n427), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n207), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n219), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n460), .A2(new_n462), .ZN(new_n866));
  INV_X1    g0666(.A(new_n689), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n460), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n866), .A2(new_n868), .A3(new_n869), .A4(new_n447), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n444), .A2(new_n302), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n442), .A2(new_n443), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT103), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT16), .B1(new_n872), .B2(KEYINPUT103), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n875), .A2(new_n408), .B1(new_n462), .B2(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n447), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n865), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n875), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n689), .B1(new_n880), .B2(new_n409), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n879), .B1(new_n471), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n870), .A2(new_n878), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n482), .B2(new_n881), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n447), .B1(new_n456), .B2(new_n464), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n456), .A2(new_n689), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n890), .A2(new_n870), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n868), .B1(new_n680), .B2(new_n479), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n865), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n883), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT104), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n893), .A2(new_n883), .A3(new_n897), .A4(new_n894), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n887), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n318), .A2(new_n691), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n680), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n689), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n870), .A2(new_n878), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n471), .B2(new_n882), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n482), .A2(new_n881), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n905), .A2(new_n865), .B1(new_n906), .B2(new_n879), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n318), .A2(new_n325), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n316), .A2(new_n692), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n318), .B(new_n325), .C1(new_n316), .C2(new_n692), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n691), .B(new_n825), .C1(new_n669), .C2(new_n673), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n820), .B(KEYINPUT102), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n903), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT105), .B1(new_n901), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n919), .B(new_n916), .C1(new_n899), .C2(new_n900), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n484), .A2(new_n719), .A3(new_n726), .A4(new_n727), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n684), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT106), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n740), .A2(new_n926), .A3(new_n741), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT106), .B1(new_n743), .B2(KEYINPUT31), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n729), .A2(new_n927), .A3(new_n744), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n825), .B1(new_n910), .B2(new_n911), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n925), .B1(new_n907), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n893), .A2(new_n883), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n929), .A4(new_n930), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n934), .A3(G330), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n484), .A2(G330), .A3(new_n929), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n932), .A2(new_n934), .A3(new_n484), .A4(new_n929), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n924), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n219), .B2(new_n750), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n924), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n864), .B1(new_n943), .B2(new_n944), .ZN(G367));
  INV_X1    g0745(.A(new_n240), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n773), .B1(new_n946), .B2(new_n337), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n253), .A2(new_n757), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n753), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT46), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n833), .A2(G116), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n840), .A2(G303), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n835), .B2(new_n787), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n783), .A2(G311), .B1(G294), .B2(new_n792), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n270), .B2(new_n794), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n266), .B1(new_n779), .B2(G317), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n956), .B1(new_n230), .B2(new_n799), .C1(new_n951), .C2(new_n950), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n953), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n792), .A2(G159), .B1(new_n795), .B2(G77), .ZN(new_n959));
  INV_X1    g0759(.A(new_n799), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(G68), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(new_n836), .C2(new_n843), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n439), .B1(new_n779), .B2(G137), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n202), .B2(new_n800), .C1(new_n787), .C2(new_n207), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n962), .B(new_n964), .C1(G150), .C2(new_n840), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  AOI21_X1  g0767(.A(new_n949), .B1(new_n967), .B2(new_n772), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n660), .A2(new_n692), .ZN(new_n969));
  MUX2_X1   g0769(.A(new_n663), .B(new_n720), .S(new_n969), .Z(new_n970));
  OAI21_X1  g0770(.A(new_n968), .B1(new_n816), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n519), .A2(new_n528), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n543), .B1(new_n972), .B2(new_n692), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n532), .A2(new_n691), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n710), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT45), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n709), .A2(new_n973), .A3(new_n974), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT44), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n977), .A2(new_n705), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n705), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n984));
  INV_X1    g0784(.A(new_n704), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n984), .C1(new_n985), .C2(new_n707), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n697), .B(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n748), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT108), .B(KEYINPUT41), .Z(new_n989));
  XOR2_X1   g0789(.A(new_n713), .B(new_n989), .Z(new_n990));
  AOI21_X1  g0790(.A(new_n752), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n975), .A2(new_n699), .A3(new_n707), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n992), .A2(KEYINPUT42), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n531), .B1(new_n973), .B2(new_n652), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n992), .A2(KEYINPUT42), .B1(new_n994), .B2(new_n692), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n993), .A2(new_n995), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n996), .B(new_n997), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n705), .A2(new_n975), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n971), .B1(new_n991), .B2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n987), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n748), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n713), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT112), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT112), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1006), .A3(new_n713), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(new_n748), .C2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n704), .A2(new_n771), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n762), .A2(new_n712), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(G107), .B2(new_n946), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n712), .C1(G68), .C2(G77), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT110), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT110), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n341), .A2(G50), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT50), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n758), .B1(new_n250), .B2(G45), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n753), .B1(new_n1020), .B2(new_n774), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n836), .A2(new_n810), .B1(new_n226), .B2(new_n800), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n960), .A2(new_n338), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n802), .B2(new_n341), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n266), .B1(new_n778), .B2(new_n371), .C1(new_n270), .C2(new_n794), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n840), .B2(G50), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(new_n203), .C2(new_n787), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n266), .B1(new_n779), .B2(G326), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n799), .A2(new_n835), .B1(new_n800), .B2(new_n797), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT111), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n783), .A2(G322), .B1(G311), .B2(new_n792), .ZN(new_n1032));
  INV_X1    g0832(.A(G317), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n787), .B2(new_n554), .C1(new_n1033), .C2(new_n790), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT49), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1029), .B1(new_n544), .B2(new_n794), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1028), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1021), .B1(new_n1041), .B2(new_n772), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1002), .A2(new_n752), .B1(new_n1009), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1008), .A2(new_n1043), .ZN(G393));
  OAI22_X1  g0844(.A1(new_n790), .A2(new_n810), .B1(new_n836), .B2(new_n371), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n802), .A2(new_n207), .B1(new_n799), .B2(new_n226), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G68), .B2(new_n833), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n266), .B1(new_n778), .B2(new_n843), .C1(new_n222), .C2(new_n794), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n787), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n342), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1046), .A2(new_n1048), .A3(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n439), .B1(new_n778), .B2(new_n788), .C1(new_n230), .C2(new_n794), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G116), .A2(new_n960), .B1(new_n792), .B2(G303), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n835), .B2(new_n800), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(G294), .C2(new_n1050), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n790), .A2(new_n785), .B1(new_n836), .B2(new_n1033), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n831), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n260), .A2(new_n758), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n774), .B1(G97), .B2(new_n240), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n756), .B(new_n1060), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n975), .B2(new_n816), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n713), .B1(new_n1003), .B2(new_n982), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n982), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n748), .B2(new_n1002), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1064), .B1(new_n751), .B2(new_n982), .C1(new_n1065), .C2(new_n1067), .ZN(G390));
  AND2_X1   g0868(.A1(new_n826), .A2(G330), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n929), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n912), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n820), .B1(new_n725), .B2(new_n824), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n745), .A2(new_n912), .A3(new_n1069), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n914), .B1(new_n717), .B2(new_n826), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n745), .A2(new_n1069), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n1071), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n929), .A2(new_n912), .A3(new_n1069), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n922), .A2(new_n684), .A3(new_n936), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n900), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1076), .B2(new_n1071), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n887), .A2(new_n896), .A3(new_n898), .A4(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n933), .C1(new_n1073), .C2(new_n1071), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1086), .A2(new_n1087), .A3(new_n1074), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1079), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1079), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1086), .A2(new_n1087), .A3(new_n1074), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1090), .A2(new_n713), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT113), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1090), .A2(KEYINPUT113), .A3(new_n713), .A4(new_n1096), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(KEYINPUT39), .A2(new_n886), .B1(new_n895), .B2(KEYINPUT104), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n769), .A3(new_n898), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n753), .B1(new_n832), .B2(new_n342), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT114), .ZN(new_n1105));
  INV_X1    g0905(.A(G137), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n802), .A2(new_n1106), .B1(new_n799), .B2(new_n810), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G50), .B2(new_n795), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n779), .A2(G125), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n439), .B(new_n1109), .C1(G128), .C2(new_n783), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT53), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n800), .A2(new_n371), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1108), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT115), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1050), .A2(new_n1115), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n846), .B2(new_n790), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n960), .A2(G77), .B1(new_n795), .B2(G68), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n230), .B2(new_n802), .C1(new_n836), .C2(new_n835), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n266), .B(new_n806), .C1(G294), .C2(new_n779), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n270), .B2(new_n787), .C1(new_n544), .C2(new_n790), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1113), .A2(new_n1117), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1105), .B1(new_n1122), .B2(new_n772), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1101), .A2(new_n752), .B1(new_n1103), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1099), .A2(new_n1100), .A3(new_n1124), .ZN(G378));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1084), .B1(new_n1102), .B2(new_n898), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n919), .B1(new_n1127), .B2(new_n916), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n901), .A2(KEYINPUT105), .A3(new_n917), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n377), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n679), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n689), .B1(new_n396), .B2(new_n391), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1132), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n679), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1134), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1135), .B1(new_n679), .B2(new_n1130), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n377), .B(new_n1132), .C1(new_n677), .C2(new_n678), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(G330), .A3(new_n932), .A4(new_n934), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n935), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1128), .A2(new_n1129), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1143), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n918), .B2(new_n920), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT118), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1082), .B(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1126), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1082), .B(KEYINPUT118), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1096), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(KEYINPUT57), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n713), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1146), .A2(new_n1148), .A3(new_n752), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n753), .B1(new_n832), .B2(G50), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G41), .B(new_n266), .C1(new_n779), .C2(G283), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n202), .B2(new_n794), .C1(new_n226), .C2(new_n800), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT116), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n961), .B1(new_n270), .B2(new_n802), .C1(new_n836), .C2(new_n544), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n790), .A2(new_n230), .B1(new_n787), .B2(new_n337), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT58), .Z(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n269), .B2(new_n486), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n266), .B2(G41), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n790), .A2(new_n1169), .B1(new_n787), .B2(new_n1106), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n783), .A2(G125), .B1(G150), .B2(new_n960), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n846), .B2(new_n802), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n833), .C2(new_n1115), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n795), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n779), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1166), .B(new_n1168), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT117), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n831), .B1(new_n1180), .B2(KEYINPUT117), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1159), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1142), .B2(new_n770), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1158), .A2(new_n1184), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1157), .A2(KEYINPUT119), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT119), .B1(new_n1157), .B2(new_n1185), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(G375));
  INV_X1    g0988(.A(new_n1081), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1071), .A2(new_n769), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n753), .B1(new_n832), .B2(G68), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n266), .B1(new_n795), .B2(G77), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n790), .B2(new_n835), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1023), .B1(new_n544), .B2(new_n802), .C1(new_n836), .C2(new_n797), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n800), .A2(new_n270), .B1(new_n778), .B2(new_n554), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(KEYINPUT120), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(KEYINPUT120), .B2(new_n1195), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1193), .B(new_n1197), .C1(G107), .C2(new_n1050), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n836), .A2(new_n846), .B1(new_n810), .B2(new_n800), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G50), .B2(new_n960), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n266), .B1(new_n778), .B2(new_n1169), .C1(new_n202), .C2(new_n794), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n840), .B2(G137), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1050), .A2(G150), .B1(new_n792), .B2(new_n1115), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1199), .A2(KEYINPUT121), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1200), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1191), .B1(new_n1208), .B2(new_n772), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1189), .A2(new_n752), .B1(new_n1190), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1083), .A2(new_n990), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT122), .Z(G381));
  NAND3_X1  g1014(.A1(new_n1008), .A2(new_n818), .A3(new_n1043), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1097), .A2(new_n1124), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(G381), .A2(new_n1215), .A3(G384), .A4(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(G390), .A2(G387), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(new_n1187), .C2(new_n1186), .ZN(G407));
  INV_X1    g1019(.A(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n690), .A2(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n1186), .C2(new_n1187), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(G213), .A3(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT123), .ZN(G409));
  NAND3_X1  g1025(.A1(new_n1157), .A2(G378), .A3(new_n1185), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1155), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n990), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1158), .A2(new_n1184), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1220), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1081), .A2(KEYINPUT60), .A3(new_n1082), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1083), .A2(new_n713), .A3(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1212), .A2(KEYINPUT60), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1210), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(new_n854), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n854), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1232), .A2(new_n1221), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1232), .A2(new_n1245), .A3(new_n1221), .A4(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1222), .A2(G2897), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1237), .A2(new_n1238), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n713), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1227), .B2(new_n1126), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1230), .B1(new_n1252), .B2(new_n1156), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1185), .B1(new_n1228), .B2(new_n1227), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1253), .A2(G378), .B1(new_n1254), .B2(new_n1220), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1250), .B1(new_n1255), .B2(new_n1222), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1232), .A2(new_n1221), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1250), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1260), .A2(new_n1243), .A3(new_n1261), .A4(new_n1246), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  AND2_X1   g1063(.A1(G390), .A2(G387), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1215), .C1(new_n1264), .C2(new_n1218), .ZN(new_n1265));
  OR2_X1    g1065(.A1(G390), .A2(G387), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G390), .A2(G387), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1008), .A2(new_n818), .A3(new_n1043), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n818), .B1(new_n1008), .B2(new_n1043), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1266), .B(new_n1267), .C1(new_n1268), .C2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1258), .A2(new_n1262), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1241), .A2(new_n1274), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1275), .A2(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(KEYINPUT63), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1260), .A3(new_n1271), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1278), .ZN(G405));
  NOR3_X1   g1079(.A1(new_n1186), .A2(new_n1187), .A3(new_n1216), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1226), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1239), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1187), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1253), .A2(KEYINPUT119), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1220), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1226), .A3(new_n1240), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1282), .A2(new_n1271), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1282), .A2(new_n1271), .A3(new_n1286), .A4(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1272), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .ZN(G402));
endmodule


