

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  XNOR2_X1 U323 ( .A(n546), .B(KEYINPUT54), .ZN(n547) );
  XNOR2_X1 U324 ( .A(n548), .B(n547), .ZN(n570) );
  XNOR2_X1 U325 ( .A(n363), .B(n421), .ZN(n364) );
  XOR2_X1 U326 ( .A(KEYINPUT36), .B(n464), .Z(n586) );
  XNOR2_X1 U327 ( .A(n365), .B(n364), .ZN(n371) );
  NOR2_X1 U328 ( .A1(n555), .A2(n554), .ZN(n565) );
  XNOR2_X1 U329 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n457) );
  XOR2_X1 U330 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n292) );
  XNOR2_X1 U331 ( .A(KEYINPUT1), .B(KEYINPUT95), .ZN(n291) );
  XNOR2_X1 U332 ( .A(n292), .B(n291), .ZN(n312) );
  XOR2_X1 U333 ( .A(G155GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U334 ( .A(G29GAT), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U336 ( .A(KEYINPUT6), .B(G57GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U339 ( .A(n298), .B(n297), .Z(n310) );
  XOR2_X1 U340 ( .A(KEYINPUT2), .B(KEYINPUT94), .Z(n300) );
  XNOR2_X1 U341 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n427) );
  XOR2_X1 U343 ( .A(n427), .B(KEYINPUT5), .Z(n302) );
  NAND2_X1 U344 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n308) );
  XOR2_X1 U346 ( .A(G134GAT), .B(KEYINPUT79), .Z(n352) );
  XOR2_X1 U347 ( .A(n352), .B(G85GAT), .Z(n306) );
  XOR2_X1 U348 ( .A(G127GAT), .B(KEYINPUT0), .Z(n304) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n407) );
  XNOR2_X1 U351 ( .A(n407), .B(G162GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U355 ( .A(n312), .B(n311), .Z(n514) );
  XOR2_X1 U356 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n314) );
  XNOR2_X1 U357 ( .A(G92GAT), .B(KEYINPUT32), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U359 ( .A(KEYINPUT75), .B(KEYINPUT72), .Z(n316) );
  NAND2_X1 U360 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U362 ( .A(n317), .B(KEYINPUT31), .Z(n323) );
  XOR2_X1 U363 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U364 ( .A(KEYINPUT73), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n439) );
  XOR2_X1 U366 ( .A(KEYINPUT74), .B(G85GAT), .Z(n321) );
  XNOR2_X1 U367 ( .A(G99GAT), .B(G106GAT), .ZN(n320) );
  XNOR2_X1 U368 ( .A(n321), .B(n320), .ZN(n361) );
  XNOR2_X1 U369 ( .A(n439), .B(n361), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n325) );
  XNOR2_X1 U371 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n324), .B(KEYINPUT13), .ZN(n384) );
  XOR2_X1 U373 ( .A(n325), .B(n384), .Z(n327) );
  XOR2_X1 U374 ( .A(G120GAT), .B(G71GAT), .Z(n396) );
  XOR2_X1 U375 ( .A(G176GAT), .B(G64GAT), .Z(n414) );
  XNOR2_X1 U376 ( .A(n396), .B(n414), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n577) );
  XOR2_X1 U379 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n331) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G29GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U382 ( .A(KEYINPUT7), .B(n332), .ZN(n366) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n334) );
  XNOR2_X1 U384 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U386 ( .A(G22GAT), .B(G197GAT), .Z(n336) );
  XNOR2_X1 U387 ( .A(G50GAT), .B(G36GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U389 ( .A(G8GAT), .B(G113GAT), .Z(n338) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G141GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n381) );
  XOR2_X1 U394 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n342) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n381), .B(n343), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U399 ( .A(n347), .B(n346), .Z(n348) );
  XOR2_X1 U400 ( .A(n366), .B(n348), .Z(n479) );
  INV_X1 U401 ( .A(n479), .ZN(n573) );
  NAND2_X1 U402 ( .A1(n577), .A2(n573), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n349), .B(KEYINPUT76), .ZN(n469) );
  XOR2_X1 U404 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n351) );
  XNOR2_X1 U405 ( .A(KEYINPUT64), .B(KEYINPUT11), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n353), .B(n352), .ZN(n355) );
  AND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n358) );
  INV_X1 U410 ( .A(n358), .ZN(n357) );
  INV_X1 U411 ( .A(KEYINPUT80), .ZN(n356) );
  NAND2_X1 U412 ( .A1(n357), .A2(n356), .ZN(n360) );
  NAND2_X1 U413 ( .A1(n358), .A2(KEYINPUT80), .ZN(n359) );
  NAND2_X1 U414 ( .A1(n360), .A2(n359), .ZN(n365) );
  XNOR2_X1 U415 ( .A(n361), .B(KEYINPUT78), .ZN(n363) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n362), .B(G92GAT), .ZN(n421) );
  INV_X1 U418 ( .A(n366), .ZN(n369) );
  XOR2_X1 U419 ( .A(G162GAT), .B(KEYINPUT77), .Z(n368) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n432) );
  XNOR2_X1 U422 ( .A(n369), .B(n432), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n371), .B(n370), .ZN(n541) );
  INV_X1 U424 ( .A(KEYINPUT81), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n541), .B(n372), .ZN(n464) );
  XOR2_X1 U426 ( .A(KEYINPUT86), .B(KEYINPUT15), .Z(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n373) );
  XNOR2_X1 U428 ( .A(n374), .B(n373), .ZN(n391) );
  XOR2_X1 U429 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n376) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT14), .B(n377), .ZN(n389) );
  XOR2_X1 U433 ( .A(KEYINPUT85), .B(G64GAT), .Z(n379) );
  XNOR2_X1 U434 ( .A(G211GAT), .B(G78GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U436 ( .A(n380), .B(G71GAT), .Z(n383) );
  XNOR2_X1 U437 ( .A(n381), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U439 ( .A(n385), .B(n384), .Z(n387) );
  XOR2_X1 U440 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U441 ( .A(G8GAT), .B(G183GAT), .Z(n417) );
  XNOR2_X1 U442 ( .A(n428), .B(n417), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n526) );
  NOR2_X1 U446 ( .A1(n464), .A2(n526), .ZN(n392) );
  XNOR2_X1 U447 ( .A(KEYINPUT16), .B(n392), .ZN(n454) );
  INV_X1 U448 ( .A(n514), .ZN(n569) );
  XOR2_X1 U449 ( .A(G190GAT), .B(G134GAT), .Z(n394) );
  XNOR2_X1 U450 ( .A(G43GAT), .B(G99GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U453 ( .A1(G227GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n411) );
  XOR2_X1 U455 ( .A(G183GAT), .B(KEYINPUT89), .Z(n400) );
  XNOR2_X1 U456 ( .A(G176GAT), .B(KEYINPUT91), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U458 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n402) );
  XNOR2_X1 U459 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n406) );
  XNOR2_X1 U463 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n413), .B(n407), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n555) );
  INV_X1 U468 ( .A(n555), .ZN(n519) );
  XNOR2_X1 U469 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n412), .B(G211GAT), .ZN(n440) );
  XNOR2_X1 U471 ( .A(n413), .B(n440), .ZN(n425) );
  XNOR2_X1 U472 ( .A(G204GAT), .B(G218GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U474 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U475 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U477 ( .A(n420), .B(KEYINPUT98), .Z(n423) );
  XNOR2_X1 U478 ( .A(n421), .B(KEYINPUT99), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n544) );
  XOR2_X1 U481 ( .A(n544), .B(KEYINPUT100), .Z(n426) );
  XNOR2_X1 U482 ( .A(KEYINPUT27), .B(n426), .ZN(n516) );
  NOR2_X1 U483 ( .A1(n519), .A2(n516), .ZN(n443) );
  XOR2_X1 U484 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U487 ( .A(n431), .B(KEYINPUT24), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(KEYINPUT22), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n436) );
  XNOR2_X1 U491 ( .A(G106GAT), .B(KEYINPUT23), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n549) );
  XNOR2_X1 U496 ( .A(n549), .B(KEYINPUT28), .ZN(n518) );
  NAND2_X1 U497 ( .A1(n443), .A2(n518), .ZN(n444) );
  NOR2_X1 U498 ( .A1(n569), .A2(n444), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n445), .B(KEYINPUT101), .ZN(n453) );
  NAND2_X1 U500 ( .A1(n544), .A2(n519), .ZN(n446) );
  NAND2_X1 U501 ( .A1(n549), .A2(n446), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT25), .B(n447), .Z(n450) );
  NOR2_X1 U503 ( .A1(n549), .A2(n519), .ZN(n448) );
  XOR2_X1 U504 ( .A(KEYINPUT26), .B(n448), .Z(n568) );
  OR2_X1 U505 ( .A1(n568), .A2(n516), .ZN(n449) );
  NAND2_X1 U506 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n569), .A2(n451), .ZN(n452) );
  NAND2_X1 U508 ( .A1(n453), .A2(n452), .ZN(n465) );
  NAND2_X1 U509 ( .A1(n454), .A2(n465), .ZN(n455) );
  XNOR2_X1 U510 ( .A(n455), .B(KEYINPUT102), .ZN(n480) );
  NOR2_X1 U511 ( .A1(n469), .A2(n480), .ZN(n461) );
  NAND2_X1 U512 ( .A1(n514), .A2(n461), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(G1324GAT) );
  NAND2_X1 U514 ( .A1(n461), .A2(n544), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U516 ( .A(G15GAT), .B(KEYINPUT35), .Z(n460) );
  NAND2_X1 U517 ( .A1(n461), .A2(n519), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(G1326GAT) );
  XOR2_X1 U519 ( .A(G22GAT), .B(KEYINPUT103), .Z(n463) );
  INV_X1 U520 ( .A(n518), .ZN(n496) );
  NAND2_X1 U521 ( .A1(n461), .A2(n496), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(G1327GAT) );
  NAND2_X1 U523 ( .A1(n526), .A2(n465), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n586), .A2(n466), .ZN(n468) );
  XNOR2_X1 U525 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n468), .B(n467), .ZN(n492) );
  NOR2_X1 U527 ( .A1(n469), .A2(n492), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT38), .ZN(n477) );
  NAND2_X1 U529 ( .A1(n477), .A2(n514), .ZN(n473) );
  XNOR2_X1 U530 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT39), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(G1328GAT) );
  NAND2_X1 U533 ( .A1(n477), .A2(n544), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U535 ( .A1(n477), .A2(n519), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n475), .B(KEYINPUT40), .ZN(n476) );
  XNOR2_X1 U537 ( .A(G43GAT), .B(n476), .ZN(G1330GAT) );
  NAND2_X1 U538 ( .A1(n496), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G50GAT), .B(n478), .ZN(G1331GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n482) );
  XNOR2_X1 U541 ( .A(KEYINPUT41), .B(n577), .ZN(n561) );
  NAND2_X1 U542 ( .A1(n561), .A2(n479), .ZN(n491) );
  NOR2_X1 U543 ( .A1(n480), .A2(n491), .ZN(n487) );
  NAND2_X1 U544 ( .A1(n487), .A2(n514), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U546 ( .A(G57GAT), .B(n483), .Z(G1332GAT) );
  XOR2_X1 U547 ( .A(G64GAT), .B(KEYINPUT107), .Z(n485) );
  NAND2_X1 U548 ( .A1(n487), .A2(n544), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n485), .B(n484), .ZN(G1333GAT) );
  NAND2_X1 U550 ( .A1(n519), .A2(n487), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n486), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n489) );
  NAND2_X1 U553 ( .A1(n487), .A2(n496), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U555 ( .A(G78GAT), .B(n490), .ZN(G1335GAT) );
  NOR2_X1 U556 ( .A1(n492), .A2(n491), .ZN(n497) );
  NAND2_X1 U557 ( .A1(n514), .A2(n497), .ZN(n493) );
  XNOR2_X1 U558 ( .A(G85GAT), .B(n493), .ZN(G1336GAT) );
  NAND2_X1 U559 ( .A1(n497), .A2(n544), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n494), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U561 ( .A1(n519), .A2(n497), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n495), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n499) );
  NAND2_X1 U564 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n500), .ZN(G1339GAT) );
  NOR2_X1 U567 ( .A1(n586), .A2(n526), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(KEYINPUT45), .ZN(n504) );
  INV_X1 U569 ( .A(n577), .ZN(n502) );
  NOR2_X1 U570 ( .A1(n573), .A2(n502), .ZN(n503) );
  AND2_X1 U571 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(KEYINPUT111), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n573), .A2(n561), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(KEYINPUT46), .ZN(n507) );
  NAND2_X1 U575 ( .A1(n507), .A2(n526), .ZN(n508) );
  NOR2_X1 U576 ( .A1(n541), .A2(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(KEYINPUT48), .ZN(n545) );
  NAND2_X1 U581 ( .A1(n514), .A2(n545), .ZN(n515) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(KEYINPUT112), .B(n517), .Z(n533) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U585 ( .A1(n533), .A2(n520), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n529), .A2(n573), .ZN(n523) );
  XOR2_X1 U587 ( .A(G113GAT), .B(KEYINPUT113), .Z(n521) );
  XNOR2_X1 U588 ( .A(KEYINPUT114), .B(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U591 ( .A1(n529), .A2(n561), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  INV_X1 U593 ( .A(n526), .ZN(n580) );
  NAND2_X1 U594 ( .A1(n529), .A2(n580), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U598 ( .A1(n529), .A2(n464), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U600 ( .A(G134GAT), .B(n532), .Z(G1343GAT) );
  NOR2_X1 U601 ( .A1(n533), .A2(n568), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(KEYINPUT116), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n540), .A2(n573), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n535), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n537) );
  NAND2_X1 U606 ( .A1(n561), .A2(n540), .ZN(n536) );
  XNOR2_X1 U607 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n538), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n540), .A2(n580), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n539), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U611 ( .A(G162GAT), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U612 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n543), .B(n542), .ZN(G1347GAT) );
  XOR2_X1 U614 ( .A(G169GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U615 ( .A1(n545), .A2(n544), .ZN(n548) );
  INV_X1 U616 ( .A(KEYINPUT118), .ZN(n546) );
  AND2_X1 U617 ( .A1(n569), .A2(n549), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n570), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U621 ( .A(KEYINPUT55), .B(n553), .Z(n554) );
  NAND2_X1 U622 ( .A1(n565), .A2(n573), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(n560), .Z(n563) );
  NAND2_X1 U628 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n580), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n464), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  INV_X1 U636 ( .A(n568), .ZN(n572) );
  AND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n585) );
  INV_X1 U639 ( .A(n585), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  OR2_X1 U644 ( .A1(n585), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G218GAT), .B(n589), .Z(G1355GAT) );
endmodule

