//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  XNOR2_X1  g000(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n191), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT94), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G237), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G214), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT94), .A3(G131), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n205), .A3(new_n202), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n196), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT71), .A2(G140), .ZN(new_n208));
  OAI21_X1  g022(.A(G125), .B1(KEYINPUT71), .B2(G140), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G125), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  OAI221_X1 g025(.A(KEYINPUT16), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT16), .A2(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(G146), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT19), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G125), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n211), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n209), .A2(new_n208), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(new_n225), .B2(KEYINPUT19), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n207), .B(new_n215), .C1(new_n216), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT18), .A2(G131), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT92), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n203), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n201), .A2(KEYINPUT92), .A3(new_n202), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G146), .B1(new_n223), .B2(new_n224), .ZN(new_n233));
  INV_X1    g047(.A(new_n216), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n217), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n228), .B(KEYINPUT93), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n201), .A3(new_n202), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n190), .B1(new_n227), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n232), .A2(new_n236), .A3(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT17), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n196), .B2(new_n204), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n196), .A2(new_n204), .A3(new_n206), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n242), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT16), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n223), .A2(new_n224), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n214), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n215), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n248), .A2(new_n249), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT73), .A3(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n241), .B1(new_n245), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n240), .B1(new_n256), .B2(new_n190), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT95), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n187), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n261));
  INV_X1    g075(.A(new_n259), .ZN(new_n262));
  INV_X1    g076(.A(new_n190), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n263), .B(new_n241), .C1(new_n245), .C2(new_n255), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n261), .B(new_n262), .C1(new_n264), .C2(new_n240), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G478), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT15), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G143), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n272), .A2(G143), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n200), .A2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n200), .A2(G128), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n273), .C1(new_n274), .C2(new_n271), .ZN(new_n280));
  XNOR2_X1  g094(.A(G116), .B(G122), .ZN(new_n281));
  INV_X1    g095(.A(G107), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n278), .B(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT9), .B(G234), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G217), .A3(new_n198), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G122), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT14), .B1(new_n291), .B2(G116), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT14), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(G122), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(G116), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G107), .ZN(new_n299));
  OAI21_X1  g113(.A(G134), .B1(new_n276), .B2(new_n277), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n279), .A2(new_n273), .A3(new_n271), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n302), .A3(new_n283), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n298), .B1(new_n297), .B2(G107), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n286), .B(new_n290), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n297), .A2(G107), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT96), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n300), .A2(new_n301), .B1(new_n282), .B2(new_n281), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n299), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n290), .B1(new_n310), .B2(new_n286), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n270), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT97), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n286), .B1(new_n303), .B2(new_n304), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n289), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n305), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT97), .A3(new_n270), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n269), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G952), .ZN(new_n320));
  AOI211_X1 g134(.A(G953), .B(new_n320), .C1(G234), .C2(G237), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT21), .B(G898), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n270), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n312), .A2(new_n268), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n319), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n256), .A2(new_n190), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n270), .B1(new_n328), .B2(new_n264), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G475), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n266), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT98), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n260), .A2(new_n265), .B1(new_n329), .B2(G475), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT98), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(new_n327), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(G221), .B1(new_n287), .B2(G902), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G469), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n198), .A2(G227), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT80), .ZN(new_n342));
  XNOR2_X1  g156(.A(G110), .B(G140), .ZN(new_n343));
  XOR2_X1   g157(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n282), .A2(G104), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n189), .B2(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n282), .A2(KEYINPUT3), .A3(G104), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G101), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n348), .A2(new_n349), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT82), .B(G101), .ZN(new_n356));
  INV_X1    g170(.A(new_n346), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT83), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n350), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(new_n352), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n246), .A2(KEYINPUT64), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G146), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n366), .A3(new_n200), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n246), .A2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT0), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(new_n272), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT0), .A2(G128), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n246), .B2(G143), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n200), .A2(KEYINPUT65), .A3(G146), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n365), .A2(G146), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n246), .A2(KEYINPUT64), .ZN(new_n380));
  OAI21_X1  g194(.A(G143), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(new_n381), .A3(new_n371), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n363), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n359), .A2(new_n361), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n378), .A2(new_n381), .A3(new_n387), .A4(G128), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n200), .B1(new_n364), .B2(new_n366), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n376), .A2(new_n377), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(G143), .B2(new_n246), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n389), .A2(new_n390), .B1(new_n272), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g207(.A(G104), .B(G107), .Z(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n397));
  OAI21_X1  g211(.A(G128), .B1(new_n389), .B2(new_n387), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n369), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n359), .A2(new_n361), .B1(G101), .B2(new_n394), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n396), .A2(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT11), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n271), .B2(G137), .ZN(new_n404));
  INV_X1    g218(.A(G137), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT11), .A3(G134), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n271), .A2(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G131), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n406), .A3(new_n205), .A4(new_n407), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n385), .A2(new_n402), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n412), .B1(new_n385), .B2(new_n402), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n340), .B(new_n345), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n385), .A2(new_n402), .A3(new_n412), .ZN(new_n416));
  AND4_X1   g230(.A1(new_n360), .A2(new_n355), .A3(new_n356), .A4(new_n357), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n360), .B1(new_n350), .B2(new_n356), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n395), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n399), .A3(new_n388), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n396), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT12), .B1(new_n421), .B2(new_n411), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n423), .B(new_n412), .C1(new_n420), .C2(new_n396), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n416), .B(new_n344), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n396), .A2(new_n397), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n400), .A2(new_n401), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT4), .B1(new_n417), .B2(new_n418), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n350), .A2(new_n351), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n383), .B1(new_n432), .B2(new_n353), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n411), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n416), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n340), .B1(new_n435), .B2(new_n345), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n339), .B(new_n270), .C1(new_n426), .C2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n413), .A2(new_n345), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n416), .B1(new_n422), .B2(new_n424), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n344), .B(KEYINPUT81), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n438), .A2(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G469), .B1(new_n441), .B2(G902), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n338), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n336), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT76), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT22), .B(G137), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n215), .A2(new_n235), .ZN(new_n449));
  XOR2_X1   g263(.A(KEYINPUT74), .B(G110), .Z(new_n450));
  AND2_X1   g264(.A1(KEYINPUT67), .A2(G119), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT67), .A2(G119), .ZN(new_n452));
  OAI21_X1  g266(.A(G128), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G119), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G128), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(KEYINPUT23), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n451), .A2(new_n452), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n272), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n450), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n453), .A2(new_n456), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT24), .B(G110), .Z(new_n464));
  OAI22_X1  g278(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n449), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n457), .A2(new_n460), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n468), .A2(G110), .B1(new_n463), .B2(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n252), .A2(new_n254), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT77), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n471), .B1(new_n467), .B2(new_n470), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n448), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n470), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT77), .ZN(new_n476));
  INV_X1    g290(.A(new_n448), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G234), .ZN(new_n480));
  AOI21_X1  g294(.A(G902), .B1(new_n480), .B2(G217), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT79), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n270), .A3(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G217), .B1(new_n480), .B2(G902), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT70), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n484), .A2(new_n486), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n474), .A2(KEYINPUT25), .A3(new_n478), .A4(new_n270), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(KEYINPUT78), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n483), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n411), .A2(new_n382), .A3(new_n374), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n407), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n271), .A2(G137), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(new_n410), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT1), .B1(new_n216), .B2(new_n200), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n502), .A2(G128), .B1(new_n368), .B2(new_n367), .ZN(new_n503));
  NOR4_X1   g317(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT1), .A4(new_n272), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n411), .A2(new_n382), .A3(new_n374), .A4(KEYINPUT66), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G116), .B1(new_n451), .B2(new_n452), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n294), .A2(G119), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g326(.A(KEYINPUT2), .B(G113), .Z(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n510), .A3(new_n511), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n411), .A2(new_n382), .A3(new_n374), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n519), .A2(new_n505), .A3(KEYINPUT30), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n509), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(new_n505), .A3(new_n517), .A4(new_n521), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n191), .A2(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT31), .ZN(new_n531));
  INV_X1    g345(.A(new_n529), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n507), .A2(new_n518), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n524), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n517), .A2(new_n495), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT28), .B1(new_n536), .B2(new_n505), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n532), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT31), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n523), .A2(new_n539), .A3(new_n524), .A4(new_n529), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G472), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n270), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n541), .A2(KEYINPUT32), .A3(new_n542), .A4(new_n270), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n519), .A2(new_n505), .A3(new_n521), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n518), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n533), .B1(new_n548), .B2(new_n524), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n537), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n550), .A2(KEYINPUT29), .A3(new_n529), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n270), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n535), .A2(new_n537), .A3(new_n532), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n529), .B1(new_n523), .B2(new_n524), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT29), .ZN(new_n555));
  OAI21_X1  g369(.A(G472), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n545), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n383), .A2(new_n210), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT88), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n383), .A2(KEYINPUT88), .A3(new_n210), .ZN(new_n563));
  INV_X1    g377(.A(new_n210), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n399), .A2(new_n564), .A3(new_n388), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G224), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n562), .A2(new_n570), .A3(new_n563), .A4(new_n565), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT5), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(G116), .C1(new_n451), .C2(new_n452), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G113), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n510), .A2(KEYINPUT5), .A3(new_n511), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n516), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n401), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(G110), .B(G122), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT86), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n431), .A2(new_n354), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n430), .B2(new_n431), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n580), .B(new_n583), .C1(new_n585), .C2(new_n517), .ZN(new_n586));
  INV_X1    g400(.A(new_n578), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n515), .B1(new_n587), .B2(new_n576), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n419), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n363), .B2(new_n518), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n581), .B(KEYINPUT86), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT87), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n586), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT6), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n580), .B1(new_n585), .B2(new_n517), .ZN(new_n595));
  INV_X1    g409(.A(new_n592), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT6), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n573), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n576), .A2(KEYINPUT89), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT89), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n575), .B2(G113), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n600), .A2(new_n587), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n401), .B1(new_n603), .B2(new_n516), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n583), .A2(KEYINPUT8), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT8), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n591), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n579), .A2(new_n419), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n568), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n562), .A2(new_n563), .A3(new_n565), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n565), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n610), .B2(new_n568), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n609), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n586), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n270), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n559), .B1(new_n599), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(G902), .B1(new_n615), .B2(new_n586), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n597), .B1(KEYINPUT6), .B2(new_n593), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n619), .B(new_n558), .C1(new_n620), .C2(new_n573), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(KEYINPUT90), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(G214), .B1(G237), .B2(G902), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT85), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n599), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n558), .A4(new_n619), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n622), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n444), .A2(new_n494), .A3(new_n557), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(new_n356), .Z(G3));
  INV_X1    g446(.A(new_n483), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n491), .A2(KEYINPUT78), .A3(new_n492), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n487), .A2(new_n489), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n437), .A2(new_n442), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n337), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n541), .A2(new_n270), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(G472), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n543), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n621), .A2(KEYINPUT99), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n618), .ZN(new_n644));
  OAI211_X1 g458(.A(KEYINPUT99), .B(new_n559), .C1(new_n599), .C2(new_n617), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n624), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n266), .A2(new_n330), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n317), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n316), .A2(KEYINPUT33), .A3(new_n305), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n267), .A2(G902), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n314), .A2(new_n318), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n267), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n325), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n642), .A2(new_n646), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT34), .B(G104), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  OR3_X1    g476(.A1(new_n257), .A2(new_n187), .A3(new_n259), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n260), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n330), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n319), .A2(new_n326), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n325), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n642), .A2(new_n646), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT35), .B(G107), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  INV_X1    g484(.A(new_n482), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n475), .B(new_n672), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n490), .A2(new_n493), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n641), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(new_n444), .A3(new_n630), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n634), .B2(new_n635), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n557), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n644), .A2(new_n645), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n625), .A3(new_n443), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n324), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n321), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n665), .A2(new_n666), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n272), .ZN(G30));
  INV_X1    g507(.A(new_n666), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n647), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n688), .B(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n443), .A2(new_n698), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n624), .B(new_n695), .C1(new_n699), .C2(KEYINPUT40), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n532), .B1(new_n523), .B2(new_n524), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n548), .A2(new_n524), .A3(new_n532), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n270), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n545), .A2(new_n546), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n674), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n622), .A2(new_n628), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT38), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n700), .A2(new_n706), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n647), .A2(new_n657), .A3(new_n688), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n684), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT102), .B(G146), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G48));
  NAND3_X1  g530(.A1(new_n557), .A2(new_n494), .A3(new_n659), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n270), .B1(new_n426), .B2(new_n436), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n719), .A2(new_n337), .A3(new_n437), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n646), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n557), .A2(new_n494), .A3(new_n667), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n721), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n294), .ZN(G18));
  NAND3_X1  g541(.A1(new_n557), .A2(new_n680), .A3(new_n336), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n454), .ZN(G21));
  NAND2_X1  g544(.A1(new_n636), .A2(KEYINPUT104), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n532), .B1(new_n549), .B2(new_n537), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n531), .A2(new_n540), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NOR2_X1   g550(.A1(G472), .A2(G902), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n542), .B1(new_n541), .B2(new_n270), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n731), .A2(new_n733), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n325), .ZN(new_n744));
  INV_X1    g558(.A(new_n695), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n646), .A2(new_n720), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n291), .ZN(G24));
  AND2_X1   g562(.A1(new_n646), .A2(new_n720), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n740), .A2(new_n741), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n680), .A2(new_n738), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n647), .A2(new_n753), .A3(new_n657), .A4(new_n688), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n749), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G125), .ZN(G27));
  AND3_X1   g571(.A1(new_n545), .A2(KEYINPUT108), .A3(new_n546), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT108), .B1(new_n545), .B2(new_n546), .ZN(new_n759));
  INV_X1    g573(.A(new_n556), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n731), .A2(new_n733), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n707), .A2(new_n625), .A3(new_n443), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(KEYINPUT42), .A3(new_n755), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n557), .A2(new_n494), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n755), .A3(new_n765), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT42), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n768), .A2(KEYINPUT106), .A3(new_n765), .A4(new_n755), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n624), .B1(new_n622), .B2(new_n628), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n557), .A2(new_n775), .A3(new_n494), .A4(new_n443), .ZN(new_n776));
  INV_X1    g590(.A(new_n755), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT42), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n767), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n205), .ZN(G33));
  NAND3_X1  g597(.A1(new_n768), .A2(new_n690), .A3(new_n765), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  INV_X1    g599(.A(new_n775), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n647), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n641), .A3(new_n680), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n786), .B1(new_n793), .B2(KEYINPUT44), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n441), .A2(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n441), .A2(KEYINPUT45), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(G469), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(G469), .A2(G902), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n437), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n797), .B2(new_n798), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n337), .B(new_n698), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n794), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT109), .B(G137), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G39));
  OAI21_X1  g622(.A(new_n337), .B1(new_n800), .B2(new_n801), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(KEYINPUT47), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n786), .A2(new_n557), .A3(new_n494), .A4(new_n713), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G140), .ZN(G42));
  INV_X1    g628(.A(new_n762), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n647), .A2(new_n787), .A3(new_n624), .A4(new_n338), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n719), .A2(new_n437), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT110), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT110), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n705), .B(new_n709), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  INV_X1    g638(.A(new_n713), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n681), .B(new_n683), .C1(new_n690), .C2(new_n825), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n624), .B(new_n695), .C1(new_n644), .C2(new_n645), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n638), .A2(new_n689), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n706), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(new_n756), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n721), .B1(new_n717), .B2(new_n725), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n747), .A2(new_n832), .A3(new_n729), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n755), .A2(new_n742), .A3(new_n680), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n775), .A2(new_n443), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT112), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n751), .A2(new_n765), .A3(new_n837), .A4(new_n755), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT111), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n647), .B2(new_n666), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n658), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n787), .A2(new_n333), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n840), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n325), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n638), .A2(new_n641), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n494), .A4(new_n630), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n631), .A3(new_n676), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n665), .A2(new_n694), .A3(new_n689), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n557), .A2(new_n680), .A3(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n776), .A2(new_n691), .B1(new_n850), .B2(new_n835), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n831), .A2(new_n833), .A3(new_n839), .A4(new_n852), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n764), .A2(new_n766), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n826), .A2(new_n756), .A3(new_n858), .A4(new_n829), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(new_n857), .A3(KEYINPUT53), .A4(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT114), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n836), .A2(new_n838), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n336), .A2(new_n443), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n629), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n768), .B2(new_n675), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n765), .A2(new_n557), .A3(new_n680), .A4(new_n849), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n784), .A3(new_n867), .A4(new_n847), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n859), .A3(new_n831), .A4(new_n833), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n862), .B1(new_n870), .B2(new_n782), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n824), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  INV_X1    g691(.A(new_n720), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n709), .A2(new_n625), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n743), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n687), .B1(new_n789), .B2(new_n790), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n876), .B(new_n877), .C1(new_n880), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n877), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n879), .A2(new_n881), .A3(new_n885), .A4(new_n882), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n886), .C1(new_n876), .C2(new_n877), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n882), .A2(new_n720), .A3(new_n775), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n494), .A2(new_n321), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n878), .A2(new_n889), .A3(new_n786), .A4(new_n705), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n647), .A2(new_n657), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n751), .A2(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n881), .A2(new_n775), .A3(new_n882), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n810), .A2(new_n811), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n337), .B1(new_n818), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n896), .B2(new_n818), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n875), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n883), .A2(new_n721), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT119), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n320), .B(G953), .C1(new_n890), .C2(new_n843), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT48), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n888), .B2(new_n763), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n888), .A2(new_n763), .A3(new_n906), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n904), .B(new_n905), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT118), .B1(new_n895), .B2(new_n898), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n894), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n895), .A2(KEYINPUT118), .A3(new_n898), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n875), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n893), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT117), .B(new_n875), .C1(new_n893), .C2(new_n899), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n902), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n860), .A2(new_n871), .A3(new_n824), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n874), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n823), .B1(new_n919), .B2(new_n920), .ZN(G75));
  OR3_X1    g735(.A1(new_n198), .A2(KEYINPUT120), .A3(G952), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT120), .B1(new_n198), .B2(G952), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT121), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT56), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n860), .A2(new_n871), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(G902), .ZN(new_n929));
  INV_X1    g743(.A(G210), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n620), .B(new_n572), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n933), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(G51));
  AOI211_X1 g750(.A(new_n270), .B(new_n797), .C1(new_n860), .C2(new_n871), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n798), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n824), .B1(new_n860), .B2(new_n871), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n918), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n426), .A2(new_n436), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n937), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT122), .B1(new_n943), .B2(new_n924), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(new_n924), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n852), .A2(new_n833), .A3(new_n839), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n830), .A2(KEYINPUT52), .ZN(new_n948));
  INV_X1    g762(.A(new_n859), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT53), .B1(new_n950), .B2(new_n857), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n870), .A2(new_n782), .A3(new_n862), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT54), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n860), .A2(new_n871), .A3(new_n824), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n941), .B1(new_n955), .B2(new_n938), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n945), .B(new_n946), .C1(new_n956), .C2(new_n937), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n944), .A2(new_n957), .ZN(G54));
  INV_X1    g772(.A(new_n257), .ZN(new_n959));
  NAND2_X1  g773(.A1(KEYINPUT58), .A2(G475), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n929), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n929), .B2(new_n960), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n924), .B1(new_n961), .B2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(new_n649), .A2(new_n650), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n918), .B2(new_n939), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT123), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(new_n967), .C1(new_n918), .C2(new_n939), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n925), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n966), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n874), .B2(new_n918), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n964), .B2(new_n974), .ZN(G63));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT60), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n928), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n926), .B1(new_n979), .B2(new_n673), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n479), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(KEYINPUT61), .A3(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  OAI21_X1  g800(.A(G953), .B1(new_n323), .B2(new_n567), .ZN(new_n987));
  NOR4_X1   g801(.A1(new_n848), .A2(new_n747), .A3(new_n832), .A4(new_n729), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n990), .B2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n620), .B1(G898), .B2(new_n198), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n509), .A2(new_n522), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n226), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n842), .A2(new_n844), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT125), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n786), .A2(new_n699), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n768), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n806), .A2(new_n813), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n711), .A2(new_n756), .A3(new_n826), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT62), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(new_n1005), .A3(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT126), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n994), .B(new_n997), .C1(new_n1009), .C2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(G953), .B1(new_n1013), .B2(new_n1006), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT127), .B1(new_n1014), .B2(new_n996), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n997), .B1(G900), .B2(G953), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n794), .A2(new_n805), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n763), .A2(new_n827), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n802), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n813), .A2(new_n756), .A3(new_n784), .A4(new_n826), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n782), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1016), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1010), .A2(new_n1015), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1024), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1010), .A2(new_n1015), .A3(new_n1026), .A4(new_n1022), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  INV_X1    g844(.A(new_n530), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n554), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n861), .B2(new_n873), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1030), .B1(new_n1021), .B2(new_n989), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n523), .A2(new_n524), .A3(new_n532), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n946), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1009), .A2(new_n990), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n1030), .ZN(new_n1039));
  AOI211_X1 g853(.A(new_n1033), .B(new_n1037), .C1(new_n701), .C2(new_n1039), .ZN(G57));
endmodule


