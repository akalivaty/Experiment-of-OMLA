//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT31), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT64), .B(new_n192), .C1(new_n193), .C2(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(G137), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n191), .B1(new_n198), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n197), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(G134), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT64), .B1(new_n206), .B2(new_n192), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n202), .B(new_n191), .C1(new_n205), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(new_n201), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n196), .B2(new_n197), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(new_n191), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n204), .B1(new_n209), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n220), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT0), .B(G128), .Z(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n212), .A2(new_n210), .A3(new_n191), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n203), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n216), .A2(new_n226), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT1), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n218), .A2(new_n220), .A3(new_n232), .A4(G128), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n224), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n191), .B1(new_n206), .B2(new_n201), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n209), .B2(new_n213), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G119), .ZN(new_n242));
  OR3_X1    g056(.A1(new_n241), .A2(new_n242), .A3(KEYINPUT66), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n231), .A2(new_n240), .A3(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(KEYINPUT68), .A2(G953), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT68), .A2(G953), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(G210), .A3(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT26), .B(G101), .Z(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g067(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT70), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n253), .B(new_n255), .Z(new_n256));
  AND2_X1   g070(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n231), .A2(KEYINPUT30), .A3(new_n240), .ZN(new_n258));
  INV_X1    g072(.A(new_n226), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n240), .B1(new_n229), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n245), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n189), .B(new_n190), .C1(new_n257), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n246), .A3(new_n256), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT71), .B1(new_n265), .B2(KEYINPUT31), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n256), .B(KEYINPUT73), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n246), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n245), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n260), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n269), .B1(new_n246), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n268), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n257), .A2(new_n263), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n187), .B(new_n188), .C1(new_n267), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n275), .B(new_n278), .C1(new_n264), .C2(new_n266), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n231), .A2(new_n240), .A3(new_n245), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n258), .B2(new_n262), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n287), .B2(new_n256), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n263), .A2(new_n246), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n290));
  INV_X1    g104(.A(new_n256), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n274), .ZN(new_n293));
  INV_X1    g107(.A(new_n268), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n270), .A3(new_n294), .ZN(new_n295));
  AND4_X1   g109(.A1(new_n285), .A2(new_n288), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n245), .B1(new_n231), .B2(new_n240), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT28), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n291), .A2(new_n285), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n270), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(KEYINPUT75), .A3(new_n270), .A4(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n188), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G472), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n282), .A2(new_n284), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n236), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g121(.A(G104), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT80), .B1(new_n308), .B2(G107), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(G107), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n308), .A2(KEYINPUT80), .A3(G107), .ZN(new_n312));
  OAI21_X1  g126(.A(G101), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(new_n308), .B2(G107), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  INV_X1    g129(.A(G107), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G104), .ZN(new_n317));
  INV_X1    g131(.A(G101), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n314), .A2(new_n317), .A3(new_n318), .A4(new_n310), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT82), .B1(new_n307), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT10), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n232), .B1(G143), .B2(new_n217), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n223), .B1(new_n323), .B2(new_n234), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n322), .B1(new_n324), .B2(new_n233), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n319), .A4(new_n313), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n233), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n218), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n323), .A2(KEYINPUT81), .ZN(new_n332));
  OAI21_X1  g146(.A(G128), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n333), .B2(new_n223), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n322), .B1(new_n334), .B2(new_n320), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n314), .A2(new_n317), .A3(new_n310), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(G101), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n319), .A2(KEYINPUT4), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n341), .A3(G101), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n226), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n328), .A2(new_n335), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n216), .A3(new_n230), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n321), .A2(new_n327), .B1(new_n340), .B2(new_n343), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n215), .B(new_n203), .C1(new_n227), .C2(new_n228), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n347), .B(new_n335), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n249), .A2(G227), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G140), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n346), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n348), .A2(new_n349), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n237), .A2(new_n320), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n334), .B2(new_n320), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT12), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n214), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n350), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G469), .B1(new_n362), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(G469), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT12), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n216), .A2(new_n230), .A3(new_n357), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n359), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n353), .B1(new_n355), .B2(new_n345), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n350), .A2(KEYINPUT83), .A3(new_n353), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n353), .B1(new_n346), .B2(new_n350), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n364), .B(new_n188), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT84), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n379), .B(new_n380), .C1(new_n363), .C2(new_n374), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G210), .B1(G237), .B2(G902), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n243), .A2(new_n342), .A3(new_n244), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n242), .A2(KEYINPUT5), .ZN(new_n386));
  INV_X1    g200(.A(G116), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n387), .A2(KEYINPUT5), .A3(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G113), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n241), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n242), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n385), .A2(new_n339), .B1(new_n320), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT85), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n236), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n259), .B2(new_n397), .ZN(new_n399));
  INV_X1    g213(.A(G953), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G224), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n401), .A2(KEYINPUT7), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n396), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n392), .B1(new_n320), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n320), .B2(KEYINPUT86), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n395), .B(KEYINPUT8), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n405), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n393), .A2(new_n395), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n396), .A2(KEYINPUT6), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n399), .B(new_n401), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n393), .A2(new_n416), .A3(new_n395), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n384), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n384), .A3(new_n418), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n383), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n378), .A2(new_n381), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  INV_X1    g240(.A(G140), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(G125), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n397), .A2(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(G146), .B(new_n428), .C1(new_n431), .C2(new_n426), .ZN(new_n432));
  XNOR2_X1  g246(.A(G125), .B(G140), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n217), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT23), .B1(new_n234), .B2(G119), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n436));
  INV_X1    g250(.A(G119), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(G128), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n435), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G110), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G119), .B(G128), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT24), .B(G110), .Z(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT79), .B1(new_n439), .B2(new_n440), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n432), .B(new_n434), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n432), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(KEYINPUT16), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n449), .A2(KEYINPUT78), .A3(G146), .A4(new_n428), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n428), .B1(new_n431), .B2(new_n426), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n217), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n443), .A2(new_n442), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n439), .B(KEYINPUT77), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n249), .A2(G221), .A3(G234), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT22), .B(G137), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n446), .B2(new_n456), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n425), .B1(new_n465), .B2(new_n188), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n425), .B(new_n188), .C1(new_n461), .C2(new_n463), .ZN(new_n468));
  INV_X1    g282(.A(G217), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(G234), .B2(new_n188), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n470), .A2(G902), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n467), .A2(new_n472), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n308), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT19), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n431), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n433), .A2(KEYINPUT89), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n217), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n248), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT68), .A2(G953), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(G214), .A3(new_n250), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n219), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n249), .A2(G143), .A3(G214), .A4(new_n250), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n191), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n191), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n485), .B(new_n432), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(KEYINPUT18), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT18), .A2(G131), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n481), .A2(new_n482), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n434), .B1(new_n497), .B2(new_n217), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n478), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n492), .A2(new_n491), .A3(KEYINPUT17), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n453), .B1(KEYINPUT17), .B2(new_n491), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n498), .A2(new_n496), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n502), .B1(new_n494), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(new_n478), .ZN(new_n505));
  INV_X1    g319(.A(G475), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n188), .ZN(new_n507));
  OAI211_X1 g321(.A(KEYINPUT90), .B(new_n476), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n493), .A2(new_n499), .ZN(new_n510));
  INV_X1    g324(.A(new_n478), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n491), .A2(KEYINPUT17), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(new_n450), .A3(new_n448), .A4(new_n452), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n492), .A2(new_n491), .A3(KEYINPUT17), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n478), .B(new_n499), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n507), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n509), .B1(new_n517), .B2(new_n475), .ZN(new_n518));
  INV_X1    g332(.A(new_n517), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n508), .B(new_n518), .C1(KEYINPUT20), .C2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n504), .A2(new_n478), .ZN(new_n521));
  INV_X1    g335(.A(new_n516), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n188), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G475), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n219), .A2(G128), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n234), .A2(G143), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G134), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(new_n527), .A3(new_n193), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G116), .B(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n316), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n387), .A2(G122), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(KEYINPUT14), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n387), .A2(G122), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n535), .B1(new_n537), .B2(KEYINPUT14), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n316), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT91), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n536), .A2(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G107), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n531), .A4(new_n533), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n532), .B(new_n316), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT13), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n526), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n527), .A2(KEYINPUT13), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n526), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n530), .C1(new_n193), .C2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n376), .A2(new_n469), .A3(G953), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n545), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n552), .B1(new_n545), .B2(new_n551), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n188), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  OAI221_X1 g372(.A(new_n188), .B1(KEYINPUT15), .B2(new_n556), .C1(new_n553), .C2(new_n554), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(G234), .A2(G237), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(G952), .A3(new_n400), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT92), .ZN(new_n563));
  INV_X1    g377(.A(new_n249), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(G902), .A3(new_n561), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT21), .B(G898), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n525), .A2(new_n560), .A3(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n306), .A2(new_n424), .A3(new_n474), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NOR2_X1   g385(.A1(new_n187), .A2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n283), .A2(new_n188), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n283), .B2(new_n188), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n378), .A2(new_n381), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n576), .A2(new_n474), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT33), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n581), .C1(new_n553), .C2(new_n554), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n545), .A2(new_n551), .ZN(new_n583));
  INV_X1    g397(.A(new_n552), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n545), .A2(new_n551), .A3(new_n552), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(KEYINPUT94), .A3(new_n579), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n556), .A2(G902), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n588), .A2(new_n589), .B1(new_n556), .B2(new_n555), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n520), .B2(new_n524), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n423), .A2(new_n592), .A3(new_n568), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n578), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XOR2_X1   g409(.A(KEYINPUT34), .B(G104), .Z(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  NAND2_X1  g411(.A1(new_n517), .A2(new_n475), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n508), .A2(new_n518), .A3(new_n598), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n523), .A2(G475), .B1(new_n558), .B2(new_n559), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n568), .B(KEYINPUT96), .Z(new_n601));
  AND4_X1   g415(.A1(new_n422), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n578), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT97), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT35), .B(G107), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n462), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT98), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(new_n457), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n473), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n466), .B2(new_n471), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n424), .A2(new_n576), .A3(new_n569), .A4(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT37), .B(G110), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT99), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n612), .B(new_n614), .ZN(G12));
  XOR2_X1   g429(.A(new_n563), .B(KEYINPUT100), .Z(new_n616));
  INV_X1    g430(.A(G900), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n566), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n599), .A2(new_n600), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT101), .A4(new_n619), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n622), .A2(new_n611), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n306), .A2(new_n424), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XOR2_X1   g440(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n618), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n577), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT40), .Z(new_n630));
  INV_X1    g444(.A(new_n297), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n294), .B1(new_n246), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n265), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n188), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n282), .A2(new_n284), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n421), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n419), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n525), .A2(new_n560), .ZN(new_n641));
  NOR4_X1   g455(.A1(new_n640), .A2(new_n383), .A3(new_n611), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n630), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT104), .B(G143), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G45));
  NAND2_X1  g459(.A1(new_n591), .A2(new_n619), .ZN(new_n646));
  INV_X1    g460(.A(new_n611), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n306), .A2(new_n424), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  OAI21_X1  g464(.A(new_n188), .B1(new_n372), .B2(new_n373), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(G469), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n377), .A3(new_n374), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT105), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n306), .A2(new_n654), .A3(new_n593), .A4(new_n474), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT41), .B(G113), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G15));
  NAND4_X1  g471(.A1(new_n306), .A2(new_n654), .A3(new_n474), .A4(new_n602), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G116), .ZN(G18));
  NAND4_X1  g473(.A1(new_n422), .A2(new_n377), .A3(new_n652), .A4(new_n374), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n569), .A2(new_n611), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n306), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G119), .ZN(G21));
  AOI21_X1  g478(.A(new_n187), .B1(new_n283), .B2(new_n188), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n265), .A2(KEYINPUT31), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n278), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n298), .A2(new_n270), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n268), .ZN(new_n669));
  AOI211_X1 g483(.A(G472), .B(G902), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n422), .A2(new_n601), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n641), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n654), .A2(new_n671), .A3(new_n474), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(G122), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G24));
  NOR3_X1   g490(.A1(new_n665), .A2(new_n670), .A3(new_n647), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n591), .A2(new_n678), .A3(new_n619), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n591), .B2(new_n619), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n660), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT108), .B(G125), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G27));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n375), .A2(new_n377), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n637), .A2(new_n419), .A3(new_n383), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n685), .A2(KEYINPUT42), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n266), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n265), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n279), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(KEYINPUT109), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n284), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n696), .B(new_n698), .C1(KEYINPUT110), .C2(new_n282), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n282), .A2(KEYINPUT110), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n305), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n690), .B(new_n474), .C1(new_n699), .C2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n306), .A2(new_n474), .A3(new_n685), .A4(new_n689), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n702), .A2(new_n705), .A3(KEYINPUT111), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n191), .ZN(G33));
  AND2_X1   g525(.A1(new_n622), .A2(new_n623), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n306), .A2(new_n474), .A3(new_n712), .A4(new_n689), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G134), .ZN(G36));
  INV_X1    g528(.A(new_n525), .ZN(new_n715));
  INV_X1    g529(.A(new_n590), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n717), .B(KEYINPUT43), .Z(new_n718));
  OAI211_X1 g532(.A(new_n718), .B(new_n611), .C1(new_n574), .C2(new_n575), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n687), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n720), .B2(new_n719), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n362), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n364), .A2(new_n188), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(KEYINPUT112), .A3(new_n374), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(G469), .C1(new_n724), .C2(G902), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n731), .A2(KEYINPUT113), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(KEYINPUT113), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT112), .B1(new_n728), .B2(new_n374), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n377), .B(new_n628), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n722), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT114), .B(G137), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G39));
  OAI21_X1  g554(.A(new_n377), .B1(new_n734), .B2(new_n735), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n306), .A2(new_n474), .A3(new_n646), .A4(new_n688), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT115), .Z(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G140), .ZN(G42));
  AND2_X1   g563(.A1(new_n652), .A2(new_n374), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT49), .Z(new_n751));
  NOR2_X1   g565(.A1(new_n380), .A2(new_n383), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n640), .A2(new_n474), .A3(new_n752), .ZN(new_n753));
  OR4_X1    g567(.A1(new_n636), .A2(new_n751), .A3(new_n717), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n718), .A2(new_n616), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n750), .A2(new_n377), .A3(new_n687), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n677), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n474), .A2(new_n563), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n636), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n715), .A2(new_n590), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n671), .A2(new_n474), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n755), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n750), .A2(new_n383), .A3(new_n377), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n640), .A3(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n765), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n766), .B1(new_n765), .B2(new_n771), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n762), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n764), .A2(new_n687), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT116), .Z(new_n776));
  NAND2_X1  g590(.A1(new_n750), .A2(new_n380), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n743), .A2(new_n744), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n778), .B2(KEYINPUT118), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(KEYINPUT118), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT51), .B(new_n774), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n699), .A2(new_n701), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n474), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n757), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n760), .A2(new_n592), .ZN(new_n788));
  OAI211_X1 g602(.A(G952), .B(new_n400), .C1(new_n765), .C2(new_n660), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n776), .A2(new_n778), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n774), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n781), .B(new_n790), .C1(KEYINPUT51), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n380), .B1(new_n363), .B2(new_n374), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n647), .A3(new_n619), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n796), .A2(new_n423), .A3(new_n641), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n636), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n625), .A2(new_n649), .A3(new_n682), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n686), .A2(new_n379), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(KEYINPUT84), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n422), .A2(new_n802), .A3(new_n624), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n804), .A2(new_n306), .B1(new_n677), .B2(new_n681), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n649), .A4(new_n798), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n655), .A2(new_n658), .A3(new_n674), .A4(new_n663), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n715), .A2(new_n560), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n672), .B1(new_n809), .B2(new_n592), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n576), .A2(new_n577), .A3(new_n474), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n570), .A2(new_n612), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n677), .A2(new_n685), .A3(new_n689), .ZN(new_n813));
  AOI211_X1 g627(.A(new_n618), .B(new_n560), .C1(G475), .C2(new_n523), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n599), .A2(new_n687), .A3(new_n611), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n306), .A2(new_n577), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n713), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n808), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n807), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n794), .B1(new_n819), .B2(new_n710), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n812), .A2(new_n817), .A3(new_n794), .ZN(new_n822));
  INV_X1    g636(.A(new_n808), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n807), .A2(new_n822), .A3(new_n706), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n807), .A2(new_n818), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n708), .A2(new_n709), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n819), .A2(new_n710), .A3(new_n794), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n825), .B1(new_n830), .B2(new_n821), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n793), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(G952), .A2(G953), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n754), .B1(new_n832), .B2(new_n833), .ZN(G75));
  XNOR2_X1  g648(.A(new_n415), .B(KEYINPUT55), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n414), .A2(new_n417), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT120), .Z(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n188), .B1(new_n820), .B2(new_n824), .ZN(new_n840));
  AOI211_X1 g654(.A(KEYINPUT56), .B(new_n839), .C1(new_n840), .C2(G210), .ZN(new_n841));
  INV_X1    g655(.A(new_n824), .ZN(new_n842));
  OAI211_X1 g656(.A(G210), .B(G902), .C1(new_n828), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n836), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(G210), .ZN(new_n847));
  AOI211_X1 g661(.A(new_n847), .B(new_n188), .C1(new_n820), .C2(new_n824), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n839), .B1(new_n848), .B2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n843), .A2(new_n844), .A3(new_n838), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n850), .A3(new_n835), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n249), .A2(G952), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n846), .A2(new_n851), .A3(new_n853), .ZN(G51));
  NAND2_X1  g668(.A1(new_n820), .A2(new_n824), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n825), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n726), .B(KEYINPUT57), .Z(new_n858));
  OAI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(new_n373), .B2(new_n372), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(G469), .A3(new_n724), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n852), .B1(new_n859), .B2(new_n860), .ZN(G54));
  AND2_X1   g675(.A1(KEYINPUT58), .A2(G475), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n840), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n505), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n853), .B1(new_n863), .B2(new_n505), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n863), .B2(new_n505), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G60));
  NAND2_X1  g682(.A1(G478), .A2(G902), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT59), .Z(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n588), .B1(new_n831), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n588), .A2(new_n871), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n873), .B(new_n853), .C1(new_n857), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n856), .B2(new_n825), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT122), .B1(new_n876), .B2(new_n852), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n872), .B1(new_n875), .B2(new_n877), .ZN(G63));
  XOR2_X1   g692(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n469), .A2(new_n188), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n880), .B(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n855), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n609), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n853), .B1(new_n883), .B2(new_n465), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n879), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n883), .A2(new_n465), .ZN(new_n888));
  INV_X1    g702(.A(new_n879), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n853), .A3(new_n884), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n887), .A2(new_n890), .ZN(G66));
  INV_X1    g705(.A(G224), .ZN(new_n892));
  OAI21_X1  g706(.A(G953), .B1(new_n567), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n808), .A2(new_n812), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n564), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n839), .B1(G898), .B2(new_n249), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(G69));
  AND2_X1   g711(.A1(new_n805), .A2(new_n649), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n643), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n745), .A2(new_n747), .B1(new_n722), .B2(new_n737), .ZN(new_n902));
  INV_X1    g716(.A(new_n629), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n688), .B1(new_n809), .B2(new_n592), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n306), .A3(new_n474), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n249), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n260), .A2(new_n261), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n258), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n483), .A2(new_n484), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n909), .B(new_n910), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(G227), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n564), .B1(new_n913), .B2(new_n617), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n249), .A2(G900), .ZN(new_n917));
  INV_X1    g731(.A(new_n641), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n783), .A2(new_n737), .A3(new_n422), .A4(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n898), .A2(new_n713), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n902), .A2(new_n827), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n917), .B1(new_n921), .B2(new_n249), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n912), .B(new_n916), .C1(new_n911), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n249), .ZN(new_n924));
  INV_X1    g738(.A(new_n917), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n911), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n911), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n906), .B2(new_n249), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n915), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n923), .A2(new_n929), .ZN(G72));
  NAND2_X1  g744(.A1(G472), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT63), .Z(new_n932));
  INV_X1    g746(.A(new_n894), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n921), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n289), .A2(new_n256), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n852), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n288), .A2(new_n265), .A3(new_n292), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n932), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n936), .B1(new_n830), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n901), .A2(new_n894), .A3(new_n902), .A4(new_n905), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n940), .A2(KEYINPUT126), .A3(new_n932), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT126), .B1(new_n940), .B2(new_n932), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n289), .A2(new_n256), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n939), .A2(new_n944), .ZN(G57));
endmodule


