

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U562 ( .A1(G651), .A2(n641), .ZN(n661) );
  AND2_X1 U563 ( .A1(n1013), .A2(n788), .ZN(n527) );
  AND2_X1 U564 ( .A1(n740), .A2(G1996), .ZN(n714) );
  NOR2_X1 U565 ( .A1(n719), .A2(n1021), .ZN(n722) );
  INV_X1 U566 ( .A(KEYINPUT98), .ZN(n720) );
  AND2_X1 U567 ( .A1(n716), .A2(n715), .ZN(n740) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U569 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n753) );
  XNOR2_X1 U570 ( .A(n754), .B(n753), .ZN(n768) );
  INV_X1 U571 ( .A(n792), .ZN(n789) );
  INV_X1 U572 ( .A(KEYINPUT101), .ZN(n778) );
  INV_X1 U573 ( .A(KEYINPUT33), .ZN(n790) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n711) );
  AND2_X1 U575 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U576 ( .A(n711), .B(KEYINPUT64), .ZN(n715) );
  INV_X1 U577 ( .A(KEYINPUT17), .ZN(n531) );
  NAND2_X1 U578 ( .A1(n894), .A2(G138), .ZN(n557) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n540), .Z(n655) );
  INV_X1 U580 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n528), .A2(G2104), .ZN(n529) );
  XNOR2_X1 U582 ( .A(n529), .B(KEYINPUT65), .ZN(n555) );
  NAND2_X1 U583 ( .A1(G101), .A2(n555), .ZN(n530) );
  XOR2_X1 U584 ( .A(n530), .B(KEYINPUT23), .Z(n534) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  XNOR2_X2 U586 ( .A(n532), .B(n531), .ZN(n894) );
  NAND2_X1 U587 ( .A1(n894), .A2(G137), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n539) );
  AND2_X1 U589 ( .A1(G2105), .A2(G2104), .ZN(n899) );
  NAND2_X1 U590 ( .A1(G113), .A2(n899), .ZN(n537) );
  INV_X1 U591 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n535), .ZN(n900) );
  NAND2_X1 U593 ( .A1(G125), .A2(n900), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X2 U595 ( .A1(n539), .A2(n538), .ZN(G160) );
  INV_X1 U596 ( .A(G651), .ZN(n545) );
  NOR2_X1 U597 ( .A1(G543), .A2(n545), .ZN(n540) );
  NAND2_X1 U598 ( .A1(G63), .A2(n655), .ZN(n542) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n641) );
  NAND2_X1 U600 ( .A1(G51), .A2(n661), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT6), .B(n543), .ZN(n550) );
  NOR2_X1 U603 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U604 ( .A1(n654), .A2(G89), .ZN(n544) );
  XNOR2_X1 U605 ( .A(n544), .B(KEYINPUT4), .ZN(n547) );
  NOR2_X1 U606 ( .A1(n641), .A2(n545), .ZN(n652) );
  NAND2_X1 U607 ( .A1(G76), .A2(n652), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U609 ( .A(n548), .B(KEYINPUT5), .Z(n549) );
  NOR2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT74), .B(n551), .Z(n552) );
  XNOR2_X1 U612 ( .A(KEYINPUT7), .B(n552), .ZN(G168) );
  NAND2_X1 U613 ( .A1(G114), .A2(n899), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G126), .A2(n900), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n561) );
  INV_X1 U616 ( .A(KEYINPUT89), .ZN(n559) );
  BUF_X1 U617 ( .A(n555), .Z(n895) );
  NAND2_X1 U618 ( .A1(G102), .A2(n895), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n559), .B(n558), .ZN(n560) );
  NOR2_X2 U621 ( .A1(n561), .A2(n560), .ZN(G164) );
  NAND2_X1 U622 ( .A1(G64), .A2(n655), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n562), .B(KEYINPUT68), .ZN(n565) );
  NAND2_X1 U624 ( .A1(G52), .A2(n661), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n563), .Z(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U627 ( .A1(G90), .A2(n654), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G77), .A2(n652), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U631 ( .A1(n570), .A2(n569), .ZN(G171) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G82), .ZN(G220) );
  XOR2_X1 U636 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n840) );
  NAND2_X1 U640 ( .A1(n840), .A2(G567), .ZN(n572) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  XOR2_X1 U642 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n574) );
  NAND2_X1 U643 ( .A1(G56), .A2(n655), .ZN(n573) );
  XNOR2_X1 U644 ( .A(n574), .B(n573), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n654), .A2(G81), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U648 ( .A1(G68), .A2(n652), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n579), .B(n578), .ZN(n580) );
  NOR2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n661), .A2(G43), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n1021) );
  INV_X1 U654 ( .A(G860), .ZN(n603) );
  OR2_X1 U655 ( .A1(n1021), .A2(n603), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G54), .A2(n661), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G92), .A2(n654), .ZN(n585) );
  NAND2_X1 U660 ( .A1(G79), .A2(n652), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n655), .A2(G66), .ZN(n586) );
  XOR2_X1 U663 ( .A(KEYINPUT72), .B(n586), .Z(n587) );
  NOR2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U666 ( .A(n591), .B(KEYINPUT15), .ZN(n592) );
  XOR2_X2 U667 ( .A(KEYINPUT73), .B(n592), .Z(n1018) );
  OR2_X1 U668 ( .A1(n1018), .A2(G868), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G65), .A2(n655), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G53), .A2(n661), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G91), .A2(n654), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G78), .A2(n652), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n1005) );
  INV_X1 U677 ( .A(n1005), .ZN(G299) );
  NAND2_X1 U678 ( .A1(G868), .A2(G286), .ZN(n602) );
  INV_X1 U679 ( .A(G868), .ZN(n674) );
  NAND2_X1 U680 ( .A1(G299), .A2(n674), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U683 ( .A1(n604), .A2(n1018), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U685 ( .A1(G868), .A2(n1021), .ZN(n608) );
  NAND2_X1 U686 ( .A1(G868), .A2(n1018), .ZN(n606) );
  NOR2_X1 U687 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U689 ( .A(KEYINPUT75), .B(n609), .Z(G282) );
  NAND2_X1 U690 ( .A1(n895), .A2(G99), .ZN(n610) );
  XNOR2_X1 U691 ( .A(KEYINPUT77), .B(n610), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n899), .A2(G111), .ZN(n611) );
  XOR2_X1 U693 ( .A(KEYINPUT76), .B(n611), .Z(n612) );
  NOR2_X1 U694 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U695 ( .A(n614), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G135), .A2(n894), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n900), .A2(G123), .ZN(n617) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n978) );
  XOR2_X1 U701 ( .A(G2096), .B(n978), .Z(n620) );
  NOR2_X1 U702 ( .A1(G2100), .A2(n620), .ZN(n621) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n621), .ZN(G156) );
  NAND2_X1 U704 ( .A1(G559), .A2(n1018), .ZN(n622) );
  XNOR2_X1 U705 ( .A(n622), .B(n1021), .ZN(n669) );
  NOR2_X1 U706 ( .A1(n669), .A2(G860), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G93), .A2(n654), .ZN(n624) );
  NAND2_X1 U708 ( .A1(G67), .A2(n655), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G80), .A2(n652), .ZN(n626) );
  NAND2_X1 U711 ( .A1(G55), .A2(n661), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n627) );
  OR2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n673) );
  XOR2_X1 U714 ( .A(n629), .B(n673), .Z(G145) );
  NAND2_X1 U715 ( .A1(G88), .A2(n654), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G75), .A2(n652), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n661), .A2(G50), .ZN(n632) );
  XOR2_X1 U719 ( .A(KEYINPUT82), .B(n632), .Z(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n655), .A2(G62), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(G303) );
  INV_X1 U723 ( .A(G303), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G49), .A2(n661), .ZN(n638) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U727 ( .A(KEYINPUT80), .B(n639), .ZN(n640) );
  NOR2_X1 U728 ( .A1(n655), .A2(n640), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n641), .A2(G87), .ZN(n642) );
  NAND2_X1 U730 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U731 ( .A1(n652), .A2(G72), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G60), .A2(n655), .ZN(n645) );
  NAND2_X1 U733 ( .A1(G47), .A2(n661), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U735 ( .A1(G85), .A2(n654), .ZN(n646) );
  XOR2_X1 U736 ( .A(KEYINPUT66), .B(n646), .Z(n647) );
  NOR2_X1 U737 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U738 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U739 ( .A(KEYINPUT67), .B(n651), .Z(G290) );
  NAND2_X1 U740 ( .A1(G73), .A2(n652), .ZN(n653) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(n653), .Z(n660) );
  NAND2_X1 U742 ( .A1(G86), .A2(n654), .ZN(n657) );
  NAND2_X1 U743 ( .A1(G61), .A2(n655), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U745 ( .A(KEYINPUT81), .B(n658), .Z(n659) );
  NOR2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n661), .A2(G48), .ZN(n662) );
  NAND2_X1 U748 ( .A1(n663), .A2(n662), .ZN(G305) );
  XNOR2_X1 U749 ( .A(n673), .B(G166), .ZN(n664) );
  XNOR2_X1 U750 ( .A(n664), .B(G288), .ZN(n665) );
  XNOR2_X1 U751 ( .A(KEYINPUT19), .B(n665), .ZN(n667) );
  XNOR2_X1 U752 ( .A(G290), .B(n1005), .ZN(n666) );
  XNOR2_X1 U753 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U754 ( .A(n668), .B(G305), .ZN(n911) );
  XNOR2_X1 U755 ( .A(n911), .B(KEYINPUT83), .ZN(n670) );
  XNOR2_X1 U756 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G868), .A2(n671), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n672), .B(KEYINPUT84), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XOR2_X1 U766 ( .A(KEYINPUT85), .B(G44), .Z(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT3), .B(n681), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n682) );
  XOR2_X1 U769 ( .A(KEYINPUT22), .B(n682), .Z(n683) );
  NOR2_X1 U770 ( .A1(G218), .A2(n683), .ZN(n684) );
  XNOR2_X1 U771 ( .A(KEYINPUT86), .B(n684), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n685), .A2(G96), .ZN(n686) );
  XOR2_X1 U773 ( .A(KEYINPUT87), .B(n686), .Z(n844) );
  NAND2_X1 U774 ( .A1(n844), .A2(G2106), .ZN(n691) );
  NAND2_X1 U775 ( .A1(G120), .A2(G69), .ZN(n687) );
  NOR2_X1 U776 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n688), .A2(G108), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n689), .B(KEYINPUT88), .ZN(n845) );
  NAND2_X1 U779 ( .A1(G567), .A2(n845), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n846) );
  NAND2_X1 U781 ( .A1(G483), .A2(G661), .ZN(n692) );
  NOR2_X1 U782 ( .A1(n846), .A2(n692), .ZN(n843) );
  NAND2_X1 U783 ( .A1(n843), .A2(G36), .ZN(G176) );
  NAND2_X1 U784 ( .A1(G95), .A2(n895), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G107), .A2(n899), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G131), .A2(n894), .ZN(n695) );
  XNOR2_X1 U788 ( .A(KEYINPUT93), .B(n695), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n900), .A2(G119), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n906) );
  NAND2_X1 U792 ( .A1(n906), .A2(G1991), .ZN(n709) );
  NAND2_X1 U793 ( .A1(G117), .A2(n899), .ZN(n701) );
  NAND2_X1 U794 ( .A1(G129), .A2(n900), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n895), .A2(G105), .ZN(n702) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(n702), .Z(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U799 ( .A(n705), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U800 ( .A1(G141), .A2(n894), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n884) );
  NAND2_X1 U802 ( .A1(n884), .A2(G1996), .ZN(n708) );
  AND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n980) );
  NAND2_X1 U804 ( .A1(G40), .A2(G160), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n710), .B(KEYINPUT90), .ZN(n713) );
  NOR2_X1 U806 ( .A1(n713), .A2(n715), .ZN(n825) );
  INV_X1 U807 ( .A(n825), .ZN(n712) );
  NOR2_X1 U808 ( .A1(n980), .A2(n712), .ZN(n818) );
  XNOR2_X1 U809 ( .A(KEYINPUT95), .B(n713), .ZN(n716) );
  XOR2_X1 U810 ( .A(KEYINPUT26), .B(n714), .Z(n718) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n755) );
  NAND2_X1 U812 ( .A1(n755), .A2(G1341), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n722), .A2(n1018), .ZN(n721) );
  XNOR2_X1 U815 ( .A(n721), .B(n720), .ZN(n728) );
  NAND2_X1 U816 ( .A1(n722), .A2(n1018), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n740), .A2(G1348), .ZN(n724) );
  NOR2_X1 U818 ( .A1(G2067), .A2(n755), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n733) );
  NAND2_X1 U822 ( .A1(n740), .A2(G2072), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT27), .ZN(n731) );
  INV_X1 U824 ( .A(G1956), .ZN(n945) );
  NOR2_X1 U825 ( .A1(n945), .A2(n740), .ZN(n730) );
  NOR2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n1005), .A2(n734), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n1005), .A2(n734), .ZN(n735) );
  XOR2_X1 U830 ( .A(n735), .B(KEYINPUT28), .Z(n736) );
  NAND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U832 ( .A(n739), .B(n738), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n740), .A2(G1961), .ZN(n741) );
  XOR2_X1 U834 ( .A(KEYINPUT96), .B(n741), .Z(n744) );
  XOR2_X1 U835 ( .A(KEYINPUT25), .B(G2078), .Z(n927) );
  NOR2_X1 U836 ( .A1(n927), .A2(n755), .ZN(n742) );
  XNOR2_X1 U837 ( .A(KEYINPUT97), .B(n742), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n750), .A2(G171), .ZN(n745) );
  NAND2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n767) );
  NAND2_X1 U841 ( .A1(G8), .A2(n755), .ZN(n792) );
  NOR2_X1 U842 ( .A1(G1966), .A2(n792), .ZN(n771) );
  NOR2_X1 U843 ( .A1(G2084), .A2(n755), .ZN(n769) );
  NOR2_X1 U844 ( .A1(n771), .A2(n769), .ZN(n747) );
  NAND2_X1 U845 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U846 ( .A(n748), .B(KEYINPUT30), .ZN(n749) );
  NOR2_X1 U847 ( .A1(n749), .A2(G168), .ZN(n752) );
  NOR2_X1 U848 ( .A1(G171), .A2(n750), .ZN(n751) );
  NOR2_X1 U849 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U850 ( .A1(G2090), .A2(n755), .ZN(n756) );
  XNOR2_X1 U851 ( .A(n756), .B(KEYINPUT100), .ZN(n758) );
  NOR2_X1 U852 ( .A1(n792), .A2(G1971), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U854 ( .A1(n759), .A2(G303), .ZN(n761) );
  AND2_X1 U855 ( .A1(n768), .A2(n761), .ZN(n760) );
  NAND2_X1 U856 ( .A1(n767), .A2(n760), .ZN(n765) );
  INV_X1 U857 ( .A(n761), .ZN(n762) );
  OR2_X1 U858 ( .A1(n762), .A2(G286), .ZN(n763) );
  AND2_X1 U859 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U861 ( .A(n766), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n767), .A2(n768), .ZN(n773) );
  AND2_X1 U863 ( .A1(G8), .A2(n769), .ZN(n770) );
  NOR2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n786) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U868 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n786), .A2(n777), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(n778), .ZN(n780) );
  AND2_X1 U871 ( .A1(n780), .A2(n792), .ZN(n784) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U873 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  NOR2_X1 U874 ( .A1(n792), .A2(n782), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n799) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n1013) );
  NOR2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  NOR2_X1 U878 ( .A1(G1971), .A2(G303), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n1012), .A2(n785), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n527), .A2(n789), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n1012), .A2(KEYINPUT33), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n795) );
  XOR2_X1 U885 ( .A(G1981), .B(G305), .Z(n1002) );
  INV_X1 U886 ( .A(n1002), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U889 ( .A(n800), .B(KEYINPUT102), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n818), .A2(n801), .ZN(n815) );
  XOR2_X1 U891 ( .A(G1986), .B(G290), .Z(n1006) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NAND2_X1 U893 ( .A1(G116), .A2(n899), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G128), .A2(n900), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U896 ( .A(KEYINPUT35), .B(n804), .ZN(n811) );
  XNOR2_X1 U897 ( .A(KEYINPUT92), .B(KEYINPUT34), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n894), .A2(G140), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n895), .A2(G104), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT91), .B(n805), .Z(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U902 ( .A(n809), .B(n808), .Z(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT36), .B(n812), .Z(n889) );
  OR2_X1 U905 ( .A1(n823), .A2(n889), .ZN(n984) );
  NAND2_X1 U906 ( .A1(n1006), .A2(n984), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n825), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n828) );
  XOR2_X1 U909 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n821) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n884), .ZN(n986) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n906), .ZN(n982) );
  NOR2_X1 U913 ( .A1(n816), .A2(n982), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n986), .A2(n819), .ZN(n820) );
  XNOR2_X1 U916 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n822), .A2(n984), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n823), .A2(n889), .ZN(n983) );
  NAND2_X1 U919 ( .A1(n824), .A2(n983), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U923 ( .A(KEYINPUT104), .B(G2454), .ZN(n838) );
  XNOR2_X1 U924 ( .A(G2430), .B(G2435), .ZN(n836) );
  XOR2_X1 U925 ( .A(G2451), .B(G2427), .Z(n831) );
  XNOR2_X1 U926 ( .A(G2438), .B(G2446), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U928 ( .A(n832), .B(G2443), .Z(n834) );
  XNOR2_X1 U929 ( .A(G1348), .B(G1341), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U932 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n839), .A2(G14), .ZN(n920) );
  XNOR2_X1 U934 ( .A(KEYINPUT105), .B(n920), .ZN(G401) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U937 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n843), .A2(n842), .ZN(G188) );
  XOR2_X1 U940 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XNOR2_X1 U941 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  NOR2_X1 U944 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n846), .ZN(G319) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n848) );
  XNOR2_X1 U948 ( .A(KEYINPUT108), .B(G2678), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2096), .B(G2100), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G227) );
  XOR2_X1 U958 ( .A(G1976), .B(G1981), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1966), .B(G1956), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n868) );
  XOR2_X1 U961 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U962 ( .A(G1996), .B(KEYINPUT112), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U964 ( .A(G1971), .B(G1961), .Z(n862) );
  XNOR2_X1 U965 ( .A(G1991), .B(G1986), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U967 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U968 ( .A(KEYINPUT110), .B(G2474), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U971 ( .A1(G124), .A2(n900), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n895), .A2(G100), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G136), .A2(n894), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G112), .A2(n899), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U978 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U979 ( .A1(G118), .A2(n899), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G130), .A2(n900), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n894), .A2(G142), .ZN(n878) );
  XOR2_X1 U983 ( .A(KEYINPUT113), .B(n878), .Z(n880) );
  NAND2_X1 U984 ( .A1(n895), .A2(G106), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U986 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(n884), .ZN(n893) );
  XOR2_X1 U989 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n887) );
  XNOR2_X1 U990 ( .A(n978), .B(KEYINPUT115), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U992 ( .A(n888), .B(G162), .Z(n891) );
  XOR2_X1 U993 ( .A(G164), .B(n889), .Z(n890) );
  XNOR2_X1 U994 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(n893), .B(n892), .Z(n909) );
  NAND2_X1 U996 ( .A1(G139), .A2(n894), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G103), .A2(n895), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U999 ( .A(KEYINPUT114), .B(n898), .ZN(n905) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n899), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n900), .ZN(n901) );
  NAND2_X1 U1002 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1003 ( .A(KEYINPUT47), .B(n903), .Z(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n972) );
  XNOR2_X1 U1005 ( .A(G160), .B(n972), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n1021), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(G171), .B(n1018), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n914), .B(G286), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n918) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(n918), .Z(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n923), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1024 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n1031) );
  INV_X1 U1025 ( .A(KEYINPUT55), .ZN(n995) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n936) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n924) );
  NAND2_X1 U1028 ( .A1(n924), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n926) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n925) );
  NOR2_X1 U1031 ( .A1(n926), .A2(n925), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G1996), .B(G32), .ZN(n929) );
  XNOR2_X1 U1033 ( .A(G27), .B(n927), .ZN(n928) );
  NOR2_X1 U1034 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1035 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1036 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(n934), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1039 ( .A(KEYINPUT119), .B(n937), .Z(n940) );
  XOR2_X1 U1040 ( .A(KEYINPUT54), .B(G34), .Z(n938) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n938), .ZN(n939) );
  NAND2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(n995), .B(n941), .ZN(n943) );
  INV_X1 U1044 ( .A(G29), .ZN(n942) );
  NAND2_X1 U1045 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n944), .ZN(n1001) );
  XNOR2_X1 U1047 ( .A(G20), .B(n945), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(G1341), .B(G19), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(G6), .B(G1981), .ZN(n946) );
  NOR2_X1 U1050 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n952) );
  XOR2_X1 U1052 ( .A(KEYINPUT59), .B(G1348), .Z(n950) );
  XNOR2_X1 U1053 ( .A(G4), .B(n950), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1055 ( .A(n953), .B(KEYINPUT60), .ZN(n956) );
  XOR2_X1 U1056 ( .A(G1966), .B(G21), .Z(n954) );
  XNOR2_X1 U1057 ( .A(KEYINPUT122), .B(n954), .ZN(n955) );
  NAND2_X1 U1058 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1059 ( .A(n957), .B(KEYINPUT123), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n964) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n962) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n959) );
  XNOR2_X1 U1063 ( .A(G1976), .B(G23), .ZN(n958) );
  NOR2_X1 U1064 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1065 ( .A(n960), .B(KEYINPUT124), .ZN(n961) );
  NAND2_X1 U1066 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1067 ( .A(n964), .B(n963), .ZN(n965) );
  NAND2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1069 ( .A(G5), .B(G1961), .ZN(n967) );
  NOR2_X1 U1070 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1071 ( .A(n969), .B(KEYINPUT61), .ZN(n971) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT121), .ZN(n970) );
  NAND2_X1 U1073 ( .A1(n971), .A2(n970), .ZN(n999) );
  XNOR2_X1 U1074 ( .A(G164), .B(G2078), .ZN(n975) );
  XNOR2_X1 U1075 ( .A(G2072), .B(n972), .ZN(n973) );
  XNOR2_X1 U1076 ( .A(n973), .B(KEYINPUT118), .ZN(n974) );
  NAND2_X1 U1077 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1078 ( .A(n976), .B(KEYINPUT50), .ZN(n993) );
  XOR2_X1 U1079 ( .A(G2084), .B(G160), .Z(n977) );
  NOR2_X1 U1080 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1081 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1082 ( .A1(n982), .A2(n981), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n984), .A2(n983), .ZN(n989) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n985) );
  NOR2_X1 U1085 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1086 ( .A(n987), .B(KEYINPUT51), .ZN(n988) );
  NOR2_X1 U1087 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1090 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  NAND2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1092 ( .A1(n997), .A2(G29), .ZN(n998) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1029) );
  XNOR2_X1 U1095 ( .A(G16), .B(KEYINPUT56), .ZN(n1027) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1098 ( .A(KEYINPUT57), .B(n1004), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1005), .B(G1956), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G303), .ZN(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  INV_X1 U1104 ( .A(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT120), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(G1348), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G171), .B(G1961), .ZN(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(G1341), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(n1031), .B(n1030), .ZN(G311) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

