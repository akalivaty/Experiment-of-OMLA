//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  XOR2_X1   g006(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT69), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n205), .A3(KEYINPUT1), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT70), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT70), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n200), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n202), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT65), .A2(G134), .ZN(new_n215));
  NOR2_X1   g029(.A1(KEYINPUT65), .A2(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G137), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n213), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n218), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT65), .A2(G134), .ZN(new_n225));
  AOI21_X1  g039(.A(G137), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n226), .B2(KEYINPUT11), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n228), .A2(new_n218), .A3(G137), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n224), .A2(G137), .A3(new_n225), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT67), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n224), .A2(new_n235), .A3(G137), .A4(new_n225), .ZN(new_n236));
  AOI21_X1  g050(.A(G131), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AND4_X1   g051(.A1(KEYINPUT68), .A2(new_n230), .A3(new_n232), .A4(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n231), .B1(new_n227), .B2(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT68), .B1(new_n239), .B2(new_n237), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n221), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT2), .B(G113), .Z(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n236), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n213), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n217), .A2(KEYINPUT66), .A3(new_n228), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT66), .B1(new_n217), .B2(new_n228), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n232), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n213), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n239), .A2(KEYINPUT68), .A3(new_n237), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n195), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n211), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n256), .B2(new_n195), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n241), .B(new_n245), .C1(new_n255), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n246), .ZN(new_n266));
  OAI21_X1  g080(.A(G131), .B1(new_n251), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n238), .B2(new_n240), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n262), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n245), .B1(new_n269), .B2(new_n241), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n194), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n253), .A2(new_n254), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n263), .B1(new_n274), .B2(new_n267), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n212), .A2(new_n220), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n253), .B2(new_n254), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n241), .C1(new_n255), .C2(new_n263), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n245), .A3(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT72), .B(new_n194), .C1(new_n265), .C2(new_n270), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n192), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT30), .B(new_n241), .C1(new_n255), .C2(new_n263), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n268), .A2(new_n262), .B1(new_n274), .B2(new_n221), .ZN(new_n286));
  XOR2_X1   g100(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(new_n244), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n192), .A3(new_n264), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT31), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n288), .A2(new_n291), .A3(new_n192), .A4(new_n264), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n187), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT32), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(G472), .A3(G902), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n284), .B2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n271), .A2(new_n272), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n281), .A2(new_n273), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n192), .A3(new_n283), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n264), .ZN(new_n303));
  INV_X1    g117(.A(new_n192), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n241), .B1(new_n255), .B2(new_n263), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n244), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n273), .B1(new_n308), .B2(new_n264), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n273), .B2(new_n281), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n192), .A2(KEYINPUT29), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G472), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(new_n297), .C1(new_n284), .C2(new_n293), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n296), .A2(new_n299), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G107), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G104), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n320));
  INV_X1    g134(.A(G104), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G107), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(G104), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G101), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G101), .B1(new_n322), .B2(new_n319), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n212), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n195), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n201), .B1(new_n333), .B2(new_n260), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n334), .A3(new_n330), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n255), .A2(KEYINPUT12), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n335), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n268), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT10), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n210), .A2(new_n211), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n201), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n321), .A2(G107), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n324), .B2(new_n325), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n320), .B1(new_n322), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n348), .B(G101), .C1(new_n350), .C2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(new_n262), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n350), .B2(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n329), .A3(KEYINPUT4), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n335), .A2(KEYINPUT80), .A3(new_n343), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT80), .B1(new_n335), .B2(new_n343), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n347), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n342), .B1(new_n360), .B2(new_n268), .ZN(new_n361));
  INV_X1    g175(.A(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n335), .A2(KEYINPUT80), .A3(new_n343), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n346), .A2(new_n344), .B1(new_n354), .B2(new_n356), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n255), .A2(new_n364), .A3(KEYINPUT81), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n341), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G227), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT78), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G140), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n361), .A2(new_n366), .B1(new_n268), .B2(new_n360), .ZN(new_n375));
  INV_X1    g189(.A(new_n373), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT82), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n360), .A2(new_n268), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n367), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n376), .B1(new_n341), .B2(new_n367), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n381), .B(G469), .C1(new_n385), .C2(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n341), .A2(new_n367), .A3(new_n376), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n376), .B2(new_n375), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n379), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n380), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n331), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n393));
  INV_X1    g207(.A(G116), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n394), .A2(KEYINPUT5), .A3(G119), .ZN(new_n395));
  INV_X1    g209(.A(G113), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n242), .A2(new_n243), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n356), .A2(new_n244), .A3(new_n353), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G125), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n259), .B2(new_n261), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n212), .B2(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n369), .A2(G224), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n416), .A3(new_n406), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n409), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n244), .A2(new_n353), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n419), .A2(new_n356), .B1(new_n392), .B2(new_n401), .ZN(new_n420));
  INV_X1    g234(.A(new_n413), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(KEYINPUT7), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n420), .A2(new_n405), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n329), .A2(KEYINPUT85), .A3(new_n330), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(new_n400), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n405), .B(KEYINPUT8), .Z(new_n426));
  AOI21_X1  g240(.A(new_n426), .B1(new_n424), .B2(new_n400), .ZN(new_n427));
  INV_X1    g241(.A(new_n422), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n425), .A2(new_n427), .B1(new_n413), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n418), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G210), .B1(G237), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n418), .A2(new_n430), .A3(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G214), .B1(G237), .B2(G902), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT83), .Z(new_n438));
  XOR2_X1   g252(.A(new_n438), .B(KEYINPUT84), .Z(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT9), .B(G234), .ZN(new_n440));
  OAI21_X1  g254(.A(G221), .B1(new_n440), .B2(G902), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n391), .A2(new_n436), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT16), .ZN(new_n444));
  INV_X1    g258(.A(G140), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(G125), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(G125), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n410), .A2(G140), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(G146), .B(new_n446), .C1(new_n449), .C2(new_n444), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n448), .A3(new_n197), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n452));
  INV_X1    g266(.A(G119), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(G128), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .A4(new_n208), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(G128), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT76), .B(G110), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(new_n209), .B2(new_n453), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT24), .B(G110), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n450), .B(new_n451), .C1(new_n459), .C2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n446), .B1(new_n449), .B2(new_n444), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n197), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n450), .ZN(new_n466));
  INV_X1    g280(.A(G110), .ZN(new_n467));
  OAI221_X1 g281(.A(new_n466), .B1(new_n460), .B2(new_n461), .C1(new_n457), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT22), .B(G137), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n463), .A2(new_n468), .A3(new_n472), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n389), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT25), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT77), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n476), .B(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(G234), .B2(new_n389), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n474), .A2(new_n475), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n482), .A2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n491));
  OAI21_X1  g305(.A(G131), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n493));
  INV_X1    g307(.A(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n369), .A3(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n199), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n213), .A3(new_n489), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n466), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n492), .A2(KEYINPUT91), .A3(new_n493), .A4(new_n497), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n213), .B1(new_n496), .B2(new_n489), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n321), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n508));
  OAI211_X1 g322(.A(G131), .B(new_n508), .C1(new_n490), .C2(new_n491), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n449), .A2(G146), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n451), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(G131), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n496), .A2(new_n489), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT88), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n509), .A2(new_n511), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n505), .A2(new_n507), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n507), .B1(new_n505), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n389), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G475), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n505), .A2(new_n507), .A3(new_n518), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT89), .ZN(new_n524));
  INV_X1    g338(.A(new_n497), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n503), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n492), .A2(KEYINPUT89), .A3(new_n497), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT19), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT19), .B1(new_n447), .B2(new_n448), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n197), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n526), .A2(new_n450), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(KEYINPUT90), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n507), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT90), .B1(new_n518), .B2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n523), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n536), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n522), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n543));
  INV_X1    g357(.A(new_n540), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT89), .B1(new_n492), .B2(new_n497), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n530), .A2(new_n450), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n527), .B1(new_n515), .B2(new_n517), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n507), .B1(new_n548), .B2(KEYINPUT90), .ZN(new_n549));
  INV_X1    g363(.A(new_n535), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n519), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n538), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n544), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n522), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n543), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G478), .ZN(new_n560));
  INV_X1    g374(.A(G122), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G116), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n394), .A2(G122), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT14), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G107), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT94), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G116), .B(G122), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n564), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n561), .A2(G116), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n318), .B1(new_n571), .B2(KEYINPUT14), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n207), .A2(G143), .A3(new_n208), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n199), .A2(G128), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n215), .A2(new_n216), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n578), .A3(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n318), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n574), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT93), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n199), .A2(KEYINPUT13), .A3(G128), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n575), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G134), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n568), .B(new_n318), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n575), .A2(new_n578), .A3(KEYINPUT93), .A4(new_n576), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n586), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n440), .A2(new_n481), .A3(G953), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(new_n594), .A3(new_n596), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n584), .A2(new_n594), .A3(new_n596), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n584), .B2(new_n594), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n389), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n560), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n560), .B1(new_n600), .B2(KEYINPUT95), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(G234), .A2(G237), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(G952), .A3(new_n369), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G902), .A3(G953), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT21), .B(G898), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n558), .A2(new_n610), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n317), .A2(new_n443), .A3(new_n488), .A4(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  AND3_X1   g434(.A1(new_n278), .A2(new_n245), .A3(new_n280), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n193), .B1(new_n308), .B2(new_n264), .ZN(new_n622));
  OAI22_X1  g436(.A1(new_n621), .A2(KEYINPUT28), .B1(new_n622), .B2(KEYINPUT72), .ZN(new_n623));
  INV_X1    g437(.A(new_n283), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n304), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n290), .A2(new_n292), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(G472), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(KEYINPUT96), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n438), .B1(new_n434), .B2(new_n435), .ZN(new_n632));
  INV_X1    g446(.A(new_n617), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n598), .A2(new_n599), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT33), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G478), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n604), .A2(G478), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(G478), .B2(G902), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n635), .A2(new_n558), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n391), .A2(new_n488), .A3(new_n441), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n631), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT34), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G6));
  INV_X1    g461(.A(new_n644), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n553), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n604), .A2(new_n605), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n636), .A2(KEYINPUT95), .A3(new_n389), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n608), .B1(new_n653), .B2(new_n560), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(G475), .B2(new_n521), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n635), .A2(KEYINPUT97), .A3(new_n650), .A4(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n650), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(new_n634), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n630), .A2(new_n648), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n542), .A2(KEYINPUT92), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n556), .B1(new_n555), .B2(new_n522), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n610), .A2(new_n617), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n473), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n469), .B(new_n669), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n480), .A2(new_n482), .B1(new_n485), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n630), .A2(new_n443), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  XNOR2_X1  g491(.A(new_n612), .B(KEYINPUT99), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(new_n615), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n650), .A2(new_n610), .A3(new_n522), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT100), .ZN(new_n684));
  INV_X1    g498(.A(new_n632), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n391), .A2(new_n441), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n317), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n436), .B(KEYINPUT38), .ZN(new_n691));
  INV_X1    g505(.A(new_n438), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n610), .A3(new_n692), .A4(new_n671), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n391), .A2(new_n441), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n681), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n667), .B(new_n693), .C1(new_n696), .C2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n303), .A2(new_n192), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n265), .A2(new_n270), .ZN(new_n699));
  AOI21_X1  g513(.A(G902), .B1(new_n699), .B2(new_n304), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n628), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n294), .B2(new_n295), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n299), .A2(new_n316), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n697), .B(new_n706), .C1(KEYINPUT40), .C2(new_n696), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  AOI211_X1 g522(.A(new_n641), .B(new_n681), .C1(new_n543), .C2(new_n557), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n317), .A2(new_n688), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  NAND2_X1  g525(.A1(new_n317), .A2(new_n488), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n367), .A2(new_n382), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n373), .ZN(new_n715));
  AOI211_X1 g529(.A(G469), .B(G902), .C1(new_n715), .C2(new_n387), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n379), .B1(new_n388), .B2(new_n389), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n441), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n643), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  AOI21_X1  g537(.A(new_n719), .B1(new_n656), .B2(new_n659), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n718), .A2(new_n727), .A3(new_n441), .A4(new_n632), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n341), .A2(new_n367), .A3(new_n376), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n376), .B1(new_n367), .B2(new_n382), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n389), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n441), .A3(new_n390), .A4(new_n632), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT101), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n673), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n317), .A2(new_n735), .A3(KEYINPUT102), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT102), .B1(new_n317), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n453), .ZN(G21));
  NAND2_X1  g553(.A1(new_n632), .A2(new_n610), .ZN(new_n740));
  NOR4_X1   g554(.A1(new_n719), .A2(new_n667), .A3(new_n617), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT104), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n389), .B1(new_n284), .B2(new_n293), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n290), .B(new_n292), .C1(new_n310), .C2(new_n192), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n187), .B(KEYINPUT103), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n743), .A2(G472), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n742), .B1(new_n746), .B2(new_n488), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n488), .B(new_n748), .C1(new_n627), .C2(new_n628), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(KEYINPUT104), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n741), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  AND2_X1   g566(.A1(new_n733), .A2(KEYINPUT101), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n733), .A2(KEYINPUT101), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n709), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n746), .A2(new_n672), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT105), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n709), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n728), .B2(new_n734), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n748), .B1(new_n627), .B2(new_n628), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n671), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G125), .ZN(G27));
  OAI21_X1  g579(.A(KEYINPUT106), .B1(new_n383), .B2(new_n384), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n377), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(G469), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n379), .A2(new_n389), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n390), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n434), .A2(new_n435), .A3(new_n692), .ZN(new_n774));
  INV_X1    g588(.A(new_n441), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n773), .B1(new_n772), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n709), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n295), .A2(new_n294), .B1(new_n313), .B2(G472), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n487), .B1(new_n781), .B2(new_n298), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT42), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n712), .B2(new_n779), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  INV_X1    g601(.A(new_n778), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT100), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n683), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n487), .B1(new_n684), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n790), .A2(new_n317), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  NAND2_X1  g611(.A1(new_n667), .A2(new_n642), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT43), .Z(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n631), .A3(new_n672), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n774), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(G469), .B1(new_n385), .B2(KEYINPUT45), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n766), .A2(new_n768), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n805), .B1(new_n806), .B2(KEYINPUT45), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n804), .B1(new_n807), .B2(new_n770), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n390), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n807), .A2(new_n804), .A3(new_n770), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n441), .B(new_n695), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n802), .A2(new_n803), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(KEYINPUT111), .B(G137), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(G39));
  INV_X1    g631(.A(new_n317), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n758), .A2(new_n488), .A3(new_n774), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n441), .B1(new_n809), .B2(new_n810), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT47), .B(new_n441), .C1(new_n809), .C2(new_n810), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(new_n445), .ZN(G42));
  NAND3_X1  g640(.A1(new_n488), .A2(new_n439), .A3(new_n441), .ZN(new_n827));
  INV_X1    g641(.A(new_n718), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n798), .B(new_n827), .C1(KEYINPUT49), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT112), .Z(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(KEYINPUT49), .ZN(new_n831));
  OR4_X1    g645(.A1(new_n691), .A2(new_n830), .A3(new_n706), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n299), .A2(new_n316), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n684), .A2(new_n391), .A3(new_n441), .A4(new_n686), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n709), .A2(new_n391), .A3(new_n441), .A4(new_n686), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n835), .A2(new_n781), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n667), .A2(new_n740), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n681), .A2(new_n775), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n772), .A3(new_n671), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n835), .B2(new_n702), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(new_n764), .A3(KEYINPUT52), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(new_n843), .B2(new_n764), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n786), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n751), .B1(new_n736), .B2(new_n737), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n317), .B(new_n488), .C1(new_n724), .C2(new_n720), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n418), .A2(new_n430), .A3(new_n432), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n432), .B1(new_n418), .B2(new_n430), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n633), .B(new_n439), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n558), .A2(new_n642), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n667), .A2(new_n610), .A3(new_n852), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n558), .A2(new_n856), .A3(new_n642), .A4(new_n852), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n630), .A2(new_n858), .A3(new_n648), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n848), .A2(new_n619), .A3(new_n675), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n847), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n681), .B1(new_n521), .B2(G475), .ZN(new_n864));
  INV_X1    g678(.A(new_n649), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n654), .B(new_n864), .C1(new_n865), .C2(new_n541), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n863), .B1(new_n866), .B2(new_n774), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n849), .A2(new_n850), .A3(new_n438), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n607), .A2(new_n609), .A3(new_n864), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT114), .A4(new_n650), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n671), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(new_n441), .A3(new_n391), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n317), .A2(KEYINPUT115), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT115), .B1(new_n317), .B2(new_n872), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n795), .B(new_n793), .C1(new_n778), .C2(new_n777), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n876), .A2(new_n818), .B1(new_n779), .B2(new_n756), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n862), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n317), .A2(new_n872), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n317), .A2(new_n872), .A3(KEYINPUT115), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n780), .A2(new_n761), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(KEYINPUT116), .A3(new_n796), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n861), .A2(new_n878), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n834), .B1(new_n846), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n861), .A2(new_n878), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n786), .A2(KEYINPUT53), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n843), .A2(new_n764), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n843), .A2(new_n764), .A3(KEYINPUT52), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n888), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n834), .B1(new_n783), .B2(new_n785), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n844), .B2(new_n845), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n886), .A3(KEYINPUT117), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n833), .B(new_n887), .C1(new_n896), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n786), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n893), .B2(new_n894), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT53), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n889), .A2(new_n902), .A3(new_n834), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT54), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n900), .A2(KEYINPUT118), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT118), .B1(new_n900), .B2(new_n906), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n719), .A2(new_n774), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n705), .A2(new_n488), .A3(new_n613), .A4(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT120), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n667), .A3(new_n641), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n799), .B(new_n679), .C1(new_n750), .C2(new_n747), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n774), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n823), .A2(new_n824), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n828), .A2(new_n441), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n799), .A2(new_n679), .A3(new_n910), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n761), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n913), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n719), .A2(new_n691), .A3(new_n692), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT50), .Z(new_n924));
  OAI21_X1  g738(.A(new_n909), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT51), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n909), .B(new_n927), .C1(new_n921), .C2(new_n924), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n912), .A2(new_n558), .A3(new_n642), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n753), .A2(new_n754), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n914), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n919), .A2(new_n782), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT48), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n369), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n926), .A2(new_n928), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n907), .A2(new_n908), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(G952), .A2(G953), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n832), .B1(new_n937), .B2(new_n938), .ZN(G75));
  NOR2_X1   g753(.A1(new_n369), .A2(G952), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT122), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT56), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n889), .A2(new_n895), .A3(new_n888), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT117), .B1(new_n898), .B2(new_n886), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n887), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(G902), .ZN(new_n948));
  INV_X1    g762(.A(G210), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n409), .A2(new_n417), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT121), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT55), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(new_n415), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n943), .B(new_n954), .C1(new_n948), .C2(new_n949), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n942), .B1(new_n956), .B2(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n770), .B(KEYINPUT57), .ZN(new_n959));
  INV_X1    g773(.A(new_n900), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n833), .B1(new_n946), .B2(new_n887), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n388), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n944), .A2(new_n945), .B1(new_n903), .B2(new_n834), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(new_n389), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n807), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n940), .B1(new_n963), .B2(new_n966), .ZN(G54));
  AND2_X1   g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n965), .A2(new_n536), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n536), .B1(new_n965), .B2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n940), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT59), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n637), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n960), .B2(new_n961), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n941), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n907), .B2(new_n908), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(new_n637), .ZN(G63));
  NAND2_X1  g793(.A1(G217), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT60), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n947), .A2(new_n670), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n484), .B1(new_n964), .B2(new_n981), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n984), .A3(new_n941), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n983), .A2(new_n984), .A3(KEYINPUT61), .A4(new_n941), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(G66));
  INV_X1    g803(.A(G224), .ZN(new_n990));
  OAI21_X1  g804(.A(G953), .B1(new_n616), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT123), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n861), .B2(G953), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n952), .B1(G898), .B2(new_n369), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G69));
  OAI21_X1  g809(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n528), .A2(new_n529), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(G900), .A2(G953), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n838), .B1(new_n757), .B2(new_n763), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1001));
  INV_X1    g815(.A(new_n796), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n901), .A2(new_n825), .A3(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n813), .A2(new_n839), .A3(new_n782), .A4(new_n814), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1001), .A2(new_n1003), .A3(new_n815), .A4(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n998), .B(new_n999), .C1(new_n1005), .C2(G953), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n558), .A2(new_n642), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n558), .B2(new_n654), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n868), .B1(new_n1008), .B2(KEYINPUT125), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n1009), .B(new_n696), .C1(KEYINPUT125), .C2(new_n1008), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n825), .B1(new_n713), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n815), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1001), .A2(new_n707), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1001), .A2(new_n1015), .A3(new_n707), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1006), .B1(new_n1017), .B2(new_n998), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n369), .B1(G227), .B2(G900), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(new_n1006), .B2(KEYINPUT126), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(G72));
  OR3_X1    g837(.A1(new_n1005), .A2(new_n860), .A3(new_n847), .ZN(new_n1024));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(KEYINPUT63), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT127), .ZN(new_n1027));
  AOI211_X1 g841(.A(new_n192), .B(new_n303), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1014), .A2(new_n861), .A3(new_n1016), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n698), .B1(new_n1029), .B2(new_n1027), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n303), .A2(new_n304), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1026), .B1(new_n1031), .B2(new_n289), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n904), .A2(new_n905), .A3(new_n1032), .ZN(new_n1033));
  NOR4_X1   g847(.A1(new_n1028), .A2(new_n1030), .A3(new_n940), .A4(new_n1033), .ZN(G57));
endmodule


