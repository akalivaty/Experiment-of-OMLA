//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n468), .A2(new_n460), .A3(new_n464), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n473), .B1(new_n477), .B2(new_n464), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n461), .B2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n479), .A2(G137), .A3(new_n464), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(new_n483), .A3(G125), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n472), .A2(new_n478), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G160));
  AND3_X1   g063(.A1(new_n479), .A2(G2105), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n479), .A2(new_n464), .A3(new_n481), .ZN(new_n491));
  INV_X1    g066(.A(G136), .ZN(new_n492));
  OR3_X1    g067(.A1(new_n491), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G100), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT71), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  AND4_X1   g071(.A1(new_n490), .A2(new_n493), .A3(new_n495), .A4(new_n496), .ZN(G162));
  NAND3_X1  g072(.A1(new_n479), .A2(G126), .A3(new_n481), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n464), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n464), .A2(G102), .A3(G2104), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n481), .A3(new_n483), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n479), .A2(KEYINPUT4), .A3(new_n481), .A4(new_n503), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n500), .A2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT73), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n512), .B(new_n514), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT72), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(G88), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(new_n531), .A3(G651), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n519), .A2(new_n522), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(G166));
  NAND2_X1  g109(.A1(new_n521), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n527), .A2(new_n529), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n540), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n515), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT74), .B(G52), .Z(new_n548));
  AOI22_X1  g123(.A1(G651), .A2(new_n547), .B1(new_n521), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT75), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n544), .A2(KEYINPUT75), .A3(new_n549), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(G171));
  NAND2_X1  g128(.A1(new_n540), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT76), .B(G43), .ZN(new_n558));
  AOI22_X1  g133(.A1(G651), .A2(new_n557), .B1(new_n521), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n520), .A2(G53), .A3(G543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n569), .A2(KEYINPUT9), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n515), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n568), .B2(new_n570), .ZN(new_n576));
  INV_X1    g151(.A(G91), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n527), .A2(new_n529), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n572), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  OR2_X1    g155(.A1(new_n533), .A2(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n533), .A2(KEYINPUT78), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT79), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n528), .A2(G74), .ZN(new_n586));
  AOI22_X1  g161(.A1(G651), .A2(new_n586), .B1(new_n521), .B2(G49), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n527), .A2(new_n529), .A3(new_n588), .A4(G87), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n585), .A2(new_n587), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n540), .A2(G86), .B1(G48), .B2(new_n521), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G651), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n515), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n599), .A2(KEYINPUT80), .A3(G651), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n596), .B1(new_n595), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(new_n602), .ZN(G305));
  XOR2_X1   g178(.A(KEYINPUT82), .B(G85), .Z(new_n604));
  NAND2_X1  g179(.A1(new_n540), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n515), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(G651), .A2(new_n608), .B1(new_n521), .B2(G47), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n540), .A2(new_n611), .A3(G92), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G66), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n515), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(G651), .A2(new_n615), .B1(new_n521), .B2(G54), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT10), .B1(new_n578), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n612), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n621));
  NAND4_X1  g196(.A1(new_n612), .A2(new_n621), .A3(new_n618), .A4(new_n616), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n624), .B2(G171), .ZN(G284));
  OAI21_X1  g201(.A(new_n625), .B1(new_n624), .B2(G171), .ZN(G321));
  NAND2_X1  g202(.A1(G299), .A2(new_n624), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G168), .B2(new_n624), .ZN(G280));
  XOR2_X1   g204(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g205(.A(new_n623), .ZN(new_n631));
  XOR2_X1   g206(.A(KEYINPUT85), .B(G559), .Z(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(G860), .B2(new_n632), .ZN(G148));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g212(.A(new_n476), .B1(new_n465), .B2(new_n471), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  INV_X1    g216(.A(new_n491), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n489), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(new_n464), .B2(G111), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2435), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2438), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT14), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(G14), .ZN(G401));
  XOR2_X1   g237(.A(G2067), .B(G2678), .Z(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n665), .B(KEYINPUT86), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n666), .B2(new_n664), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n664), .A2(new_n665), .ZN(new_n672));
  MUX2_X1   g247(.A(new_n672), .B(new_n664), .S(new_n666), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n668), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2096), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n681), .A2(new_n683), .A3(new_n685), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n688), .B(new_n689), .C1(new_n687), .C2(new_n686), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(G1986), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT22), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  NAND2_X1  g271(.A1(new_n642), .A2(G141), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n489), .A2(G129), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT26), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G105), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n468), .A2(new_n464), .A3(new_n469), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT70), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n702), .B1(new_n704), .B2(new_n470), .ZN(new_n705));
  OAI21_X1  g280(.A(G29), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT27), .B(G1996), .Z(new_n712));
  NAND2_X1  g287(.A1(G162), .A2(G29), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G29), .B2(G35), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT29), .B(G2090), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n711), .A2(new_n712), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G299), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT100), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT23), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1956), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT91), .B(G2067), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n728));
  INV_X1    g303(.A(G26), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G29), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n642), .A2(G140), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT90), .ZN(new_n733));
  OR2_X1    g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G116), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n467), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n489), .A2(G128), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n731), .B1(new_n738), .B2(G29), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n727), .B(new_n730), .C1(new_n739), .C2(new_n728), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n719), .A2(G4), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n631), .B2(new_n719), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G1348), .ZN(new_n743));
  AND4_X1   g318(.A1(new_n717), .A2(new_n725), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(KEYINPUT24), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(KEYINPUT24), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n707), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n707), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT94), .Z(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G2084), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n711), .A2(new_n712), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G33), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n642), .A2(G139), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n755), .B(new_n758), .C1(new_n464), .C2(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  OAI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(new_n707), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n750), .A2(G2084), .B1(new_n762), .B2(G2072), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n730), .B1(new_n739), .B2(new_n728), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(new_n726), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n744), .A2(new_n753), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G5), .A2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G171), .B2(G16), .ZN(new_n768));
  MUX2_X1   g343(.A(new_n767), .B(new_n768), .S(KEYINPUT97), .Z(new_n769));
  OAI22_X1  g344(.A1(new_n769), .A2(G1961), .B1(new_n714), .B2(new_n716), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n719), .A2(G19), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n561), .B2(new_n719), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  INV_X1    g348(.A(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT99), .B1(new_n774), .B2(G29), .ZN(new_n775));
  OR3_X1    g350(.A1(new_n774), .A2(KEYINPUT99), .A3(G29), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n775), .B(new_n776), .C1(G164), .C2(new_n707), .ZN(new_n777));
  INV_X1    g352(.A(G2078), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n766), .A2(new_n770), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n762), .A2(G2072), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G22), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G166), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1971), .ZN(new_n786));
  MUX2_X1   g361(.A(G6), .B(G305), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT88), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n787), .A2(new_n789), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G23), .ZN(new_n793));
  NAND2_X1  g368(.A1(G288), .A2(KEYINPUT89), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT89), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n585), .A2(new_n795), .A3(new_n587), .A4(new_n589), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n793), .B1(new_n797), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n792), .A2(KEYINPUT34), .A3(new_n800), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G290), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G16), .B2(G24), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n707), .A2(G25), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n642), .A2(G131), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n489), .A2(G119), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n707), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT87), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n808), .A2(new_n809), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n810), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n783), .B1(new_n805), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g400(.A(KEYINPUT36), .B(new_n823), .C1(new_n803), .C2(new_n804), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n781), .B(new_n782), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n769), .A2(G1961), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT30), .B(G28), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n829), .A2(new_n707), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n647), .B2(new_n707), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT96), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n719), .A2(G21), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G168), .B2(new_n719), .ZN(new_n836));
  INV_X1    g411(.A(G1966), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n828), .A2(new_n834), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT98), .Z(new_n840));
  NOR2_X1   g415(.A1(new_n742), .A2(G1348), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n827), .A2(new_n840), .A3(new_n841), .ZN(G311));
  NOR2_X1   g417(.A1(new_n825), .A2(new_n826), .ZN(new_n843));
  INV_X1    g418(.A(new_n781), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n840), .ZN(new_n846));
  INV_X1    g421(.A(new_n841), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n782), .ZN(G150));
  NAND2_X1  g423(.A1(new_n540), .A2(G93), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n515), .B2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(G651), .A2(new_n852), .B1(new_n521), .B2(G55), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n631), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n561), .B1(new_n856), .B2(new_n857), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n560), .B1(new_n849), .B2(new_n853), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n863), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT102), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n859), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n861), .B1(new_n870), .B2(new_n872), .ZN(G145));
  XNOR2_X1  g448(.A(G160), .B(new_n647), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G162), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n738), .A2(G164), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n701), .A2(new_n705), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n738), .A2(G164), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n761), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(new_n760), .A3(new_n880), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT103), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n639), .B(new_n816), .ZN(new_n887));
  INV_X1    g462(.A(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(new_n464), .B2(G118), .ZN(new_n890));
  OAI22_X1  g465(.A1(new_n491), .A2(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(G130), .B2(new_n489), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n887), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n884), .A2(new_n894), .A3(new_n760), .A4(new_n880), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n886), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n886), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n876), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n886), .A2(new_n895), .ZN(new_n899));
  INV_X1    g474(.A(new_n893), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n886), .A2(new_n893), .A3(new_n895), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n875), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT40), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n898), .A2(new_n903), .A3(new_n907), .A4(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(G395));
  XNOR2_X1  g484(.A(new_n634), .B(new_n866), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n619), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n619), .A2(G299), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n912), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  INV_X1    g495(.A(new_n797), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n533), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n797), .A2(G166), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G305), .B(G290), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n925), .A3(new_n923), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n916), .A2(new_n931), .A3(new_n918), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n920), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n920), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g511(.A(new_n935), .B1(G868), .B2(new_n858), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  INV_X1    g513(.A(new_n865), .ZN(new_n939));
  INV_X1    g514(.A(new_n857), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT101), .B1(new_n849), .B2(new_n853), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n560), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n552), .ZN(new_n943));
  OAI21_X1  g518(.A(G168), .B1(new_n943), .B2(new_n550), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n551), .A2(G286), .A3(new_n552), .ZN(new_n945));
  AND4_X1   g520(.A1(new_n939), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n939), .A2(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n917), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n943), .A2(G168), .A3(new_n550), .ZN(new_n949));
  AOI21_X1  g524(.A(G286), .B1(new_n551), .B2(new_n552), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n949), .A2(new_n950), .B1(new_n864), .B2(new_n865), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n942), .A2(new_n944), .A3(new_n939), .A4(new_n945), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n951), .B(new_n952), .C1(new_n914), .C2(new_n913), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n948), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n929), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n927), .A2(new_n928), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(new_n954), .A3(new_n948), .A4(new_n953), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n958), .A3(new_n904), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n956), .A2(new_n958), .A3(new_n962), .A4(new_n904), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n938), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT106), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(KEYINPUT44), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n738), .B(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n878), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n500), .B2(new_n508), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT68), .B1(new_n485), .B2(G2105), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n473), .B(new_n464), .C1(new_n484), .C2(new_n474), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G101), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n704), .B2(new_n470), .ZN(new_n984));
  INV_X1    g559(.A(new_n482), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n982), .A2(new_n986), .A3(G40), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n979), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n975), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n816), .B(new_n820), .Z(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n988), .A2(new_n974), .A3(new_n878), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT107), .Z(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(G290), .B(G1986), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n591), .C1(new_n601), .C2(new_n602), .ZN(new_n998));
  XOR2_X1   g573(.A(KEYINPUT111), .B(G86), .Z(new_n999));
  NAND3_X1  g574(.A1(new_n527), .A2(new_n529), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n521), .A2(G48), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1000), .A2(KEYINPUT112), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT112), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n595), .A2(new_n600), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n998), .B1(new_n1005), .B2(new_n997), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n987), .B2(new_n977), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n998), .B(KEYINPUT49), .C1(new_n1005), .C2(new_n997), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n794), .B2(new_n796), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n1014), .B2(new_n1009), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1013), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1010), .B(new_n1016), .C1(new_n921), .C2(new_n1013), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  INV_X1    g594(.A(G40), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n487), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT45), .B(new_n976), .C1(new_n500), .C2(new_n508), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n979), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n1024));
  INV_X1    g599(.A(G1971), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n977), .A2(KEYINPUT50), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT109), .B(G2090), .Z(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n976), .C1(new_n500), .C2(new_n508), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1021), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT110), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1019), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(G303), .B2(G8), .ZN(new_n1037));
  AOI211_X1 g612(.A(KEYINPUT55), .B(new_n1019), .C1(new_n581), .C2(new_n582), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1018), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(new_n1033), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1042), .A2(new_n1019), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n987), .B1(KEYINPUT50), .B2(new_n977), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n1045));
  INV_X1    g620(.A(G2084), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1032), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1023), .A2(new_n837), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1021), .A2(new_n1029), .A3(new_n1046), .A4(new_n1032), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT114), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1051), .A2(G8), .A3(G168), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1040), .A2(KEYINPUT115), .A3(new_n1043), .A4(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1041), .A2(KEYINPUT108), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1021), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT110), .A3(new_n1030), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1033), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1039), .A3(G8), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1054), .A2(new_n1062), .A3(new_n1052), .A4(new_n1043), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT63), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1053), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1068), .A2(new_n1040), .A3(KEYINPUT63), .A4(new_n1052), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1062), .A2(new_n1018), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n998), .B1(new_n1072), .B2(G288), .ZN(new_n1073));
  XOR2_X1   g648(.A(new_n1009), .B(KEYINPUT113), .Z(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1054), .A2(new_n1062), .A3(new_n1043), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT124), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1047), .A2(G168), .A3(new_n1050), .A4(new_n1048), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(G8), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1051), .A2(G286), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1080), .A2(G8), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n979), .A2(new_n1022), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT53), .A3(new_n778), .A4(new_n1021), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1023), .B2(G2078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1021), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1092));
  INV_X1    g667(.A(G1961), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1095), .A2(new_n1096), .A3(G171), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1095), .B2(G171), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1080), .A2(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(KEYINPUT51), .B2(new_n1082), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1101), .B(KEYINPUT62), .C1(new_n1103), .C2(new_n1081), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1087), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1056), .A2(G1956), .B1(new_n1023), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G299), .A2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT57), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT61), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1110), .B(KEYINPUT57), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1088), .A2(new_n1021), .A3(new_n1106), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1092), .A2(new_n724), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1114), .A2(new_n1115), .A3(KEYINPUT61), .A4(new_n1116), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n987), .A2(G2067), .A3(new_n977), .ZN(new_n1121));
  INV_X1    g696(.A(G1348), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1092), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n623), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n631), .A2(KEYINPUT60), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(KEYINPUT58), .B(G1341), .Z(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n987), .B2(new_n977), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(G1996), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1021), .A2(new_n979), .A3(new_n1022), .A4(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT119), .B(new_n1129), .C1(new_n987), .C2(new_n977), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1137));
  AND3_X1   g712(.A1(new_n1136), .A2(new_n561), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1136), .B2(new_n561), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1120), .A2(new_n1128), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1117), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(new_n1123), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1114), .B(KEYINPUT117), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n631), .B1(new_n1144), .B2(new_n1108), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1085), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1095), .A2(G171), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT121), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT54), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1095), .A2(new_n1096), .A3(G171), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1094), .A2(KEYINPUT122), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1092), .A2(new_n1153), .A3(new_n1093), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1020), .B1(new_n485), .B2(G2105), .ZN(new_n1156));
  NOR4_X1   g731(.A1(new_n984), .A2(new_n985), .A3(new_n1090), .A4(G2078), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n979), .A2(new_n1022), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1155), .A2(G301), .A3(new_n1091), .A4(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1095), .A2(G301), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1155), .A2(new_n1091), .A3(new_n1160), .ZN(new_n1164));
  OAI211_X1 g739(.A(KEYINPUT54), .B(new_n1163), .C1(new_n1164), .C2(G301), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1146), .A2(new_n1147), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1078), .B1(new_n1105), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n996), .B1(new_n1076), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n733), .A2(new_n972), .A3(new_n737), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n989), .A2(new_n993), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n817), .A2(new_n820), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(KEYINPUT126), .B(new_n1170), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1175), .A2(new_n988), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n973), .A2(new_n878), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n988), .ZN(new_n1179));
  NAND2_X1  g754(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1180));
  NOR2_X1   g755(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n988), .B2(new_n974), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n988), .A2(new_n974), .A3(new_n1181), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1179), .B(new_n1180), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n1184), .B(KEYINPUT47), .Z(new_n1185));
  NAND3_X1  g760(.A1(new_n988), .A2(new_n809), .A3(new_n806), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT48), .Z(new_n1187));
  NOR2_X1   g762(.A1(new_n994), .A2(new_n1187), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1177), .A2(new_n1185), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1169), .A2(new_n1189), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g765(.A1(G401), .A2(G229), .A3(G227), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n905), .A2(G319), .A3(new_n967), .A4(new_n1192), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


