//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT64), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n203), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n201), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n210), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n211), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G20), .B2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n211), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n257), .A2(G150), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(KEYINPUT68), .B1(G20), .B2(new_n204), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n252), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n251), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(G50), .B1(new_n211), .B2(G1), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(G50), .B2(new_n269), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  OAI21_X1  g0077(.A(G274), .B1(new_n277), .B2(new_n210), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AND2_X1   g0082(.A1(G1), .A2(G13), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n280), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT66), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n284), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n280), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(G226), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G222), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n295), .B1(new_n224), .B2(new_n293), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n289), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G200), .B2(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n276), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT10), .B1(new_n304), .B2(KEYINPUT72), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n306), .ZN(new_n308));
  INV_X1    g0108(.A(new_n301), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n275), .B1(new_n309), .B2(G169), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(KEYINPUT69), .B1(new_n311), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(KEYINPUT69), .B2(new_n310), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n288), .B1(G244), .B2(new_n291), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT70), .A2(G107), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n296), .A2(new_n219), .B1(new_n319), .B2(new_n293), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G232), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n324), .A2(new_n325), .A3(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n299), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n314), .A2(G190), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT15), .B(G87), .Z(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n262), .B1(new_n211), .B2(new_n224), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n254), .A2(new_n256), .ZN(new_n332));
  INV_X1    g0132(.A(new_n261), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n251), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G77), .B1(new_n211), .B2(G1), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n335), .B1(G77), .B2(new_n269), .C1(new_n272), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n314), .A2(new_n327), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G200), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n314), .A2(new_n327), .A3(KEYINPUT71), .A4(new_n311), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(G169), .B1(new_n314), .B2(new_n327), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(new_n338), .B2(G179), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n328), .A2(new_n339), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n307), .A2(new_n308), .A3(new_n313), .A4(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n332), .A2(new_n201), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n262), .A2(new_n224), .B1(new_n211), .B2(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n251), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT11), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n269), .B2(G68), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT12), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n203), .B1(new_n268), .B2(G20), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n356), .A2(new_n357), .B1(new_n271), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n351), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n285), .A2(KEYINPUT66), .A3(new_n286), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n291), .A2(G238), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n321), .A2(new_n323), .A3(G226), .A4(new_n294), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n321), .A2(new_n323), .A3(G232), .A4(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G97), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n369), .C1(new_n253), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n299), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n372), .A2(new_n367), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n363), .A2(KEYINPUT73), .B1(G238), .B2(new_n291), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT14), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(G169), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n374), .A2(new_n378), .A3(G179), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n379), .B2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n360), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n360), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n379), .B2(new_n302), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n374), .B2(new_n378), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n333), .B1(new_n268), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n271), .B1(new_n270), .B2(new_n333), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G58), .A2(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n207), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(G159), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n332), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  AND2_X1   g0202(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n403), .A2(new_n404), .A3(new_n253), .ZN(new_n405));
  INV_X1    g0205(.A(new_n321), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n402), .B(new_n211), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT75), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n322), .ZN(new_n410));
  NAND2_X1  g0210(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G33), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(G20), .B1(new_n412), .B2(new_n321), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n402), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n401), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n402), .A2(G20), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n253), .B1(new_n403), .B2(new_n404), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n323), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n324), .B2(new_n211), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n399), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT16), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT76), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n415), .B(new_n251), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(G33), .B1(new_n410), .B2(new_n411), .ZN(new_n426));
  INV_X1    g0226(.A(new_n323), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n416), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n402), .B1(new_n293), .B2(G20), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n399), .B1(new_n430), .B2(G68), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n431), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n394), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n281), .A2(new_n287), .B1(new_n325), .B2(new_n290), .ZN(new_n434));
  AND2_X1   g0234(.A1(G226), .A2(G1698), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n412), .A2(new_n321), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT77), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n412), .A2(new_n438), .A3(new_n321), .A4(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G87), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n412), .A2(G223), .A3(new_n294), .A4(new_n321), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n437), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n434), .B1(new_n442), .B2(new_n299), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G179), .ZN(new_n444));
  INV_X1    g0244(.A(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n443), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT18), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n433), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n443), .A2(G200), .ZN(new_n452));
  AOI211_X1 g0252(.A(G190), .B(new_n434), .C1(new_n442), .C2(new_n299), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n433), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n443), .A2(new_n302), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(G200), .B2(new_n443), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT76), .B1(new_n431), .B2(KEYINPUT16), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n423), .A2(new_n424), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n203), .B1(new_n413), .B2(new_n402), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n403), .A2(new_n404), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n406), .B1(new_n461), .B2(G33), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT7), .B1(new_n462), .B2(G20), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n252), .B1(new_n464), .B2(new_n401), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n457), .A2(KEYINPUT17), .A3(new_n394), .A4(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n448), .A2(new_n450), .A3(new_n455), .A4(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n346), .A2(new_n392), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT83), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G257), .A2(G1698), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(new_n227), .B2(G1698), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(new_n412), .A3(new_n321), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n324), .A2(G303), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n289), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G270), .A3(new_n289), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n285), .A2(new_n482), .A3(new_n477), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n475), .A2(new_n484), .A3(new_n311), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n211), .C1(G33), .C2(new_n370), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n251), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n487), .A2(KEYINPUT20), .A3(new_n251), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n268), .A2(G13), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n268), .A2(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n269), .A2(new_n497), .A3(new_n210), .A4(new_n250), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n500), .A3(G116), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT82), .B1(new_n498), .B2(new_n488), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n494), .A2(new_n496), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n470), .B1(new_n485), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n481), .A2(new_n483), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n462), .A2(new_n472), .B1(G303), .B2(new_n324), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n289), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n503), .A2(new_n509), .A3(KEYINPUT21), .A4(G169), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n485), .A2(new_n503), .A3(new_n470), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n505), .A2(new_n506), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT84), .B1(new_n513), .B2(new_n504), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n503), .A2(new_n509), .A3(G169), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n503), .B1(G200), .B2(new_n509), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n302), .B2(new_n509), .ZN(new_n519));
  AND4_X1   g0319(.A1(new_n512), .A2(new_n514), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G250), .A2(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G257), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n412), .A3(new_n321), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G294), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n289), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n480), .A2(new_n289), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n227), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n483), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n445), .ZN(new_n531));
  INV_X1    g0331(.A(new_n483), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n311), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n412), .A2(KEYINPUT22), .A3(G87), .A4(new_n321), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n211), .B1(new_n318), .B2(KEYINPUT23), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT22), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n324), .B2(new_n220), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n538), .B1(new_n535), .B2(new_n536), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT24), .B1(new_n549), .B2(new_n546), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n252), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  XOR2_X1   g0351(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n552));
  NOR2_X1   g0352(.A1(new_n269), .A2(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n498), .A2(new_n226), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n531), .B(new_n534), .C1(new_n551), .C2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n541), .B1(new_n540), .B2(new_n547), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n549), .A2(new_n546), .A3(KEYINPUT24), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n251), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n524), .A2(new_n525), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n299), .ZN(new_n563));
  INV_X1    g0363(.A(new_n528), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n564), .A3(new_n302), .A4(new_n483), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n533), .B2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n566), .A3(new_n556), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n319), .B1(new_n428), .B2(new_n429), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT6), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n569), .A2(new_n370), .A3(G107), .ZN(new_n570));
  XNOR2_X1  g0370(.A(G97), .B(G107), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(new_n211), .B1(new_n224), .B2(new_n332), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n251), .B1(new_n568), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n498), .A2(G97), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G97), .B2(new_n270), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT78), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n578), .C1(G97), .C2(new_n270), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n483), .B1(new_n527), .B2(new_n522), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(KEYINPUT4), .A2(G244), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n321), .A2(new_n323), .A3(new_n584), .A4(new_n294), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n321), .A2(new_n323), .A3(G250), .A4(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n486), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n462), .A2(G244), .A3(new_n294), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n311), .B(new_n583), .C1(new_n590), .C2(new_n289), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n412), .A2(new_n321), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n294), .A2(G244), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n587), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n289), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n445), .B1(new_n596), .B2(new_n582), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n581), .A2(new_n591), .A3(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(G190), .B(new_n583), .C1(new_n590), .C2(new_n289), .ZN(new_n599));
  OAI21_X1  g0399(.A(G200), .B1(new_n596), .B2(new_n582), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n574), .A4(new_n580), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n558), .A2(new_n567), .A3(new_n598), .A4(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G87), .A2(G97), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n316), .A2(new_n604), .A3(new_n317), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n211), .B1(new_n253), .B2(new_n370), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n262), .A2(KEYINPUT19), .A3(new_n370), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n211), .A2(G68), .ZN(new_n609));
  OAI22_X1  g0409(.A1(new_n607), .A2(new_n608), .B1(new_n592), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI221_X1 g0412(.A(KEYINPUT81), .B1(new_n592), .B2(new_n609), .C1(new_n607), .C2(new_n608), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n251), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n329), .A2(new_n269), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n499), .A2(new_n329), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(G238), .A2(G1698), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n225), .B2(G1698), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n412), .A3(new_n321), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G116), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n299), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n289), .B(G250), .C1(G1), .C2(new_n476), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n285), .A2(new_n477), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n445), .B1(new_n624), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n289), .B1(new_n621), .B2(new_n622), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n630), .A2(new_n311), .A3(new_n627), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT80), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n630), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G179), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT80), .ZN(new_n635));
  OAI21_X1  g0435(.A(G169), .B1(new_n630), .B2(new_n627), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n618), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n624), .A2(G190), .A3(new_n628), .ZN(new_n639));
  OAI21_X1  g0439(.A(G200), .B1(new_n630), .B2(new_n627), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n498), .A2(new_n220), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n641), .A2(new_n643), .A3(new_n616), .A4(new_n614), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n602), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n469), .A2(new_n520), .A3(new_n646), .ZN(G372));
  AND3_X1   g0447(.A1(new_n433), .A2(new_n449), .A3(new_n446), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n449), .B1(new_n433), .B2(new_n446), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n341), .A2(new_n344), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n385), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n455), .A2(new_n467), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n391), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n307), .A3(new_n308), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n313), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n567), .A2(new_n598), .A3(new_n601), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n634), .A2(new_n636), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n618), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n644), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT86), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n601), .A2(new_n598), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n252), .B1(new_n610), .B2(new_n611), .ZN(new_n664));
  AOI211_X1 g0464(.A(new_n642), .B(new_n615), .C1(new_n664), .C2(new_n613), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n641), .B1(new_n618), .B2(new_n659), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT86), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n663), .A2(new_n666), .A3(new_n667), .A4(new_n567), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n513), .A2(new_n504), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n517), .A3(new_n558), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n662), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n660), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n661), .B2(new_n598), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n581), .A2(new_n591), .A3(new_n597), .ZN(new_n675));
  XNOR2_X1  g0475(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n638), .A2(new_n644), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n672), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n469), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n657), .A2(new_n681), .ZN(G369));
  NAND2_X1  g0482(.A1(new_n669), .A2(new_n517), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n268), .A2(new_n211), .A3(G13), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n684), .B2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n503), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT89), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n683), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n514), .A2(new_n517), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n512), .A3(new_n519), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n696), .B2(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT90), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n699), .B(new_n694), .C1(new_n696), .C2(new_n693), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(G330), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n691), .B1(new_n551), .B2(new_n557), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n567), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n558), .ZN(new_n704));
  INV_X1    g0504(.A(new_n558), .ZN(new_n705));
  INV_X1    g0505(.A(new_n691), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n691), .B1(new_n695), .B2(new_n512), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n711), .A2(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n605), .A2(G116), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n215), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n715), .A2(new_n268), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT91), .ZN(new_n719));
  INV_X1    g0519(.A(new_n208), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n718), .A2(new_n719), .B1(new_n720), .B2(new_n717), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n719), .B2(new_n718), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  AOI211_X1 g0523(.A(KEYINPUT29), .B(new_n691), .C1(new_n671), .C2(new_n679), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n514), .A2(new_n512), .A3(new_n517), .A4(new_n558), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n663), .A3(new_n567), .A4(new_n666), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n638), .A2(new_n644), .A3(new_n675), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n676), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n666), .A2(KEYINPUT26), .A3(new_n675), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n672), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n726), .B1(new_n730), .B2(KEYINPUT92), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT92), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n732), .B(new_n672), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n706), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n724), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n520), .A2(new_n646), .A3(new_n706), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n633), .A2(new_n529), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n596), .A2(new_n582), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n485), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n737), .A2(KEYINPUT30), .A3(new_n485), .A4(new_n738), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n738), .A2(new_n533), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n475), .A2(new_n484), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n633), .A3(G179), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n691), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n739), .A2(new_n740), .B1(new_n743), .B2(new_n745), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n706), .B1(new_n751), .B2(new_n742), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT31), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n736), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G330), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n735), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n723), .B1(new_n757), .B2(G1), .ZN(G364));
  NAND2_X1  g0558(.A1(new_n211), .A2(G13), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n268), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n717), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n701), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n698), .A2(new_n700), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(G330), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n210), .B1(G20), .B2(new_n445), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n462), .A2(new_n716), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n248), .A2(new_n476), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n476), .C2(new_n209), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n716), .A2(new_n324), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT93), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G355), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G116), .B2(new_n215), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n772), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n763), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n211), .A2(new_n311), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n302), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n211), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n293), .B1(new_n785), .B2(new_n224), .C1(new_n787), .C2(new_n370), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G190), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n783), .A2(G190), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G68), .A2(new_n790), .B1(new_n792), .B2(G50), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n211), .A2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n220), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n783), .A2(G190), .A3(new_n388), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  AOI211_X1 g0598(.A(new_n788), .B(new_n796), .C1(G58), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n794), .A2(new_n784), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n800), .A2(KEYINPUT95), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(KEYINPUT95), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n398), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n794), .A2(new_n302), .A3(G200), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT96), .Z(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G107), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n799), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT97), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n790), .ZN(new_n812));
  OR2_X1    g0612(.A1(KEYINPUT33), .A2(G317), .ZN(new_n813));
  NAND2_X1  g0613(.A1(KEYINPUT33), .A2(G317), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n787), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G294), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  INV_X1    g0618(.A(G322), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n324), .B1(new_n785), .B2(new_n818), .C1(new_n819), .C2(new_n797), .ZN(new_n820));
  INV_X1    g0620(.A(new_n803), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(G329), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n792), .A2(G326), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n795), .B(KEYINPUT98), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n807), .A2(G283), .B1(G303), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n817), .A2(new_n822), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n809), .A2(new_n810), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n811), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n782), .B1(new_n828), .B2(new_n771), .ZN(new_n829));
  INV_X1    g0629(.A(new_n770), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n697), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g0631(.A1(new_n767), .A2(KEYINPUT99), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(KEYINPUT99), .B1(new_n767), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  AOI21_X1  g0635(.A(new_n691), .B1(new_n671), .B2(new_n679), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n344), .A2(new_n340), .A3(new_n337), .A4(new_n691), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n337), .A2(new_n691), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n345), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n836), .B(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n755), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n764), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n768), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n771), .A2(new_n768), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n763), .B1(G77), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n324), .B1(new_n785), .B2(new_n488), .C1(new_n849), .C2(new_n797), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n821), .B2(G311), .ZN(new_n851));
  INV_X1    g0651(.A(G283), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n812), .A2(new_n852), .B1(new_n370), .B2(new_n787), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G303), .B2(new_n792), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n807), .A2(G87), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n824), .A2(G107), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n851), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n785), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n792), .A2(G137), .B1(new_n858), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  INV_X1    g0660(.A(new_n798), .ZN(new_n861));
  INV_X1    g0661(.A(G143), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n859), .B1(new_n860), .B2(new_n812), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n462), .B1(new_n202), .B2(new_n787), .ZN(new_n866));
  INV_X1    g0666(.A(new_n807), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n203), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(G132), .C2(new_n821), .ZN(new_n869));
  INV_X1    g0669(.A(new_n824), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n865), .B(new_n869), .C1(new_n201), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n864), .A2(KEYINPUT34), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n857), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n848), .B1(new_n873), .B2(new_n771), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  INV_X1    g0676(.A(new_n572), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n212), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  NAND3_X1  g0681(.A1(new_n720), .A2(G77), .A3(new_n395), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n268), .B(G13), .C1(new_n882), .C2(new_n244), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n373), .A2(KEYINPUT13), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n886));
  OAI21_X1  g0686(.A(G169), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT14), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n382), .A3(new_n381), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n360), .A3(new_n706), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n415), .A2(new_n251), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT16), .B1(new_n464), .B2(new_n422), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n394), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n689), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT100), .B(new_n394), .C1(new_n892), .C2(new_n893), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n653), .B2(new_n650), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n433), .A2(new_n897), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n466), .B(new_n394), .C1(new_n453), .C2(new_n452), .ZN(new_n903));
  AND4_X1   g0703(.A1(new_n901), .A2(new_n447), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n444), .B(new_n689), .C1(new_n445), .C2(new_n443), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n896), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n906), .B2(new_n903), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n891), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n447), .A2(new_n902), .A3(new_n901), .A4(new_n903), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n906), .A2(new_n903), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n901), .ZN(new_n912));
  INV_X1    g0712(.A(new_n899), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n468), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(KEYINPUT101), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT101), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(new_n891), .C1(new_n900), .C2(new_n908), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n447), .A2(new_n902), .A3(new_n903), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(new_n901), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n902), .B1(new_n653), .B2(new_n650), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n891), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n915), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n890), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n839), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n680), .A2(new_n706), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n651), .A2(new_n691), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n360), .A2(new_n691), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n385), .A2(new_n391), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n360), .B(new_n691), .C1(new_n889), .C2(new_n390), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n916), .A2(new_n931), .A3(new_n918), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n689), .B1(new_n648), .B2(new_n649), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n469), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n657), .B1(new_n735), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT102), .B1(new_n752), .B2(KEYINPUT31), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT102), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n748), .A2(new_n944), .A3(new_n749), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n736), .A2(new_n753), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n839), .B1(new_n933), .B2(new_n934), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n916), .A2(new_n918), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n923), .B2(new_n915), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n469), .A2(new_n946), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(G330), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n942), .A2(new_n957), .B1(new_n268), .B2(new_n760), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n942), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n884), .B1(new_n958), .B2(new_n959), .ZN(G367));
  INV_X1    g0760(.A(KEYINPUT42), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n695), .A2(new_n512), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n962), .A2(new_n558), .A3(new_n706), .A4(new_n704), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n581), .A2(new_n691), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n663), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n675), .A2(new_n691), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n961), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n708), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n970), .A2(new_n711), .A3(KEYINPUT42), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n598), .B1(new_n965), .B2(new_n558), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n706), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n665), .A2(new_n706), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n672), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n661), .B2(new_n976), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n975), .A2(KEYINPUT43), .A3(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT103), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n978), .B(KEYINPUT43), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT104), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n710), .A2(new_n968), .ZN(new_n984));
  AND3_X1   g0784(.A1(new_n980), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(new_n980), .B2(new_n983), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n717), .B(KEYINPUT41), .Z(new_n988));
  NAND3_X1  g0788(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n963), .A2(new_n707), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n991), .B2(new_n968), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(KEYINPUT44), .A3(new_n968), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n712), .B2(new_n967), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n989), .A2(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n710), .B1(new_n996), .B2(KEYINPUT105), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n989), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n993), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT105), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n1001), .A3(new_n709), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n970), .A2(new_n711), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT106), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n963), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n701), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n698), .A2(new_n1006), .A3(G330), .A4(new_n700), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1004), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1008), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n756), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT107), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1003), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1012), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n757), .B1(new_n1016), .B2(new_n1010), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n997), .A2(new_n1002), .ZN(new_n1018));
  OAI21_X1  g0818(.A(KEYINPUT107), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n988), .B1(new_n1020), .B2(new_n757), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n987), .B1(new_n1021), .B2(new_n762), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n772), .B1(new_n215), .B2(new_n330), .C1(new_n774), .C2(new_n239), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(new_n763), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n795), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n1025), .B2(G116), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n462), .B(new_n1026), .C1(G283), .C2(new_n858), .ZN(new_n1027));
  INV_X1    g0827(.A(G317), .ZN(new_n1028));
  INV_X1    g0828(.A(G303), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n803), .C1(new_n861), .C2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n824), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n816), .A2(new_n318), .B1(new_n790), .B2(G294), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n806), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G311), .A2(new_n792), .B1(new_n1033), .B2(G97), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n787), .A2(new_n203), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n202), .B2(new_n795), .C1(new_n862), .C2(new_n791), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n293), .B1(new_n785), .B2(new_n201), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n797), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1039), .B1(G150), .B2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n790), .A2(G159), .B1(new_n1033), .B2(G77), .ZN(new_n1042));
  INV_X1    g0842(.A(G137), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1041), .B(new_n1042), .C1(new_n803), .C2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1030), .A2(new_n1035), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT47), .Z(new_n1046));
  INV_X1    g0846(.A(new_n771), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1024), .B1(new_n830), .B2(new_n978), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1022), .A2(new_n1048), .ZN(G387));
  AOI21_X1  g0849(.A(new_n761), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n236), .A2(new_n476), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1051), .A2(new_n773), .B1(new_n715), .B2(new_n778), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n261), .A2(new_n201), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n476), .B1(new_n203), .B2(new_n224), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1054), .A2(new_n715), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1052), .A2(new_n1056), .B1(G107), .B2(new_n215), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n764), .B1(new_n1057), .B2(new_n772), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n970), .B2(new_n830), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n790), .A2(G311), .B1(new_n858), .B2(G303), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n819), .B2(new_n791), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G317), .B2(new_n798), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT108), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT48), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1062), .B(KEYINPUT108), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n816), .A2(G283), .B1(new_n1025), .B2(G294), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n592), .B1(new_n488), .B2(new_n806), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n821), .B2(G326), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n821), .A2(G150), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n812), .A2(new_n333), .B1(new_n330), .B2(new_n787), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n791), .A2(new_n398), .B1(new_n795), .B2(new_n224), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n807), .A2(G97), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n797), .A2(new_n201), .B1(new_n785), .B2(new_n203), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n592), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1085), .A2(KEYINPUT109), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1047), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(KEYINPUT109), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1059), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1050), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1011), .A2(new_n756), .A3(new_n1012), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1017), .A2(new_n1091), .A3(new_n717), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1090), .A2(new_n1092), .ZN(G393));
  INV_X1    g0893(.A(KEYINPUT110), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n710), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n709), .A2(KEYINPUT110), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n996), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n710), .A2(new_n1000), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1020), .B(new_n717), .C1(new_n1013), .C2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(KEYINPUT111), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n761), .B1(new_n1099), .B2(KEYINPUT111), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n968), .A2(new_n770), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n772), .B1(new_n370), .B2(new_n215), .C1(new_n774), .C2(new_n243), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(KEYINPUT112), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n763), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n797), .A2(new_n818), .B1(new_n791), .B2(new_n1028), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT52), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n821), .A2(G322), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n324), .B1(new_n785), .B2(new_n849), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G116), .B2(new_n816), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n790), .A2(G303), .B1(new_n1025), .B2(G283), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1110), .A2(new_n808), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n795), .A2(new_n203), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n787), .A2(new_n224), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G50), .C2(new_n790), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n592), .B1(new_n261), .B2(new_n858), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n862), .C2(new_n803), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1040), .A2(G159), .B1(new_n792), .B2(G150), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n855), .A3(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1109), .A2(new_n1114), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1107), .B1(new_n771), .B2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1101), .A2(new_n1102), .B1(new_n1103), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1100), .A2(new_n1127), .ZN(G390));
  AOI21_X1  g0928(.A(new_n929), .B1(new_n836), .B2(new_n927), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n935), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n890), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n919), .A2(new_n925), .A3(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n706), .B(new_n927), .C1(new_n731), .C2(new_n733), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n930), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n935), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n890), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n923), .B2(new_n915), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n754), .A2(new_n935), .A3(G330), .A4(new_n927), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n946), .A2(new_n947), .A3(G330), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n935), .B1(new_n841), .B2(new_n927), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1141), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n931), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n946), .A2(G330), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT114), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n839), .B1(new_n1147), .B2(KEYINPUT114), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n935), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1133), .A2(new_n1139), .A3(new_n930), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n469), .A2(G330), .A3(new_n946), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n657), .B(new_n1153), .C1(new_n940), .C2(new_n735), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1143), .A2(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n717), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n919), .A2(new_n768), .A3(new_n925), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n763), .B1(new_n261), .B2(new_n847), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n868), .B1(G87), .B2(new_n824), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n791), .A2(new_n852), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n1116), .C1(new_n318), .C2(new_n790), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n324), .B1(new_n785), .B2(new_n370), .C1(new_n488), .C2(new_n797), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n821), .B2(G294), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1162), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n812), .A2(new_n1043), .B1(new_n785), .B2(new_n1168), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(KEYINPUT115), .B1(G159), .B2(new_n816), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(KEYINPUT115), .B2(new_n1169), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT116), .Z(new_n1172));
  OAI21_X1  g0972(.A(new_n293), .B1(new_n806), .B2(new_n201), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n821), .B2(G125), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT117), .ZN(new_n1175));
  INV_X1    g0975(.A(G132), .ZN(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n797), .A2(new_n1176), .B1(new_n791), .B2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT118), .Z(new_n1179));
  NOR2_X1   g0979(.A1(new_n795), .A2(new_n860), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1167), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1161), .B1(new_n1183), .B2(new_n771), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1143), .A2(new_n762), .B1(new_n1160), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1159), .A2(new_n1185), .ZN(G378));
  NAND2_X1  g0986(.A1(new_n919), .A2(new_n925), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1136), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n936), .A2(new_n937), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n949), .A2(new_n950), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n956), .B1(new_n951), .B2(new_n948), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n307), .A2(new_n308), .A3(new_n313), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n275), .A2(new_n897), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n307), .A2(new_n308), .A3(new_n313), .A4(new_n1194), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1191), .A2(new_n1192), .A3(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1190), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1203), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1191), .A2(new_n1192), .A3(new_n1203), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n939), .A3(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1206), .A2(new_n1211), .A3(KEYINPUT121), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT121), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n761), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n764), .B1(new_n201), .B2(new_n846), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n812), .A2(new_n1176), .B1(new_n795), .B2(new_n1168), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1040), .A2(G128), .B1(new_n858), .B2(G137), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n860), .B2(new_n787), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(G125), .C2(new_n792), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT59), .Z(new_n1220));
  OR2_X1    g1020(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(KEYINPUT119), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT120), .B(G124), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n821), .A2(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G33), .B(G41), .C1(new_n1033), .C2(G159), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1221), .A2(new_n1222), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n821), .A2(G283), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n462), .A2(G41), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1040), .A2(G107), .B1(new_n858), .B2(new_n329), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(new_n1037), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n791), .A2(new_n488), .B1(new_n795), .B2(new_n224), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n812), .A2(new_n370), .B1(new_n202), .B2(new_n806), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1228), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1236), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n1226), .A2(new_n1234), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1215), .B1(new_n1047), .B2(new_n1238), .C1(new_n1203), .C2(new_n769), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT122), .B1(new_n1214), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1206), .A2(new_n1211), .A3(KEYINPUT121), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n762), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT122), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1239), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1154), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1249), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n717), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1251), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1249), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1241), .A2(new_n1248), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G375));
  OAI211_X1 g1058(.A(new_n1154), .B(new_n1146), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  OR3_X1    g1060(.A1(new_n1156), .A2(new_n1260), .A3(new_n988), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1130), .A2(new_n768), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n763), .B1(G68), .B2(new_n847), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n803), .A2(new_n1029), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n324), .B1(new_n797), .B2(new_n852), .C1(new_n319), .C2(new_n785), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n329), .A2(new_n816), .B1(new_n792), .B2(G294), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(new_n488), .C2(new_n812), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n867), .A2(new_n224), .B1(new_n370), .B2(new_n870), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n592), .B1(G150), .B2(new_n858), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1270), .B1(new_n1177), .B2(new_n803), .C1(new_n861), .C2(new_n1043), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1168), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n790), .A2(new_n1272), .B1(new_n1033), .B2(G58), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G50), .A2(new_n816), .B1(new_n792), .B2(G132), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n870), .C2(new_n398), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1268), .A2(new_n1269), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1263), .B1(new_n1276), .B2(new_n771), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1152), .A2(new_n762), .B1(new_n1262), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1261), .A2(new_n1278), .ZN(G381));
  NAND3_X1  g1079(.A1(new_n834), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1280), .A2(G384), .ZN(new_n1281));
  NOR4_X1   g1081(.A1(G378), .A2(G390), .A3(G381), .A4(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1257), .A2(new_n1282), .A3(new_n1022), .A4(new_n1048), .ZN(G407));
  INV_X1    g1083(.A(G378), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n690), .A2(G213), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(KEYINPUT123), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1257), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(G407), .A2(G213), .A3(new_n1287), .ZN(G409));
  NOR3_X1   g1088(.A1(new_n1212), .A2(new_n1213), .A3(new_n1251), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1256), .B1(new_n1289), .B2(KEYINPUT57), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1246), .A2(new_n1247), .A3(new_n1239), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1247), .B1(new_n1246), .B2(new_n1239), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1290), .B(G378), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n988), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1242), .A2(KEYINPUT124), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n761), .B1(new_n1242), .B2(KEYINPUT124), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1240), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1284), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1286), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT60), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(new_n1259), .C1(new_n1156), .C2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT125), .B1(new_n1306), .B2(new_n1260), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1253), .B1(new_n1260), .B2(KEYINPUT60), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1278), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n875), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(G384), .A3(new_n1278), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1301), .A2(new_n1302), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1286), .A2(G2897), .ZN(new_n1317));
  OR3_X1    g1117(.A1(new_n1313), .A2(KEYINPUT126), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT126), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1311), .A2(new_n1319), .A3(new_n1312), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1321), .B2(new_n1317), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1257), .B2(G378), .ZN(new_n1324));
  OAI211_X1 g1124(.A(new_n1318), .B(new_n1322), .C1(new_n1324), .C2(new_n1286), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1301), .A2(new_n1327), .A3(new_n1302), .A4(new_n1314), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1316), .A2(new_n1325), .A3(new_n1326), .A4(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1022), .A2(new_n1048), .A3(G390), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G390), .B1(new_n1022), .B2(new_n1048), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G393), .A2(G396), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1280), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(KEYINPUT127), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1331), .A2(new_n1332), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1334), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(G390), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(G387), .A2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1339), .B1(new_n1341), .B2(new_n1330), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1336), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1329), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT63), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1343), .B1(new_n1345), .B2(new_n1315), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1302), .A4(new_n1314), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1346), .A2(new_n1326), .A3(new_n1325), .A4(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1344), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(G375), .A2(new_n1284), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1313), .A3(new_n1293), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1257), .A2(G378), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1293), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1314), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1351), .A2(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1355), .B(new_n1343), .ZN(G402));
endmodule


