//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n202), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n207), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(G20), .B2(new_n203), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n252), .A2(new_n251), .ZN(new_n263));
  OAI221_X1 g0063(.A(new_n250), .B1(new_n253), .B2(new_n255), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  INV_X1    g0065(.A(G274), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n213), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n213), .A2(new_n267), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n269), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n278), .B2(new_n279), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n282), .B1(new_n224), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n251), .B1(G33), .B2(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n275), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G190), .ZN(new_n289));
  INV_X1    g0089(.A(G200), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n265), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n264), .B1(new_n288), .B2(G169), .ZN(new_n294));
  INV_X1    g0094(.A(G179), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n288), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n252), .A2(new_n251), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n260), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n257), .A2(new_n224), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT11), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(KEYINPUT68), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT12), .B1(new_n248), .B2(G68), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n248), .A2(KEYINPUT12), .A3(G68), .ZN(new_n308));
  INV_X1    g0108(.A(new_n253), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n218), .B1(new_n206), .B2(G20), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n307), .A2(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n306), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n271), .B1(new_n219), .B2(new_n274), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n233), .A2(G1698), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n280), .B(new_n316), .C1(G226), .C2(G1698), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G97), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n314), .B(new_n315), .C1(new_n319), .C2(new_n273), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n273), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT13), .B1(new_n321), .B2(new_n313), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(G169), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(G179), .A3(new_n322), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n323), .B2(G169), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n312), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n306), .A2(new_n311), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n320), .A2(G190), .A3(new_n322), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n323), .A2(G200), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n330), .A2(new_n305), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n309), .A2(G77), .A3(new_n254), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT66), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G58), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT8), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT8), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G58), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(KEYINPUT15), .B(G87), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n257), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n300), .B1(new_n224), .B2(new_n249), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n337), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT67), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n350), .B1(new_n226), .B2(new_n280), .C1(new_n284), .C2(new_n219), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n287), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n274), .A2(new_n225), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n287), .A2(new_n266), .A3(new_n269), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT65), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT65), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n348), .A2(new_n349), .B1(G200), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n357), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G190), .B1(new_n347), .B2(KEYINPUT67), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n295), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n347), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n299), .A2(new_n334), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n287), .A2(new_n270), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(G232), .B1(new_n270), .B2(new_n268), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n285), .A2(new_n281), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n272), .A2(G1698), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n370), .B(new_n371), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n287), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n290), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n271), .B1(new_n233), .B2(new_n274), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n273), .B1(new_n374), .B2(new_n375), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  XOR2_X1   g0184(.A(KEYINPUT69), .B(KEYINPUT7), .Z(new_n385));
  NAND3_X1  g0185(.A1(new_n278), .A2(new_n207), .A3(new_n279), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n279), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n218), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n338), .A2(new_n218), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n259), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n384), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n218), .B1(new_n386), .B2(KEYINPUT7), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n372), .A2(new_n373), .A3(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n385), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(G58), .B(G68), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(G20), .B1(G159), .B2(new_n259), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(new_n300), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n342), .A2(new_n254), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n403), .A2(new_n253), .B1(new_n248), .B2(new_n342), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT70), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n383), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT17), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n393), .B1(new_n397), .B2(new_n395), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n263), .B1(new_n409), .B2(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(KEYINPUT70), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n404), .A2(KEYINPUT70), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n410), .A2(new_n394), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n383), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n408), .A2(new_n414), .A3(KEYINPUT72), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT72), .B1(new_n408), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n401), .A2(new_n300), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n388), .B1(new_n396), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G68), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT16), .B1(new_n421), .B2(new_n400), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n405), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT71), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT71), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n402), .A2(new_n425), .A3(new_n405), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n369), .A2(new_n377), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G169), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(new_n295), .B2(new_n427), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n424), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT18), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n424), .A2(KEYINPUT18), .A3(new_n426), .A4(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n417), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n367), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT80), .B(G294), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G33), .ZN(new_n439));
  OAI211_X1 g0239(.A(G257), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n440));
  OAI211_X1 g0240(.A(G250), .B(new_n281), .C1(new_n372), .C2(new_n373), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n273), .B1(new_n442), .B2(KEYINPUT81), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n439), .A2(new_n440), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  INV_X1    g0246(.A(G41), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n206), .A2(G45), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n451), .B1(new_n452), .B2(G41), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(G41), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT74), .A3(new_n206), .A4(G45), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n458), .A2(new_n273), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n443), .A2(new_n445), .B1(new_n459), .B2(G264), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n450), .A2(new_n455), .A3(new_n457), .A4(new_n268), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n363), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(G264), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n287), .A3(new_n445), .ZN(new_n465));
  AND4_X1   g0265(.A1(G179), .A2(new_n463), .A3(new_n465), .A4(new_n461), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT82), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n463), .A2(new_n465), .A3(new_n461), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G169), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n460), .A2(G179), .A3(new_n461), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n280), .A2(new_n207), .A3(G87), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT24), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G20), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n207), .B2(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n226), .A2(KEYINPUT23), .A3(G20), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n474), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n300), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT25), .B1(new_n249), .B2(new_n226), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n206), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n263), .A2(new_n248), .A3(new_n487), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n485), .A2(new_n486), .B1(new_n488), .B2(new_n226), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n467), .A2(new_n472), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n467), .A2(new_n472), .A3(new_n491), .A4(KEYINPUT83), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n290), .B1(new_n460), .B2(new_n461), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n468), .A2(new_n381), .ZN(new_n497));
  OR3_X1    g0297(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n344), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n248), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n488), .A2(new_n220), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n207), .B(G68), .C1(new_n372), .C2(new_n373), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n257), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n207), .B1(new_n318), .B2(new_n504), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n220), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n507), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n503), .B(new_n506), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n501), .B(new_n502), .C1(new_n513), .C2(new_n300), .ZN(new_n514));
  OAI211_X1 g0314(.A(G244), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n515));
  OAI211_X1 g0315(.A(G238), .B(new_n281), .C1(new_n372), .C2(new_n373), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(new_n476), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT77), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT77), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .A4(new_n476), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n287), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n287), .B1(new_n221), .B2(new_n449), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n206), .A2(new_n266), .A3(G45), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(G190), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n273), .B1(new_n517), .B2(KEYINPUT77), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n520), .B1(new_n523), .B2(new_n522), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n514), .B(new_n525), .C1(new_n290), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n513), .A2(new_n300), .ZN(new_n529));
  INV_X1    g0329(.A(new_n501), .ZN(new_n530));
  INV_X1    g0330(.A(new_n488), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n500), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n521), .A2(new_n295), .A3(new_n524), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n533), .B(new_n534), .C1(G169), .C2(new_n527), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n248), .A2(G97), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n488), .B2(new_n505), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n420), .A2(G107), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n509), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n226), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n539), .B1(new_n547), .B2(new_n300), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n458), .A2(G257), .A3(new_n273), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n461), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n283), .B2(G250), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(new_n281), .C1(new_n372), .C2(new_n373), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT73), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n372), .A2(new_n373), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n281), .A2(KEYINPUT4), .A3(G244), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n559), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n280), .A2(new_n561), .A3(KEYINPUT73), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n553), .A2(new_n556), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n550), .B1(new_n287), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n548), .B1(new_n564), .B2(new_n295), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT76), .ZN(new_n566));
  INV_X1    g0366(.A(new_n550), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n287), .ZN(new_n568));
  AOI21_X1  g0368(.A(G169), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n295), .A3(new_n461), .A4(new_n549), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n545), .A2(G20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n259), .A2(G77), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n226), .B1(new_n387), .B2(new_n388), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n300), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n539), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n572), .B(new_n579), .C1(new_n564), .C2(G169), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n567), .A2(new_n568), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n583), .B(new_n548), .C1(new_n381), .C2(new_n582), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n536), .A2(new_n571), .A3(new_n581), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n458), .A2(new_n273), .ZN(new_n587));
  INV_X1    g0387(.A(G270), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n280), .A2(G257), .A3(new_n281), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n558), .A2(G303), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n284), .C2(new_n227), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n287), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n458), .A2(KEYINPUT79), .A3(G270), .A4(new_n273), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n589), .A2(new_n461), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n551), .B(new_n207), .C1(G33), .C2(new_n505), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n300), .C1(new_n207), .C2(G116), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT20), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n248), .A2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n531), .B2(G116), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n363), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT21), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n595), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n599), .A2(new_n601), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n595), .B2(G200), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n381), .B2(new_n595), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n589), .A2(new_n461), .A3(new_n594), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n295), .B1(new_n592), .B2(new_n287), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n607), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n585), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n437), .A2(new_n499), .A3(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n437), .ZN(new_n617));
  INV_X1    g0417(.A(new_n535), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n571), .A2(new_n581), .ZN(new_n619));
  XNOR2_X1  g0419(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n536), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT26), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n528), .A2(new_n535), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(new_n580), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n618), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n571), .A2(new_n581), .A3(new_n584), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n469), .A2(new_n470), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n491), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n607), .A3(new_n613), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n627), .A2(new_n630), .A3(new_n498), .A4(new_n536), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n617), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT72), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n406), .A2(new_n407), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT17), .B1(new_n413), .B2(new_n383), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n408), .A2(new_n414), .A3(KEYINPUT72), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n365), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n333), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n329), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT85), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n379), .A2(new_n380), .A3(new_n295), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n427), .B2(G169), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n413), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT85), .B1(new_n423), .B2(new_n429), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n431), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n643), .B1(new_n413), .B2(new_n645), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n423), .A2(new_n429), .A3(KEYINPUT85), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(KEYINPUT18), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n297), .B1(new_n653), .B2(new_n293), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n633), .A2(new_n654), .ZN(G369));
  AND2_X1   g0455(.A1(new_n607), .A2(new_n613), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT86), .Z(new_n659));
  INV_X1    g0459(.A(G213), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n657), .B2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G343), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n608), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n656), .A2(new_n610), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n656), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  INV_X1    g0469(.A(new_n499), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n491), .A2(new_n665), .ZN(new_n671));
  XOR2_X1   g0471(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n492), .A2(new_n664), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n656), .A2(new_n665), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n491), .A2(new_n628), .A3(new_n664), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n675), .A2(new_n679), .ZN(G399));
  NAND2_X1  g0480(.A1(new_n210), .A2(new_n447), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n510), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n216), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n632), .A2(new_n664), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(KEYINPUT29), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n624), .A2(new_n623), .A3(new_n580), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n566), .B1(new_n565), .B2(new_n570), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n572), .A2(new_n579), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n690), .A2(KEYINPUT76), .A3(new_n569), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n536), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n688), .B1(new_n692), .B2(new_n620), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT89), .B1(new_n693), .B2(new_n618), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n494), .A2(new_n495), .A3(new_n656), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n585), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT89), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n621), .B1(new_n619), .B2(new_n536), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n699), .B(new_n535), .C1(new_n700), .C2(new_n688), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n664), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n687), .B1(KEYINPUT29), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n494), .A2(new_n495), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n585), .A2(new_n614), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n706), .A2(new_n498), .A3(new_n707), .A4(new_n664), .ZN(new_n708));
  AOI21_X1  g0508(.A(G179), .B1(new_n521), .B2(new_n524), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT88), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n595), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n595), .B2(new_n709), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n468), .B(new_n582), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n463), .A2(new_n465), .A3(new_n524), .A4(new_n521), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n611), .A3(new_n612), .A4(new_n564), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n564), .A2(new_n612), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n714), .A3(KEYINPUT30), .A4(new_n611), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n713), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT31), .B1(new_n720), .B2(new_n665), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n705), .B1(new_n708), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n704), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n685), .B1(new_n727), .B2(G1), .ZN(G364));
  INV_X1    g0528(.A(new_n681), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n207), .A2(G13), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n206), .B1(new_n730), .B2(G45), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n210), .A2(new_n280), .ZN(new_n734));
  INV_X1    g0534(.A(G355), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(G116), .B2(new_n210), .ZN(new_n736));
  INV_X1    g0536(.A(G45), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n243), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n210), .A2(new_n558), .ZN(new_n739));
  INV_X1    g0539(.A(new_n216), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n736), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n251), .B1(G20), .B2(new_n363), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n733), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n505), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n558), .ZN(new_n756));
  NAND2_X1  g0556(.A1(G20), .A2(G179), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT90), .Z(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n381), .A3(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n295), .A2(G200), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT95), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n207), .B1(new_n760), .B2(KEYINPUT95), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(G190), .A3(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n756), .B1(new_n218), .B2(new_n759), .C1(new_n220), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n207), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n751), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT94), .B(G159), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(KEYINPUT32), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT32), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G190), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  OR3_X1    g0574(.A1(new_n764), .A2(new_n769), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n758), .A2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n290), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n202), .A2(new_n778), .B1(new_n780), .B2(new_n338), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n758), .A2(new_n381), .A3(new_n290), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT91), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT91), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n786), .B2(G77), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT92), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n558), .B1(new_n763), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT97), .Z(new_n791));
  INV_X1    g0591(.A(new_n438), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT33), .B(G317), .Z(new_n793));
  OAI22_X1  g0593(.A1(new_n754), .A2(new_n792), .B1(new_n759), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT96), .B(G326), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n778), .A2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(G322), .C2(new_n779), .ZN(new_n797));
  INV_X1    g0597(.A(new_n766), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G329), .B1(new_n772), .B2(G283), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n797), .B(new_n799), .C1(new_n800), .C2(new_n785), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n775), .A2(new_n788), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n749), .B1(new_n802), .B2(new_n746), .ZN(new_n803));
  INV_X1    g0603(.A(new_n745), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n668), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n733), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n669), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n668), .A2(G330), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n640), .A2(new_n664), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n358), .A2(new_n360), .B1(new_n347), .B2(new_n665), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n640), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n686), .B(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n733), .B1(new_n813), .B2(new_n725), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n725), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n746), .A2(new_n743), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n806), .B1(new_n224), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n365), .A2(new_n665), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n361), .B1(new_n348), .B2(new_n664), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n365), .ZN(new_n820));
  INV_X1    g0620(.A(new_n746), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G137), .A2(new_n777), .B1(new_n779), .B2(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n258), .B2(new_n759), .C1(new_n785), .C2(new_n767), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(new_n772), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n218), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n280), .B1(new_n827), .B2(new_n766), .C1(new_n754), .C2(new_n338), .ZN(new_n828));
  INV_X1    g0628(.A(new_n763), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n828), .C1(G50), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n825), .A2(new_n220), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n780), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(G303), .C2(new_n777), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n280), .B(new_n755), .C1(G311), .C2(new_n798), .ZN(new_n835));
  INV_X1    g0635(.A(new_n759), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(G283), .B1(new_n829), .B2(G107), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n786), .A2(G116), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n824), .A2(new_n830), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n817), .B1(new_n820), .B2(new_n744), .C1(new_n821), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n815), .A2(new_n841), .ZN(G384));
  AND2_X1   g0642(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n545), .A2(KEYINPUT35), .ZN(new_n844));
  INV_X1    g0644(.A(G116), .ZN(new_n845));
  NOR4_X1   g0645(.A1(new_n843), .A2(new_n844), .A3(new_n215), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT36), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n390), .A2(new_n216), .A3(new_n224), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT98), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n848), .A2(KEYINPUT98), .B1(new_n202), .B2(G68), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n206), .B(G13), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n404), .B1(new_n855), .B2(new_n410), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n856), .A2(new_n662), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n417), .B2(new_n434), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n424), .A2(new_n426), .A3(new_n663), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n413), .B2(new_n383), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n430), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n406), .B1(new_n856), .B2(new_n645), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n863), .B2(new_n857), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n854), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n432), .A2(new_n433), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n857), .B1(new_n868), .B2(new_n639), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n312), .A2(new_n665), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT100), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n334), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n872), .A2(new_n327), .A3(new_n328), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n334), .B2(KEYINPUT100), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n874), .A2(new_n876), .A3(new_n820), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n615), .A2(new_n499), .A3(new_n665), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n720), .A2(new_n665), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT31), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n853), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n635), .A2(new_n636), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n648), .A2(new_n886), .A3(new_n651), .ZN(new_n887));
  INV_X1    g0687(.A(new_n860), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n413), .B2(new_n383), .ZN(new_n891));
  AND4_X1   g0691(.A1(new_n890), .A2(new_n383), .A3(new_n402), .A4(new_n405), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n893), .A2(new_n649), .A3(new_n650), .A4(new_n860), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n430), .A2(new_n861), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n894), .A2(KEYINPUT37), .B1(new_n895), .B2(new_n860), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n854), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT103), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n870), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n874), .A2(new_n876), .A3(new_n820), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n708), .B2(new_n723), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n869), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n865), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(KEYINPUT40), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n885), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT104), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n878), .A2(new_n883), .ZN(new_n906));
  OR3_X1    g0706(.A1(new_n905), .A2(new_n437), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n437), .B2(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(G330), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n652), .A2(new_n662), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n874), .A2(new_n876), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n665), .B(new_n812), .C1(new_n626), .C2(new_n631), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n810), .B(KEYINPUT99), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n915), .B2(new_n871), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT101), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT39), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n899), .A2(new_n919), .A3(new_n902), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n329), .A2(new_n665), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(KEYINPUT101), .B(new_n910), .C1(new_n915), .C2(new_n871), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n654), .B1(new_n704), .B2(new_n437), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n909), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n206), .B2(new_n730), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n909), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n852), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NOR2_X1   g0732(.A1(new_n664), .A2(new_n514), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n618), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n624), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n936));
  INV_X1    g0736(.A(new_n675), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n627), .B1(new_n548), .B2(new_n664), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n565), .A2(new_n665), .A3(new_n570), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT105), .Z(new_n941));
  NOR2_X1   g0741(.A1(new_n937), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n936), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n937), .A2(new_n941), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT106), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n949), .C1(KEYINPUT43), .C2(new_n935), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n941), .A2(new_n706), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n664), .B1(new_n952), .B2(new_n619), .ZN(new_n953));
  INV_X1    g0753(.A(new_n940), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n677), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n955), .A2(KEYINPUT42), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n957), .A2(new_n958), .B1(KEYINPUT43), .B2(new_n935), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n951), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n681), .B(KEYINPUT41), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n679), .A2(KEYINPUT44), .A3(new_n954), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT44), .B1(new_n679), .B2(new_n954), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n679), .A2(KEYINPUT107), .A3(new_n954), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT107), .B1(new_n679), .B2(new_n954), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT45), .B1(new_n965), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n675), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n673), .B(new_n674), .C1(new_n656), .C2(new_n665), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n971), .A2(new_n677), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n669), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n669), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n726), .ZN(new_n976));
  INV_X1    g0776(.A(new_n969), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n977), .A2(new_n937), .A3(new_n964), .A4(new_n967), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n961), .B1(new_n979), .B2(new_n727), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n960), .B1(new_n980), .B2(new_n732), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n747), .B1(new_n210), .B2(new_n344), .C1(new_n239), .C2(new_n739), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n982), .A2(new_n733), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n778), .A2(new_n800), .B1(new_n792), .B2(new_n759), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n780), .A2(new_n789), .B1(new_n754), .B2(new_n226), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(G283), .C2(new_n786), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n825), .A2(new_n505), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n829), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT46), .B1(new_n829), .B2(G116), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n558), .B1(new_n766), .B2(new_n990), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n786), .A2(G50), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n753), .A2(G68), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n767), .B2(new_n759), .C1(new_n224), .C2(new_n825), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n777), .A2(G143), .ZN(new_n996));
  INV_X1    g0796(.A(G137), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n280), .C1(new_n997), .C2(new_n766), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n780), .A2(new_n258), .B1(new_n763), .B2(new_n338), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n995), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n986), .A2(new_n992), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n983), .B1(new_n804), .B2(new_n935), .C1(new_n1002), .C2(new_n821), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n981), .A2(new_n1003), .ZN(G387));
  INV_X1    g0804(.A(new_n975), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n673), .A2(new_n674), .A3(new_n745), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n734), .A2(new_n682), .B1(G107), .B2(new_n210), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n236), .A2(new_n737), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n682), .ZN(new_n1009));
  AOI211_X1 g0809(.A(G45), .B(new_n1009), .C1(G68), .C2(G77), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n256), .A2(G50), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n739), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1007), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n733), .B1(new_n1014), .B2(new_n748), .ZN(new_n1015));
  INV_X1    g0815(.A(G159), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n202), .A2(new_n780), .B1(new_n778), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n342), .B2(new_n836), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n558), .B(new_n987), .C1(G150), .C2(new_n798), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n786), .A2(G68), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n753), .A2(new_n500), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n829), .A2(G77), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n795), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n280), .B1(new_n798), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n759), .A2(new_n800), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT108), .B(G322), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(new_n777), .B2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n990), .B2(new_n780), .C1(new_n785), .C2(new_n789), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n753), .A2(G283), .B1(new_n829), .B2(new_n438), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1026), .B1(new_n845), .B2(new_n825), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1024), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT109), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n821), .B1(new_n1039), .B2(KEYINPUT109), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1015), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1005), .A2(new_n732), .B1(new_n1006), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n729), .B1(new_n975), .B2(new_n726), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1005), .A2(new_n727), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(G393));
  NAND3_X1  g0846(.A1(new_n970), .A2(new_n978), .A3(new_n732), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n941), .A2(new_n745), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT110), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT51), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n258), .A2(new_n778), .B1(new_n780), .B2(new_n1016), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1050), .A2(new_n1051), .B1(new_n786), .B2(new_n342), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n558), .B(new_n831), .C1(G143), .C2(new_n798), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n836), .A2(G50), .B1(new_n753), .B2(G77), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n218), .C2(new_n763), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n836), .A2(G303), .B1(new_n753), .B2(G116), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT111), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n786), .A2(G294), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n798), .A2(new_n1028), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n773), .A3(new_n558), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G283), .B2(new_n829), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1059), .B(new_n1062), .C1(new_n1058), .C2(new_n1057), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n779), .B1(new_n777), .B2(G317), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT52), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1053), .A2(new_n1056), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n746), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n747), .B1(new_n505), .B2(new_n210), .C1(new_n246), .C2(new_n739), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1049), .A2(new_n733), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n979), .A2(new_n729), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n976), .B1(new_n970), .B2(new_n978), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1047), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(G390));
  NOR2_X1   g0872(.A1(new_n913), .A2(new_n914), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n724), .A2(new_n820), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n911), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n724), .A2(new_n820), .A3(new_n912), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n819), .A2(new_n365), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n702), .A2(new_n664), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n810), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT112), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(KEYINPUT112), .A3(new_n810), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n725), .A2(new_n437), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1088), .B(new_n654), .C1(new_n437), .C2(new_n704), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1076), .A2(KEYINPUT113), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1082), .A2(new_n912), .A3(new_n1083), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n899), .A2(new_n902), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n921), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n920), .A2(new_n923), .B1(new_n915), .B2(new_n921), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1092), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1091), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1079), .A2(KEYINPUT112), .A3(new_n810), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT112), .B1(new_n1079), .B2(new_n810), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n911), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1099), .B1(new_n1105), .B2(new_n1095), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1091), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n927), .A2(new_n1087), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n1077), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1097), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1107), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1102), .A2(new_n1113), .A3(new_n729), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n754), .A2(new_n1016), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n558), .B(new_n1115), .C1(G125), .C2(new_n798), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  INV_X1    g0917(.A(KEYINPUT53), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n763), .B2(new_n258), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n829), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n786), .A2(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G128), .A2(new_n777), .B1(new_n836), .B2(G137), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n779), .A2(G132), .B1(new_n772), .B2(G50), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT114), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n558), .B1(new_n763), .B2(new_n220), .C1(new_n832), .C2(new_n766), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1126), .B(new_n826), .C1(G77), .C2(new_n753), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n780), .A2(new_n845), .B1(new_n226), .B2(new_n759), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G283), .B2(new_n777), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1127), .B(new_n1129), .C1(new_n505), .C2(new_n785), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT115), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n746), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n816), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n733), .C1(new_n342), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n920), .A2(new_n923), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n743), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT116), .Z(new_n1137));
  NAND2_X1  g0937(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n732), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n1139), .ZN(G378));
  NAND3_X1  g0940(.A1(new_n885), .A2(new_n903), .A3(G330), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n264), .A2(new_n663), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n293), .A2(new_n298), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n293), .B2(new_n298), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OR3_X1    g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1141), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n885), .A2(new_n903), .A3(new_n1149), .A4(G330), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n926), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n925), .A2(new_n924), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1155), .A2(new_n1151), .A3(new_n918), .A4(new_n1152), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n731), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1150), .A2(new_n743), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n733), .B1(G50), .B2(new_n1133), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n829), .A2(new_n1117), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1160), .B1(new_n827), .B2(new_n759), .C1(new_n780), .C2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n777), .A2(G125), .B1(new_n753), .B2(G150), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT118), .Z(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G137), .C2(new_n786), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT59), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(G33), .A2(G41), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT117), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n825), .A2(new_n767), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(G124), .C2(new_n798), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n1168), .A3(new_n1172), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n226), .A2(new_n780), .B1(new_n778), .B2(new_n845), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G97), .B2(new_n836), .ZN(new_n1175));
  AOI211_X1 g0975(.A(G41), .B(new_n280), .C1(new_n798), .C2(G283), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n772), .A2(G58), .ZN(new_n1177));
  AND4_X1   g0977(.A1(new_n994), .A2(new_n1176), .A3(new_n1022), .A4(new_n1177), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(new_n344), .C2(new_n785), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT58), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1170), .B(new_n202), .C1(G41), .C2(new_n280), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1173), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1159), .B1(new_n1184), .B2(new_n746), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1158), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1157), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT57), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1111), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n1089), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n729), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1188), .B1(new_n1193), .B2(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n961), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1111), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n777), .A2(G294), .B1(new_n829), .B2(G97), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n845), .B2(new_n759), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n779), .A2(G283), .B1(new_n753), .B2(new_n500), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n280), .B1(new_n798), .B2(G303), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n224), .C2(new_n825), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1203), .B(new_n1206), .C1(G107), .C2(new_n786), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n785), .A2(new_n258), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n836), .A2(new_n1117), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n1016), .B2(new_n763), .C1(new_n754), .C2(new_n202), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n827), .A2(new_n778), .B1(new_n780), .B2(new_n997), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1177), .B(new_n280), .C1(new_n1161), .C2(new_n766), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n746), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n806), .B1(new_n218), .B2(new_n816), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n912), .C2(new_n744), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1086), .B2(new_n731), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1201), .A2(new_n1218), .ZN(G381));
  INV_X1    g1019(.A(G378), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1221));
  INV_X1    g1021(.A(G390), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1223), .A2(G387), .A3(G375), .ZN(G407));
  NOR2_X1   g1024(.A1(new_n660), .A2(G343), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1220), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(G375), .C2(new_n1226), .ZN(G409));
  AOI21_X1  g1027(.A(G390), .B1(new_n981), .B2(new_n1003), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT122), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n981), .A2(new_n1003), .A3(G390), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(KEYINPUT123), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n981), .A2(G390), .A3(new_n1232), .A4(new_n1003), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1229), .A2(new_n1231), .A3(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(G393), .B(G396), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1228), .B2(KEYINPUT122), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1230), .A2(KEYINPUT121), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1222), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G387), .A2(KEYINPUT121), .A3(new_n1222), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G378), .B(new_n1188), .C1(new_n1193), .C2(new_n1197), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1194), .A2(new_n1200), .A3(new_n1196), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT119), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(new_n1186), .C1(new_n1195), .C2(new_n731), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT119), .B1(new_n1157), .B2(new_n1187), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1220), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1225), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1086), .A2(KEYINPUT60), .A3(new_n1089), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1253), .A2(new_n729), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT60), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1199), .B1(new_n1090), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1217), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  XOR2_X1   g1057(.A(G384), .B(KEYINPUT120), .Z(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G384), .A2(KEYINPUT120), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1217), .B(new_n1260), .C1(new_n1254), .C2(new_n1256), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G2897), .B(new_n1225), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1260), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1257), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1225), .A2(G2897), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1262), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1244), .B1(new_n1252), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT124), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(KEYINPUT124), .B(new_n1244), .C1(new_n1252), .C2(new_n1267), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1225), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1272), .B(new_n1273), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1270), .A2(new_n1271), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1252), .A2(KEYINPUT62), .A3(new_n1277), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT62), .B1(new_n1252), .B2(new_n1277), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1243), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1286), .A2(KEYINPUT63), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1288), .A2(new_n1235), .B1(new_n1236), .B2(new_n1234), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1268), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(KEYINPUT63), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1290), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1292), .ZN(G405));
  AOI21_X1  g1093(.A(new_n1195), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1192), .B(new_n729), .C1(new_n1294), .C2(KEYINPUT57), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1295), .A2(G378), .A3(new_n1188), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G378), .B1(new_n1295), .B2(new_n1188), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1278), .B1(new_n1298), .B2(KEYINPUT126), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G375), .A2(new_n1220), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1245), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  AOI211_X1 g1104(.A(KEYINPUT126), .B(KEYINPUT127), .C1(new_n1301), .C2(new_n1245), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1277), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1303), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT127), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1302), .A2(new_n1303), .A3(new_n1300), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1306), .A2(new_n1243), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1243), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


