

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X2 U323 ( .A(n476), .B(n475), .ZN(n534) );
  XNOR2_X1 U324 ( .A(n581), .B(KEYINPUT41), .ZN(n488) );
  XNOR2_X1 U325 ( .A(n404), .B(n403), .ZN(n421) );
  XNOR2_X1 U326 ( .A(G99GAT), .B(G85GAT), .ZN(n403) );
  NOR2_X2 U327 ( .A1(n539), .A2(n485), .ZN(n570) );
  XNOR2_X1 U328 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(n509) );
  XOR2_X1 U330 ( .A(KEYINPUT99), .B(n381), .Z(n291) );
  XOR2_X1 U331 ( .A(n341), .B(n340), .Z(n292) );
  XOR2_X1 U332 ( .A(G148GAT), .B(KEYINPUT75), .Z(n293) );
  XNOR2_X1 U333 ( .A(KEYINPUT108), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X1 U334 ( .A1(n529), .A2(n535), .ZN(n379) );
  NOR2_X1 U335 ( .A1(n563), .A2(n467), .ZN(n468) );
  XNOR2_X1 U336 ( .A(n429), .B(n293), .ZN(n430) );
  XNOR2_X1 U337 ( .A(n342), .B(n292), .ZN(n343) );
  XNOR2_X1 U338 ( .A(n478), .B(KEYINPUT54), .ZN(n479) );
  INV_X1 U339 ( .A(KEYINPUT28), .ZN(n346) );
  XNOR2_X1 U340 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n483) );
  XNOR2_X1 U341 ( .A(n346), .B(KEYINPUT65), .ZN(n347) );
  XNOR2_X1 U342 ( .A(n439), .B(n438), .ZN(n581) );
  XNOR2_X1 U343 ( .A(n482), .B(n347), .ZN(n537) );
  INV_X1 U344 ( .A(G43GAT), .ZN(n459) );
  XNOR2_X1 U345 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n486) );
  XNOR2_X1 U346 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U347 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(G78GAT), .B(G211GAT), .Z(n295) );
  XNOR2_X1 U350 ( .A(G127GAT), .B(G155GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n308) );
  XOR2_X1 U352 ( .A(G71GAT), .B(KEYINPUT13), .Z(n428) );
  XOR2_X1 U353 ( .A(KEYINPUT15), .B(n428), .Z(n297) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U356 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n299) );
  XNOR2_X1 U357 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U359 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G15GAT), .Z(n449) );
  XOR2_X1 U361 ( .A(G57GAT), .B(G183GAT), .Z(n303) );
  XNOR2_X1 U362 ( .A(G1GAT), .B(G8GAT), .ZN(n302) );
  XNOR2_X1 U363 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U364 ( .A(n449), .B(n304), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U366 ( .A(n308), .B(n307), .Z(n585) );
  XOR2_X1 U367 ( .A(G176GAT), .B(G120GAT), .Z(n310) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n327) );
  XOR2_X1 U370 ( .A(G71GAT), .B(G99GAT), .Z(n312) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(G15GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n313), .B(G134GAT), .Z(n315) );
  XOR2_X1 U374 ( .A(KEYINPUT0), .B(G127GAT), .Z(n357) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(n357), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U377 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n317) );
  NAND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U380 ( .A(n319), .B(n318), .Z(n325) );
  XNOR2_X1 U381 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n320), .B(KEYINPUT18), .ZN(n321) );
  XOR2_X1 U383 ( .A(n321), .B(KEYINPUT17), .Z(n323) );
  XNOR2_X1 U384 ( .A(G183GAT), .B(G190GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n375) );
  XNOR2_X1 U386 ( .A(n375), .B(KEYINPUT20), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U388 ( .A(n327), .B(n326), .Z(n539) );
  INV_X1 U389 ( .A(n539), .ZN(n527) );
  XOR2_X1 U390 ( .A(G148GAT), .B(KEYINPUT87), .Z(n329) );
  XNOR2_X1 U391 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U393 ( .A(n330), .B(KEYINPUT86), .Z(n332) );
  XNOR2_X1 U394 ( .A(G155GAT), .B(G162GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n365) );
  XOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .Z(n433) );
  XOR2_X1 U397 ( .A(G211GAT), .B(KEYINPUT21), .Z(n334) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n374) );
  XOR2_X1 U400 ( .A(n433), .B(n374), .Z(n336) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G22GAT), .ZN(n335) );
  XNOR2_X1 U402 ( .A(n336), .B(n335), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT23), .B(G204GAT), .Z(n338) );
  XNOR2_X1 U404 ( .A(G141GAT), .B(KEYINPUT24), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U406 ( .A(n339), .B(KEYINPUT22), .ZN(n342) );
  XOR2_X1 U407 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n341) );
  NAND2_X1 U408 ( .A1(G228GAT), .A2(G233GAT), .ZN(n340) );
  XOR2_X1 U409 ( .A(n365), .B(n345), .Z(n482) );
  INV_X1 U410 ( .A(n537), .ZN(n529) );
  XOR2_X1 U411 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n349) );
  XNOR2_X1 U412 ( .A(G29GAT), .B(G85GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n351) );
  XNOR2_X1 U415 ( .A(KEYINPUT1), .B(KEYINPUT90), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U417 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U418 ( .A(G134GAT), .B(KEYINPUT79), .Z(n395) );
  XOR2_X1 U419 ( .A(G120GAT), .B(G57GAT), .Z(n432) );
  XOR2_X1 U420 ( .A(n395), .B(n432), .Z(n355) );
  NAND2_X1 U421 ( .A1(G225GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U425 ( .A(n360), .B(KEYINPUT92), .Z(n363) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(G113GAT), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n361), .B(G1GAT), .ZN(n452) );
  XNOR2_X1 U428 ( .A(n452), .B(KEYINPUT91), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n388) );
  XNOR2_X1 U431 ( .A(KEYINPUT94), .B(n388), .ZN(n522) );
  XOR2_X1 U432 ( .A(G169GAT), .B(G8GAT), .Z(n451) );
  XOR2_X1 U433 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n367) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(G92GAT), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(n451), .B(n368), .Z(n370) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n373) );
  XOR2_X1 U439 ( .A(G64GAT), .B(KEYINPUT74), .Z(n372) );
  XNOR2_X1 U440 ( .A(G176GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U441 ( .A(n372), .B(n371), .ZN(n429) );
  XOR2_X1 U442 ( .A(n373), .B(n429), .Z(n377) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n477) );
  XNOR2_X1 U445 ( .A(n477), .B(KEYINPUT97), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n378), .B(KEYINPUT27), .ZN(n383) );
  NAND2_X1 U447 ( .A1(n522), .A2(n383), .ZN(n535) );
  XOR2_X1 U448 ( .A(KEYINPUT98), .B(n379), .Z(n380) );
  NOR2_X1 U449 ( .A1(n527), .A2(n380), .ZN(n381) );
  NOR2_X1 U450 ( .A1(n527), .A2(n482), .ZN(n382) );
  XNOR2_X1 U451 ( .A(n382), .B(KEYINPUT26), .ZN(n573) );
  NAND2_X1 U452 ( .A1(n573), .A2(n383), .ZN(n387) );
  INV_X1 U453 ( .A(n477), .ZN(n524) );
  NAND2_X1 U454 ( .A1(n527), .A2(n524), .ZN(n384) );
  NAND2_X1 U455 ( .A1(n482), .A2(n384), .ZN(n385) );
  XOR2_X1 U456 ( .A(KEYINPUT25), .B(n385), .Z(n386) );
  AND2_X1 U457 ( .A1(n387), .A2(n386), .ZN(n389) );
  NOR2_X1 U458 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U459 ( .A(KEYINPUT100), .B(n390), .ZN(n391) );
  NOR2_X1 U460 ( .A1(n291), .A2(n391), .ZN(n495) );
  NOR2_X1 U461 ( .A1(n585), .A2(n495), .ZN(n417) );
  XOR2_X1 U462 ( .A(KEYINPUT80), .B(G106GAT), .Z(n393) );
  XNOR2_X1 U463 ( .A(G190GAT), .B(G218GAT), .ZN(n392) );
  XNOR2_X1 U464 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U465 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U468 ( .A(n398), .B(KEYINPUT11), .Z(n406) );
  INV_X1 U469 ( .A(KEYINPUT73), .ZN(n399) );
  NAND2_X1 U470 ( .A1(n399), .A2(G92GAT), .ZN(n402) );
  INV_X1 U471 ( .A(G92GAT), .ZN(n400) );
  NAND2_X1 U472 ( .A1(n400), .A2(KEYINPUT73), .ZN(n401) );
  NAND2_X1 U473 ( .A1(n402), .A2(n401), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n421), .B(KEYINPUT78), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n406), .B(n405), .ZN(n416) );
  XOR2_X1 U476 ( .A(G43GAT), .B(G29GAT), .Z(n408) );
  XNOR2_X1 U477 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U479 ( .A(n409), .B(KEYINPUT69), .Z(n411) );
  XNOR2_X1 U480 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n446) );
  XOR2_X1 U482 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n413) );
  XNOR2_X1 U483 ( .A(G162GAT), .B(KEYINPUT9), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U485 ( .A(n446), .B(n414), .Z(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n563) );
  XNOR2_X1 U487 ( .A(KEYINPUT36), .B(n563), .ZN(n587) );
  NAND2_X1 U488 ( .A1(n417), .A2(n587), .ZN(n418) );
  XOR2_X1 U489 ( .A(KEYINPUT37), .B(n418), .Z(n521) );
  INV_X1 U490 ( .A(KEYINPUT32), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n421), .B(n419), .ZN(n420) );
  NAND2_X1 U492 ( .A1(G230GAT), .A2(G233GAT), .ZN(n422) );
  NAND2_X1 U493 ( .A1(n420), .A2(n422), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n421), .B(KEYINPUT32), .ZN(n424) );
  INV_X1 U495 ( .A(n422), .ZN(n423) );
  NAND2_X1 U496 ( .A1(n424), .A2(n423), .ZN(n425) );
  NAND2_X1 U497 ( .A1(n426), .A2(n425), .ZN(n427) );
  XOR2_X1 U498 ( .A(n428), .B(n427), .Z(n431) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n435) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n437) );
  XNOR2_X1 U503 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n436) );
  XOR2_X1 U504 ( .A(n437), .B(n436), .Z(n438) );
  XOR2_X1 U505 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n441) );
  NAND2_X1 U506 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U508 ( .A(n442), .B(KEYINPUT30), .Z(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n444) );
  XNOR2_X1 U510 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U514 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U515 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n575) );
  XNOR2_X1 U517 ( .A(n575), .B(KEYINPUT71), .ZN(n567) );
  INV_X1 U518 ( .A(n567), .ZN(n455) );
  NOR2_X1 U519 ( .A1(n581), .A2(n455), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n456), .B(KEYINPUT77), .ZN(n497) );
  NOR2_X1 U521 ( .A1(n521), .A2(n497), .ZN(n458) );
  XNOR2_X1 U522 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n457) );
  NAND2_X1 U523 ( .A1(n509), .A2(n527), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n460) );
  NOR2_X1 U525 ( .A1(n575), .A2(n488), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n465), .A2(n585), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT109), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT47), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n470) );
  NAND2_X1 U531 ( .A1(n585), .A2(n587), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n567), .A2(n581), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n534), .A2(n477), .ZN(n480) );
  INV_X1 U538 ( .A(KEYINPUT120), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n522), .A2(n481), .ZN(n574) );
  NAND2_X1 U541 ( .A1(n574), .A2(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n563), .A2(n570), .ZN(n487) );
  INV_X1 U544 ( .A(n488), .ZN(n541) );
  NAND2_X1 U545 ( .A1(n570), .A2(n541), .ZN(n492) );
  XOR2_X1 U546 ( .A(G176GAT), .B(KEYINPUT123), .Z(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(G1349GAT) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n499) );
  INV_X1 U551 ( .A(n585), .ZN(n560) );
  NOR2_X1 U552 ( .A1(n563), .A2(n560), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT16), .B(n493), .Z(n494) );
  NOR2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT101), .B(n496), .ZN(n512) );
  NOR2_X1 U556 ( .A1(n497), .A2(n512), .ZN(n503) );
  NAND2_X1 U557 ( .A1(n522), .A2(n503), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1324GAT) );
  NAND2_X1 U559 ( .A1(n524), .A2(n503), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U561 ( .A(G15GAT), .B(KEYINPUT35), .Z(n502) );
  NAND2_X1 U562 ( .A1(n503), .A2(n527), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1326GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n529), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U566 ( .A1(n509), .A2(n522), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1328GAT) );
  NAND2_X1 U570 ( .A1(n524), .A2(n509), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n529), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U574 ( .A1(n541), .A2(n575), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT105), .B(n511), .Z(n520) );
  NOR2_X1 U576 ( .A1(n512), .A2(n520), .ZN(n517) );
  NAND2_X1 U577 ( .A1(n522), .A2(n517), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n513), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n524), .A2(n517), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n527), .A2(n517), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U585 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n530) );
  NAND2_X1 U588 ( .A1(n522), .A2(n530), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n530), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(KEYINPUT106), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n530), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n532) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT112), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n553), .A2(n537), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n567), .A2(n549), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n543) );
  NAND2_X1 U606 ( .A1(n549), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT113), .Z(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n547) );
  NAND2_X1 U611 ( .A1(n549), .A2(n585), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n563), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G134GAT), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n573), .A2(n553), .ZN(n564) );
  NOR2_X1 U619 ( .A1(n575), .A2(n564), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n557) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n488), .A2(n564), .ZN(n558) );
  XOR2_X1 U626 ( .A(n559), .B(n558), .Z(G1345GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n564), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  INV_X1 U630 ( .A(n563), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n570), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1348GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n580) );
  NOR2_X1 U640 ( .A1(n580), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  INV_X1 U646 ( .A(n580), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

