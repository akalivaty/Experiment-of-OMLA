//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G71gat), .B(G78gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT97), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n202), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n207), .A2(new_n208), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G127gat), .B(G155gat), .Z(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT20), .ZN(new_n216));
  XOR2_X1   g015(.A(new_n214), .B(new_n216), .Z(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G1gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n218), .B(KEYINPUT92), .ZN(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n228), .A3(G8gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n222), .B(new_n227), .C1(new_n223), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(KEYINPUT21), .B2(new_n211), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT99), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n217), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G183gat), .B(G211gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n235), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT89), .B(G29gat), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G36gat), .ZN(new_n241));
  INV_X1    g040(.A(G29gat), .ZN(new_n242));
  INV_X1    g041(.A(G36gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT14), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT14), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(G29gat), .B2(G36gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT88), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252));
  NOR2_X1   g051(.A1(G43gat), .A2(G50gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G43gat), .A2(G50gat), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT90), .B(G50gat), .Z(new_n258));
  OAI211_X1 g057(.A(new_n252), .B(new_n255), .C1(new_n258), .C2(G43gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n256), .A2(new_n247), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n241), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n262), .A2(KEYINPUT91), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT17), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(KEYINPUT8), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G99gat), .B(G106gat), .Z(new_n274));
  OR2_X1    g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n264), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n262), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT41), .ZN(new_n280));
  AND2_X1   g079(.A1(G232gat), .A2(G233gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n277), .A2(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT101), .ZN(new_n284));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285));
  OAI22_X1  g084(.A1(new_n278), .A2(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G134gat), .B(G162gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  OAI221_X1 g088(.A(new_n289), .B1(new_n284), .B2(new_n285), .C1(new_n278), .C2(new_n283), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n282), .A2(new_n280), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n294), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n239), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n211), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n277), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n211), .A3(new_n276), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT102), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT102), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n305), .A3(new_n301), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT10), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT10), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G230gat), .ZN(new_n310));
  INV_X1    g109(.A(G233gat), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n307), .A2(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n311), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n304), .A2(new_n313), .A3(new_n306), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n312), .A2(new_n314), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n300), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT94), .B1(new_n232), .B2(new_n262), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n232), .A2(new_n262), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G229gat), .A2(G233gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n328), .B(KEYINPUT13), .Z(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(KEYINPUT95), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n229), .A2(new_n231), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n279), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT94), .A3(new_n326), .ZN(new_n333));
  INV_X1    g132(.A(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n325), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n335), .A3(new_n329), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n334), .B1(new_n331), .B2(new_n264), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT18), .B1(new_n340), .B2(new_n328), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n264), .A2(new_n331), .ZN(new_n342));
  AND4_X1   g141(.A1(KEYINPUT18), .A2(new_n342), .A3(new_n328), .A4(new_n326), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G197gat), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT11), .B(G169gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n348), .B(KEYINPUT12), .Z(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n339), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n350), .B1(new_n339), .B2(new_n344), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355));
  NAND2_X1  g154(.A1(G211gat), .A2(G218gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT22), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(G197gat), .A2(G204gat), .ZN(new_n359));
  AND2_X1   g158(.A1(G197gat), .A2(G204gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(G211gat), .B(G218gat), .Z(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n358), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT2), .ZN(new_n369));
  INV_X1    g168(.A(G141gat), .ZN(new_n370));
  INV_X1    g169(.A(G148gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT77), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G155gat), .ZN(new_n378));
  INV_X1    g177(.A(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n381), .A3(new_n368), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n374), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n375), .A2(new_n376), .ZN(new_n384));
  AND2_X1   g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n384), .A2(new_n387), .A3(new_n381), .A4(new_n369), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n367), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n389), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n363), .B2(new_n366), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n397), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n361), .A2(new_n362), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n364), .B1(new_n358), .B2(new_n365), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n392), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT81), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n390), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n393), .B1(new_n409), .B2(new_n397), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n402), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n405), .B2(KEYINPUT81), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n389), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  OAI211_X1 g212(.A(KEYINPUT82), .B(new_n395), .C1(new_n413), .C2(new_n393), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n401), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G22gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n355), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(G78gat), .B(G106gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT80), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT31), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n420), .B(G50gat), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n411), .A2(new_n414), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n423), .B2(new_n400), .ZN(new_n424));
  AOI211_X1 g223(.A(G22gat), .B(new_n401), .C1(new_n411), .C2(new_n414), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n417), .A2(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n414), .ZN(new_n427));
  INV_X1    g226(.A(new_n408), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n390), .B1(new_n398), .B2(new_n407), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n397), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n394), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT82), .B1(new_n431), .B2(new_n395), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n400), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G22gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n416), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n355), .A4(new_n421), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G183gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT27), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT27), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G183gat), .ZN(new_n441));
  INV_X1    g240(.A(G190gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT28), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G169gat), .ZN(new_n448));
  INV_X1    g247(.A(G176gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT26), .ZN(new_n450));
  NAND2_X1  g249(.A1(G183gat), .A2(G190gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT26), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(G169gat), .B2(G176gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(G169gat), .A2(G176gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n449), .A2(KEYINPUT23), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n448), .A2(new_n449), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n454), .A2(KEYINPUT23), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n461), .A2(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT24), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n438), .A2(new_n442), .ZN(new_n468));
  NAND3_X1  g267(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT25), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n464), .A2(new_n463), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n473));
  NOR2_X1   g272(.A1(G169gat), .A2(G176gat), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(KEYINPUT23), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n468), .A2(new_n469), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT65), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n451), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT66), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT24), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n476), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n458), .B1(new_n471), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G127gat), .ZN(new_n487));
  INV_X1    g286(.A(G134gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT67), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G134gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n494), .B2(G127gat), .ZN(new_n495));
  INV_X1    g294(.A(G113gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G120gat), .ZN(new_n497));
  INV_X1    g296(.A(G120gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G113gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT1), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G120gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n500), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT70), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n507), .A2(new_n508), .A3(G113gat), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G127gat), .A2(G134gat), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT1), .B1(new_n489), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n513), .A2(new_n514), .A3(new_n496), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n510), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n506), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT71), .B1(new_n486), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n456), .B1(new_n445), .B2(new_n446), .ZN(new_n520));
  INV_X1    g319(.A(new_n460), .ZN(new_n521));
  NAND2_X1  g320(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n462), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n470), .A3(new_n472), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n473), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n484), .A2(new_n477), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n474), .B1(KEYINPUT23), .B2(new_n454), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT23), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT25), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n520), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT1), .B1(new_n504), .B2(new_n500), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n500), .B2(new_n504), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n515), .A2(new_n516), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n510), .A2(new_n512), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n534), .A2(new_n495), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n532), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n486), .A2(new_n518), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G227gat), .A2(G233gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  XNOR2_X1  g344(.A(G15gat), .B(G43gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(G71gat), .B(G99gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n544), .B(KEYINPUT32), .C1(new_n545), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n538), .B1(new_n532), .B2(new_n537), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n532), .A2(new_n537), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n542), .A3(new_n539), .ZN(new_n553));
  XNOR2_X1  g352(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT34), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n553), .A2(KEYINPUT74), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n542), .B1(new_n552), .B2(new_n539), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT73), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n548), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n562), .A3(KEYINPUT32), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT72), .B1(new_n544), .B2(new_n545), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n566), .B(KEYINPUT33), .C1(new_n541), .C2(new_n543), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI221_X1 g367(.A(new_n549), .B1(new_n555), .B2(new_n557), .C1(new_n564), .C2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n549), .B1(new_n564), .B2(new_n568), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n557), .A2(new_n555), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n437), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G8gat), .B(G36gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G64gat), .B(G92gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n486), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n581));
  INV_X1    g380(.A(G226gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n311), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT29), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n367), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n532), .A2(new_n583), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n532), .A2(KEYINPUT29), .A3(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n581), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n583), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n578), .B(new_n588), .C1(new_n591), .C2(new_n586), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT30), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G225gat), .A2(G233gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT78), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n518), .A3(new_n391), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n506), .A2(new_n389), .A3(new_n517), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n600), .A2(KEYINPUT4), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(KEYINPUT4), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n597), .B(new_n599), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n506), .A2(new_n389), .A3(new_n517), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n389), .B1(new_n517), .B2(new_n506), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT5), .B1(new_n606), .B2(new_n597), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n600), .B(KEYINPUT4), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n609), .A2(KEYINPUT5), .A3(new_n597), .A4(new_n599), .ZN(new_n610));
  XNOR2_X1  g409(.A(G1gat), .B(G29gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT0), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G85gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n608), .A2(new_n610), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(new_n614), .A3(new_n610), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n615), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n614), .B1(new_n608), .B2(new_n610), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n578), .ZN(new_n623));
  INV_X1    g422(.A(new_n583), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n580), .B2(new_n581), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n367), .B1(new_n625), .B2(new_n589), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n626), .A2(new_n627), .A3(new_n588), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n626), .B2(new_n588), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n623), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n594), .A2(new_n622), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n437), .A2(new_n572), .A3(KEYINPUT86), .A4(new_n569), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n575), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT35), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT35), .ZN(new_n636));
  AND4_X1   g435(.A1(new_n636), .A2(new_n593), .A3(new_n621), .A4(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n437), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n572), .A2(new_n569), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n572), .A2(new_n569), .A3(KEYINPUT85), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n572), .A2(new_n569), .A3(KEYINPUT36), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n609), .A2(new_n599), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n650), .A2(KEYINPUT39), .A3(new_n597), .ZN(new_n651));
  INV_X1    g450(.A(new_n614), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n606), .A2(new_n597), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n653), .B(KEYINPUT39), .C1(new_n650), .C2(new_n597), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n608), .A2(new_n610), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n655), .A2(new_n656), .B1(new_n614), .B2(new_n657), .ZN(new_n658));
  OAI221_X1 g457(.A(new_n658), .B1(new_n656), .B2(new_n655), .C1(new_n594), .C2(new_n631), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n628), .A2(new_n629), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT37), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n626), .A2(new_n661), .A3(new_n588), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(KEYINPUT38), .A3(new_n623), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n591), .A2(new_n367), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n585), .A2(new_n367), .A3(new_n587), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n623), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n662), .A2(new_n664), .B1(KEYINPUT38), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n617), .B(new_n592), .C1(new_n619), .C2(new_n620), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n659), .A2(new_n673), .A3(new_n437), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n594), .A2(new_n631), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n426), .A2(KEYINPUT84), .A3(new_n436), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT84), .B1(new_n426), .B2(new_n436), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n676), .A2(new_n622), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n649), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT87), .B1(new_n645), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n643), .B1(new_n634), .B2(KEYINPUT35), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n649), .A2(new_n674), .A3(new_n679), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT87), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n354), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(KEYINPUT96), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n645), .A2(KEYINPUT87), .A3(new_n680), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n682), .B2(new_n683), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT96), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n354), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n324), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n622), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n676), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n324), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n691), .B1(new_n690), .B2(new_n354), .ZN(new_n700));
  AOI211_X1 g499(.A(KEYINPUT96), .B(new_n353), .C1(new_n688), .C2(new_n689), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n676), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G8gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n705));
  INV_X1    g504(.A(new_n702), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT42), .B1(new_n706), .B2(new_n697), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n696), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n698), .B2(new_n703), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(new_n707), .A3(KEYINPUT103), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n709), .A2(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(new_n693), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n714), .B2(new_n649), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n641), .A2(new_n642), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n717), .A2(G15gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n715), .B1(new_n714), .B2(new_n718), .ZN(G1326gat));
  NOR2_X1   g518(.A1(new_n677), .A2(new_n678), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n693), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n723), .B2(new_n724), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(G1327gat));
  NAND2_X1  g527(.A1(new_n239), .A2(new_n323), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n298), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n700), .B2(new_n701), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n731), .A2(new_n621), .A3(new_n240), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n645), .A2(new_n680), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n735), .B2(new_n299), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n298), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n690), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n729), .A2(new_n353), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n741), .A2(KEYINPUT105), .A3(new_n621), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT105), .B1(new_n741), .B2(new_n621), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n240), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n732), .A2(new_n733), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n734), .A2(new_n744), .A3(new_n745), .ZN(G1328gat));
  NOR2_X1   g545(.A1(new_n675), .A2(G36gat), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n730), .B(new_n747), .C1(new_n700), .C2(new_n701), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G36gat), .B1(new_n741), .B2(new_n675), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(new_n754), .ZN(G1329gat));
  NOR2_X1   g554(.A1(new_n731), .A2(new_n717), .ZN(new_n756));
  INV_X1    g555(.A(new_n649), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  OAI22_X1  g557(.A1(new_n756), .A2(G43gat), .B1(new_n741), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n741), .B2(new_n437), .ZN(new_n762));
  INV_X1    g561(.A(new_n437), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n739), .A2(KEYINPUT109), .A3(new_n763), .A4(new_n740), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n258), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n731), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(KEYINPUT107), .B(new_n730), .C1(new_n700), .C2(new_n701), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n720), .A2(new_n258), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n765), .A2(new_n770), .A3(KEYINPUT48), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n258), .B1(new_n741), .B2(new_n720), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT48), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT108), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n776), .B(KEYINPUT48), .C1(new_n770), .C2(new_n772), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n771), .B1(new_n775), .B2(new_n777), .ZN(G1331gat));
  NAND4_X1  g577(.A1(new_n735), .A2(new_n353), .A3(new_n300), .A4(new_n322), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n622), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n676), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT49), .B(G64gat), .Z(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(G1333gat));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n204), .A3(new_n716), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n780), .A2(new_n757), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n204), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1334gat));
  NAND2_X1  g590(.A1(new_n780), .A2(new_n721), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(G78gat), .ZN(G1335gat));
  INV_X1    g592(.A(new_n239), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(new_n354), .A3(new_n323), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n739), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n621), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n735), .A2(new_n353), .A3(new_n239), .A4(new_n299), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n322), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n622), .A2(new_n270), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(G1336gat));
  NOR3_X1   g604(.A1(new_n323), .A2(new_n675), .A3(G92gat), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n739), .A2(new_n676), .A3(new_n795), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G92gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n806), .B(KEYINPUT112), .Z(new_n811));
  AOI22_X1  g610(.A1(new_n808), .A2(G92gat), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n796), .B2(new_n649), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n717), .A2(G99gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n803), .B2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(new_n803), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n437), .A2(G106gat), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G106gat), .B1(new_n796), .B2(new_n437), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT53), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g622(.A(KEYINPUT53), .B(G106gat), .C1(new_n796), .C2(new_n720), .ZN(new_n824));
  NOR2_X1   g623(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n818), .B2(new_n820), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n823), .B1(new_n824), .B2(new_n826), .ZN(G1339gat));
  NAND2_X1  g626(.A1(new_n699), .A2(new_n353), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n339), .A2(new_n344), .A3(new_n350), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n329), .B1(new_n333), .B2(new_n335), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n830), .A2(new_n831), .B1(new_n328), .B2(new_n340), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n327), .A2(KEYINPUT115), .A3(new_n329), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n348), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n296), .A2(new_n829), .A3(new_n834), .A4(new_n297), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n307), .A2(new_n309), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n313), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n312), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n319), .B1(new_n312), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n836), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n843), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n321), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n835), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n834), .A3(new_n322), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n353), .B2(new_n847), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n298), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n239), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g652(.A(KEYINPUT116), .B(new_n848), .C1(new_n298), .C2(new_n850), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n828), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n676), .A2(new_n621), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n717), .A2(new_n721), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n858), .A2(new_n496), .A3(new_n353), .ZN(new_n859));
  INV_X1    g658(.A(new_n855), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n575), .A2(new_n633), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n860), .A2(new_n621), .A3(new_n676), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n354), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n496), .ZN(G1340gat));
  NAND4_X1  g663(.A1(new_n862), .A2(new_n507), .A3(new_n509), .A4(new_n322), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n858), .B2(new_n323), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1341gat));
  NAND3_X1  g666(.A1(new_n862), .A2(new_n487), .A3(new_n794), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n858), .B2(new_n239), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  NAND4_X1  g669(.A1(new_n862), .A2(new_n491), .A3(new_n493), .A4(new_n299), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n858), .B2(new_n298), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n621), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n757), .A2(new_n437), .A3(new_n676), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n353), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n855), .A2(new_n763), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n649), .A2(new_n856), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n828), .B1(new_n794), .B2(new_n851), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n721), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n884), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(new_n354), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G141gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n880), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n888), .A2(G141gat), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT58), .B1(new_n893), .B2(new_n879), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(new_n878), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n371), .A3(new_n322), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n886), .A2(new_n882), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(new_n649), .A3(new_n322), .A4(new_n856), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n898), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n883), .A2(new_n887), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n371), .C1(new_n904), .C2(new_n322), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n897), .B1(new_n903), .B2(new_n905), .ZN(G1345gat));
  NOR3_X1   g705(.A1(new_n878), .A2(G155gat), .A3(new_n239), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n904), .A2(new_n794), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT118), .B(new_n908), .C1(new_n909), .C2(new_n378), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n378), .B1(new_n904), .B2(new_n794), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n896), .B2(new_n299), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n298), .A2(new_n379), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n904), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n860), .A2(new_n622), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n861), .A2(new_n675), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n354), .A3(new_n461), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(KEYINPUT119), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n675), .A2(new_n622), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n855), .A2(new_n857), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT120), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n855), .A2(new_n927), .A3(new_n857), .A4(new_n924), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n926), .A2(new_n354), .A3(new_n928), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n922), .A2(new_n923), .B1(new_n448), .B2(new_n929), .ZN(G1348gat));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n449), .A3(new_n322), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n926), .A2(new_n322), .A3(new_n928), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n449), .B2(new_n932), .ZN(G1349gat));
  NAND3_X1  g732(.A1(new_n926), .A2(new_n794), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n794), .A2(new_n439), .A3(new_n441), .ZN(new_n936));
  AND4_X1   g735(.A1(new_n621), .A2(new_n855), .A3(new_n919), .A4(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n939), .B2(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n937), .B1(new_n934), .B2(G183gat), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n941), .A2(new_n945), .A3(new_n943), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n941), .B2(new_n943), .ZN(new_n947));
  OAI22_X1  g746(.A1(new_n940), .A2(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n926), .A2(new_n299), .A3(new_n928), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G190gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n952), .A3(G190gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(KEYINPUT61), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n920), .A2(new_n442), .A3(new_n299), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n954), .B(new_n955), .C1(KEYINPUT61), .C2(new_n951), .ZN(G1351gat));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n649), .A2(new_n924), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n958), .B1(new_n899), .B2(new_n900), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n960), .B2(new_n353), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(KEYINPUT125), .A3(new_n354), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(G197gat), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n649), .A2(new_n763), .A3(new_n676), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT124), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n918), .A2(new_n965), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n966), .A2(G197gat), .A3(new_n353), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n963), .A2(new_n967), .ZN(G1352gat));
  OAI21_X1  g767(.A(G204gat), .B1(new_n960), .B2(new_n323), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n323), .A2(G204gat), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  OR3_X1    g770(.A1(new_n966), .A2(KEYINPUT126), .A3(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT126), .B1(new_n966), .B2(new_n971), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n973), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(G1353gat));
  OR3_X1    g776(.A1(new_n966), .A2(G211gat), .A3(new_n239), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n959), .A2(new_n794), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  AND2_X1   g781(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n299), .B1(new_n959), .B2(KEYINPUT127), .ZN(new_n984));
  OAI21_X1  g783(.A(G218gat), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n298), .A2(G218gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n966), .B2(new_n986), .ZN(G1355gat));
endmodule


