//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  AND2_X1   g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g005(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT76), .A2(G211gat), .ZN(new_n208));
  OAI21_X1  g007(.A(G218gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n203), .B1(new_n211), .B2(KEYINPUT77), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT76), .B(G211gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT22), .B1(new_n214), .B2(G218gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n213), .B(new_n202), .C1(new_n215), .C2(new_n206), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G226gat), .A2(G233gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n227));
  INV_X1    g026(.A(G169gat), .ZN(new_n228));
  INV_X1    g027(.A(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n222), .A2(new_n227), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n238));
  AND2_X1   g037(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n232), .B1(KEYINPUT23), .B2(new_n234), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n228), .ZN(new_n247));
  NAND2_X1  g046(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT23), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n230), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n225), .A2(KEYINPUT24), .ZN(new_n254));
  XOR2_X1   g053(.A(G183gat), .B(G190gat), .Z(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(KEYINPUT24), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n243), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n232), .B2(KEYINPUT23), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n254), .ZN(new_n262));
  XNOR2_X1  g061(.A(G183gat), .B(G190gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT24), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n265), .B2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n262), .B(new_n267), .C1(new_n263), .C2(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n237), .B1(new_n259), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n219), .B1(new_n270), .B2(KEYINPUT29), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272));
  INV_X1    g071(.A(new_n219), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n257), .A2(new_n258), .B1(new_n266), .B2(new_n268), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(new_n237), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n226), .A2(new_n236), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n252), .B1(new_n249), .B2(new_n251), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n265), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT25), .B1(new_n279), .B2(new_n253), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g080(.A(new_n261), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n281), .A2(new_n268), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n277), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n272), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n218), .B(new_n271), .C1(new_n276), .C2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  OAI21_X1  g088(.A(KEYINPUT79), .B1(new_n270), .B2(new_n219), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n291), .B(new_n273), .C1(new_n274), .C2(new_n237), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n274), .B2(new_n237), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n290), .A2(new_n292), .B1(new_n219), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n286), .B(new_n289), .C1(new_n295), .C2(new_n218), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n295), .B2(new_n218), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT37), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n290), .A2(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n219), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n217), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n289), .B1(new_n303), .B2(new_n286), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n299), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n297), .B1(new_n307), .B2(KEYINPUT38), .ZN(new_n308));
  AOI221_X4 g107(.A(new_n217), .B1(new_n294), .B2(new_n219), .C1(new_n290), .C2(new_n292), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n271), .B1(new_n276), .B2(new_n285), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n217), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT91), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(KEYINPUT91), .A3(new_n217), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT38), .ZN(new_n316));
  INV_X1    g115(.A(new_n289), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n316), .B(new_n317), .C1(new_n298), .C2(KEYINPUT37), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT92), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT86), .B(KEYINPUT6), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n323));
  INV_X1    g122(.A(G141gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(G148gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G148gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT82), .A3(G141gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT83), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n329), .A2(new_n335), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G141gat), .B(G148gat), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n334), .B(new_n332), .C1(new_n341), .C2(KEYINPUT2), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G134gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G127gat), .ZN(new_n345));
  INV_X1    g144(.A(G127gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G134gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(G127gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G134gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(G113gat), .A2(G120gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(G113gat), .A2(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT69), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT1), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(KEYINPUT69), .A3(new_n354), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n352), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G113gat), .A2(G120gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n364));
  OR2_X1    g163(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n365));
  AND4_X1   g164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n343), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT1), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n358), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n363), .A2(new_n348), .B1(G134gat), .B2(new_n350), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND4_X1   g171(.A1(new_n345), .A2(new_n365), .A3(new_n347), .A4(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n362), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n372), .A2(new_n342), .A3(new_n340), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G225gat), .A2(G233gat), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n322), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n340), .A2(new_n381), .A3(new_n342), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(new_n374), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n340), .A2(new_n342), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n370), .A2(new_n371), .B1(new_n373), .B2(new_n362), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n377), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n379), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT84), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n379), .A2(new_n390), .A3(KEYINPUT84), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(G1gat), .B(G29gat), .Z(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(new_n390), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(new_n322), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n321), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n322), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n379), .A2(new_n390), .A3(KEYINPUT84), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT84), .B1(new_n379), .B2(new_n390), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n400), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT90), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n400), .A3(new_n321), .ZN(new_n410));
  INV_X1    g209(.A(new_n400), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n395), .B2(new_n404), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n320), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n415), .B2(KEYINPUT90), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT29), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n273), .B1(new_n284), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT80), .B1(new_n270), .B2(new_n219), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n275), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n312), .B1(new_n420), .B2(new_n218), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n295), .A2(new_n218), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n314), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n298), .A2(new_n317), .ZN(new_n425));
  INV_X1    g224(.A(new_n306), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .A4(new_n316), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n308), .A2(new_n319), .A3(new_n416), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n382), .A2(new_n293), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n217), .ZN(new_n432));
  INV_X1    g231(.A(G228gat), .ZN(new_n433));
  INV_X1    g232(.A(G233gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n212), .A2(new_n216), .A3(new_n417), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n387), .B1(new_n437), .B2(new_n381), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT87), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n381), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n343), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n442));
  INV_X1    g241(.A(new_n435), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n431), .B2(new_n217), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n293), .B1(new_n211), .B2(new_n203), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n215), .A2(new_n206), .A3(new_n202), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n381), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n343), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n435), .B1(new_n450), .B2(new_n432), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(G22gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(new_n455), .A3(new_n452), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(KEYINPUT88), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT88), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n446), .B2(new_n452), .ZN(new_n459));
  AOI211_X1 g258(.A(G22gat), .B(new_n451), .C1(new_n439), .C2(new_n445), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G50gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n459), .A2(new_n460), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(KEYINPUT88), .A3(new_n464), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT30), .B1(new_n297), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n296), .A2(KEYINPUT81), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n473), .A3(new_n425), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n378), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n476), .A2(KEYINPUT39), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n476), .B(KEYINPUT39), .C1(new_n378), .C2(new_n376), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n478), .A3(new_n411), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT89), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT40), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n479), .B(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n412), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n469), .B1(new_n474), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n471), .A2(new_n415), .A3(new_n473), .A4(new_n425), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n430), .A2(new_n484), .B1(new_n485), .B2(new_n469), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n388), .B1(new_n274), .B2(new_n237), .ZN(new_n491));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n383), .B(new_n277), .C1(new_n280), .C2(new_n283), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(new_n495), .B2(KEYINPUT32), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT33), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n495), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n487), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(KEYINPUT72), .A3(new_n499), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n493), .B1(new_n491), .B2(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n495), .B(KEYINPUT32), .C1(new_n498), .C2(new_n490), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n509), .B2(new_n511), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(KEYINPUT74), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n505), .A2(new_n513), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT75), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(new_n515), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n512), .B1(new_n505), .B2(new_n513), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n513), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n519), .A2(new_n518), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n505), .B2(new_n514), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n521), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  NOR4_X1   g331(.A1(new_n459), .A2(new_n460), .A3(new_n458), .A4(new_n465), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n464), .B1(new_n467), .B2(KEYINPUT88), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n461), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n535), .A3(new_n515), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT35), .B1(new_n536), .B2(new_n485), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n524), .ZN(new_n539));
  INV_X1    g338(.A(new_n416), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n535), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n486), .A2(new_n532), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT14), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n544), .A2(KEYINPUT93), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(KEYINPUT93), .B2(new_n544), .ZN(new_n546));
  XOR2_X1   g345(.A(G43gat), .B(G50gat), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n544), .A2(KEYINPUT95), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n547), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT15), .B1(new_n547), .B2(KEYINPUT94), .ZN(new_n552));
  OAI221_X1 g351(.A(new_n550), .B1(KEYINPUT95), .B2(new_n544), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(G1gat), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(G1gat), .B2(new_n555), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(G8gat), .Z(new_n559));
  NOR2_X1   g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n559), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n549), .A2(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT17), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n560), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n565), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n564), .A2(KEYINPUT17), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n559), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n568), .A2(new_n573), .A3(KEYINPUT18), .A4(new_n569), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n561), .B(new_n564), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n569), .B(KEYINPUT13), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G197gat), .ZN(new_n583));
  XOR2_X1   g382(.A(KEYINPUT11), .B(G169gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT12), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n576), .A2(new_n588), .A3(new_n577), .A4(new_n580), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT97), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(KEYINPUT97), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(KEYINPUT97), .B(new_n591), .C1(new_n594), .C2(new_n593), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n559), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n602), .B(KEYINPUT98), .Z(new_n603));
  NOR2_X1   g402(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n606), .A2(G127gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(G127gat), .ZN(new_n608));
  OR3_X1    g407(.A1(new_n603), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n330), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n610), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G99gat), .B(G106gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n629), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n636), .B1(new_n570), .B2(new_n571), .ZN(new_n637));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n564), .A3(new_n635), .ZN(new_n640));
  NAND3_X1  g439(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n638), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n642), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n650), .A2(KEYINPUT101), .A3(new_n642), .A4(new_n647), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n619), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n634), .A2(new_n600), .A3(new_n628), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n636), .B2(new_n600), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n659), .A2(KEYINPUT103), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(KEYINPUT103), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(new_n663), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n660), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  AOI211_X1 g465(.A(KEYINPUT10), .B(new_n656), .C1(new_n636), .C2(new_n600), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n600), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n632), .A2(new_n635), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n632), .A2(KEYINPUT102), .A3(new_n635), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n658), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n658), .B2(new_n657), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n664), .B(KEYINPUT104), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n666), .A2(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n542), .A2(new_n590), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n415), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g482(.A1(new_n680), .A2(new_n474), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G8gat), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n689), .A2(KEYINPUT105), .A3(new_n687), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n689), .B2(new_n687), .ZN(new_n691));
  OAI221_X1 g490(.A(new_n686), .B1(new_n687), .B2(new_n689), .C1(new_n690), .C2(new_n691), .ZN(G1325gat));
  NOR2_X1   g491(.A1(new_n542), .A2(new_n590), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n539), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n694), .A2(G15gat), .A3(new_n679), .ZN(new_n695));
  INV_X1    g494(.A(new_n532), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(G15gat), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT106), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n469), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(new_n653), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n644), .A2(new_n647), .B1(new_n650), .B2(new_n642), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n430), .A2(new_n484), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n485), .A2(new_n469), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n532), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n537), .A2(new_n541), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n678), .ZN(new_n711));
  INV_X1    g510(.A(new_n619), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n590), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(G29gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n681), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n542), .B2(new_n705), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n708), .A2(new_n709), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .A3(new_n654), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n713), .B(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724), .B2(new_n415), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n725), .ZN(G1328gat));
  INV_X1    g525(.A(new_n474), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n712), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n654), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  AOI21_X1  g531(.A(G36gat), .B1(new_n732), .B2(KEYINPUT46), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n693), .A2(new_n474), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n728), .A2(new_n736), .ZN(G1329gat));
  OAI21_X1  g536(.A(G43gat), .B1(new_n724), .B2(new_n532), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT47), .B1(new_n738), .B2(KEYINPUT109), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n694), .A2(G43gat), .A3(new_n730), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n738), .B(new_n740), .C1(KEYINPUT109), .C2(KEYINPUT47), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n722), .A2(new_n469), .A3(new_n723), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  INV_X1    g546(.A(G50gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n714), .A2(new_n748), .A3(new_n469), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1331gat));
  AND4_X1   g551(.A1(new_n720), .A2(new_n590), .A3(new_n655), .A4(new_n711), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n681), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(G57gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1332gat));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n474), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT49), .B(G64gat), .Z(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n757), .B2(new_n759), .ZN(G1333gat));
  NAND2_X1  g559(.A1(new_n753), .A2(new_n696), .ZN(new_n761));
  INV_X1    g560(.A(new_n539), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(G71gat), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n761), .A2(G71gat), .B1(new_n753), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n753), .A2(new_n469), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n542), .B2(new_n705), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n720), .A2(KEYINPUT114), .A3(new_n654), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n590), .A2(new_n771), .A3(new_n619), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n587), .A2(new_n589), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT112), .B1(new_n712), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AND4_X1   g575(.A1(KEYINPUT51), .A2(new_n769), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT115), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n775), .B1(new_n710), .B2(KEYINPUT114), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n769), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n779), .B2(new_n769), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n778), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n623), .A3(new_n681), .A4(new_n711), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n775), .A2(new_n678), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n719), .A2(new_n721), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT113), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n719), .A2(new_n721), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n681), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n786), .B1(new_n623), .B2(new_n792), .ZN(G1336gat));
  NOR3_X1   g592(.A1(new_n678), .A2(G92gat), .A3(new_n727), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT116), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n777), .B2(new_n783), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n798), .B(new_n795), .C1(new_n777), .C2(new_n783), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n789), .A2(new_n474), .A3(new_n791), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G92gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n795), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n722), .A2(new_n474), .A3(new_n787), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n805), .B2(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1337gat));
  NOR3_X1   g607(.A1(new_n762), .A2(new_n678), .A3(G99gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n789), .A2(new_n696), .A3(new_n791), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G99gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  NOR3_X1   g612(.A1(new_n678), .A2(G106gat), .A3(new_n535), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n785), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n722), .A2(new_n469), .A3(new_n787), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n816), .B2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n784), .A2(new_n780), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n789), .A2(new_n469), .A3(new_n791), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n820), .A2(new_n814), .B1(new_n821), .B2(G106gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n818), .B1(new_n819), .B2(new_n822), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n679), .A2(new_n773), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n657), .A2(new_n668), .ZN(new_n825));
  INV_X1    g624(.A(new_n658), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n673), .A4(new_n672), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n675), .A2(new_n827), .A3(KEYINPUT54), .ZN(new_n828));
  XOR2_X1   g627(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n829));
  OAI211_X1 g628(.A(new_n658), .B(new_n829), .C1(new_n667), .C2(new_n674), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n665), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT55), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n675), .A2(new_n827), .A3(KEYINPUT54), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n665), .A4(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n705), .A2(new_n587), .A3(new_n589), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n666), .A2(new_n675), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n569), .B1(new_n568), .B2(new_n573), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n578), .A2(new_n579), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n585), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n589), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n654), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n836), .A2(new_n837), .A3(new_n838), .A4(new_n843), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n678), .A2(new_n842), .A3(new_n654), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n824), .B1(new_n846), .B2(new_n619), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n474), .A2(new_n415), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n762), .A2(new_n469), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n590), .ZN(new_n853));
  INV_X1    g652(.A(new_n536), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n590), .A2(G113gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT119), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n852), .A2(new_n859), .A3(new_n678), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n850), .A2(new_n854), .A3(new_n711), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n852), .B2(new_n619), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n712), .A2(new_n346), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n855), .B2(new_n864), .ZN(G1342gat));
  AND4_X1   g664(.A1(new_n344), .A2(new_n850), .A3(new_n854), .A4(new_n654), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT120), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n851), .A3(new_n654), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n866), .A2(new_n867), .B1(G134gat), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n696), .A2(new_n535), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n850), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n324), .A3(new_n773), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n532), .A2(new_n848), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n847), .B2(new_n535), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n712), .B1(new_n844), .B2(new_n845), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT57), .B(new_n469), .C1(new_n879), .C2(new_n824), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n590), .B(new_n876), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n875), .B1(new_n881), .B2(new_n324), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT121), .B1(new_n881), .B2(new_n324), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OAI221_X1 g684(.A(new_n875), .B1(KEYINPUT121), .B2(KEYINPUT58), .C1(new_n881), .C2(new_n324), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n327), .A3(new_n711), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n876), .B1(new_n878), .B2(new_n880), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n711), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n327), .C1(new_n890), .C2(new_n711), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n874), .A2(new_n712), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n712), .A2(G155gat), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n895), .A2(new_n330), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT123), .ZN(G1346gat));
  AOI21_X1  g698(.A(G162gat), .B1(new_n874), .B2(new_n654), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n705), .A2(new_n331), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n890), .B2(new_n901), .ZN(G1347gat));
  NOR2_X1   g701(.A1(new_n847), .A2(new_n681), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n762), .A2(new_n727), .A3(new_n469), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n590), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n847), .A2(new_n681), .A3(new_n727), .A4(new_n536), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n907), .A2(new_n247), .A3(new_n248), .A4(new_n773), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1348gat));
  OAI21_X1  g708(.A(G176gat), .B1(new_n905), .B2(new_n678), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n907), .A2(new_n229), .A3(new_n711), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1349gat));
  OAI21_X1  g711(.A(G183gat), .B1(new_n905), .B2(new_n619), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n907), .A2(new_n220), .A3(new_n712), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g715(.A1(new_n907), .A2(new_n221), .A3(new_n654), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n903), .A2(new_n654), .A3(new_n904), .ZN(new_n918));
  NOR2_X1   g717(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n221), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(G1351gat));
  AND3_X1   g723(.A1(new_n903), .A2(new_n474), .A3(new_n873), .ZN(new_n925));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n773), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n532), .A2(new_n415), .A3(new_n474), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n878), .B2(new_n880), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n773), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  XOR2_X1   g731(.A(KEYINPUT126), .B(G204gat), .Z(new_n933));
  NOR2_X1   g732(.A1(new_n678), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n925), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT127), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(KEYINPUT127), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(new_n711), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n933), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n939), .B(new_n941), .C1(new_n937), .C2(new_n935), .ZN(G1353gat));
  INV_X1    g741(.A(new_n214), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n943), .A3(new_n712), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n930), .A2(new_n712), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  INV_X1    g747(.A(G218gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n925), .A2(new_n949), .A3(new_n654), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n930), .A2(new_n654), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n949), .ZN(G1355gat));
endmodule


