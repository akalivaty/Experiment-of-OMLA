

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U323 ( .A(n394), .B(KEYINPUT64), .ZN(n395) );
  XNOR2_X1 U324 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U325 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U326 ( .A(n352), .B(n295), .ZN(n298) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n411) );
  XNOR2_X1 U328 ( .A(n412), .B(n411), .ZN(n570) );
  XNOR2_X1 U329 ( .A(n396), .B(n395), .ZN(n541) );
  XNOR2_X1 U330 ( .A(n311), .B(n310), .ZN(n554) );
  XNOR2_X1 U331 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(G92GAT), .B(G85GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(G99GAT), .B(G106GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n352) );
  NAND2_X1 U336 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  INV_X1 U337 ( .A(KEYINPUT76), .ZN(n293) );
  INV_X1 U338 ( .A(n298), .ZN(n296) );
  NAND2_X1 U339 ( .A1(n296), .A2(KEYINPUT11), .ZN(n300) );
  INV_X1 U340 ( .A(KEYINPUT11), .ZN(n297) );
  NAND2_X1 U341 ( .A1(n298), .A2(n297), .ZN(n299) );
  NAND2_X1 U342 ( .A1(n300), .A2(n299), .ZN(n302) );
  XOR2_X1 U343 ( .A(G50GAT), .B(G162GAT), .Z(n435) );
  XNOR2_X1 U344 ( .A(n435), .B(KEYINPUT65), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n311) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G43GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n373) );
  XNOR2_X1 U349 ( .A(G36GAT), .B(G190GAT), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n305), .B(G218GAT), .ZN(n404) );
  XNOR2_X1 U351 ( .A(n373), .B(n404), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n307) );
  XNOR2_X1 U353 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n306) );
  XOR2_X1 U354 ( .A(n307), .B(n306), .Z(n308) );
  XNOR2_X1 U355 ( .A(KEYINPUT78), .B(n554), .ZN(n533) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G127GAT), .Z(n338) );
  XOR2_X1 U357 ( .A(n338), .B(G71GAT), .Z(n313) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U360 ( .A(n314), .B(G99GAT), .Z(n319) );
  XOR2_X1 U361 ( .A(KEYINPUT84), .B(G134GAT), .Z(n316) );
  XNOR2_X1 U362 ( .A(KEYINPUT83), .B(G120GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(KEYINPUT0), .B(n317), .Z(n419) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(n419), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U367 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n321) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(G190GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U370 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U371 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n325) );
  XNOR2_X1 U372 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U374 ( .A(G169GAT), .B(n326), .Z(n408) );
  XOR2_X1 U375 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n328) );
  XNOR2_X1 U376 ( .A(G176GAT), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n408), .B(n329), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n521) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n333) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(KEYINPUT13), .B(n334), .Z(n353) );
  XOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n336) );
  XNOR2_X1 U385 ( .A(G1GAT), .B(G64GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U387 ( .A(n338), .B(n337), .Z(n340) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U389 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U390 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n342) );
  XNOR2_X1 U391 ( .A(KEYINPUT14), .B(KEYINPUT79), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U393 ( .A(n344), .B(n343), .Z(n348) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(G155GAT), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n345), .B(G78GAT), .ZN(n436) );
  XNOR2_X1 U396 ( .A(G8GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n346), .B(G211GAT), .ZN(n399) );
  XNOR2_X1 U398 ( .A(n436), .B(n399), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U400 ( .A(n353), .B(n349), .Z(n548) );
  INV_X1 U401 ( .A(n548), .ZN(n581) );
  XNOR2_X1 U402 ( .A(n533), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U403 ( .A1(n581), .A2(n584), .ZN(n351) );
  XOR2_X1 U404 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n385) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n355) );
  XOR2_X1 U407 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n361) );
  XOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT74), .Z(n357) );
  XNOR2_X1 U410 ( .A(G176GAT), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n401) );
  XOR2_X1 U412 ( .A(G78GAT), .B(n401), .Z(n359) );
  NAND2_X1 U413 ( .A1(G230GAT), .A2(G233GAT), .ZN(n358) );
  XOR2_X1 U414 ( .A(n359), .B(n358), .Z(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n366) );
  XOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n363) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(KEYINPUT75), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U419 ( .A(G148GAT), .B(n364), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n578) );
  XOR2_X1 U421 ( .A(G113GAT), .B(G1GAT), .Z(n415) );
  XOR2_X1 U422 ( .A(G141GAT), .B(G197GAT), .Z(n368) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(G36GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n415), .B(n369), .Z(n371) );
  NAND2_X1 U426 ( .A1(G229GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(n372), .B(KEYINPUT69), .Z(n375) );
  XNOR2_X1 U429 ( .A(n373), .B(KEYINPUT30), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n383) );
  XOR2_X1 U431 ( .A(KEYINPUT68), .B(G15GAT), .Z(n377) );
  XNOR2_X1 U432 ( .A(G169GAT), .B(G22GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n379) );
  XNOR2_X1 U435 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n382) );
  XOR2_X1 U438 ( .A(n383), .B(n382), .Z(n542) );
  INV_X1 U439 ( .A(n542), .ZN(n574) );
  AND2_X1 U440 ( .A1(n578), .A2(n574), .ZN(n384) );
  AND2_X1 U441 ( .A1(n385), .A2(n384), .ZN(n393) );
  XNOR2_X1 U442 ( .A(n578), .B(KEYINPUT41), .ZN(n560) );
  NAND2_X1 U443 ( .A1(n542), .A2(n560), .ZN(n387) );
  XOR2_X1 U444 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n386) );
  XOR2_X1 U445 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U446 ( .A(KEYINPUT109), .B(n548), .Z(n566) );
  INV_X1 U447 ( .A(n554), .ZN(n388) );
  NOR2_X1 U448 ( .A1(n566), .A2(n388), .ZN(n389) );
  NAND2_X1 U449 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(KEYINPUT47), .ZN(n392) );
  NOR2_X1 U451 ( .A1(n393), .A2(n392), .ZN(n396) );
  INV_X1 U452 ( .A(KEYINPUT48), .ZN(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n398) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U456 ( .A(n400), .B(n399), .Z(n403) );
  XNOR2_X1 U457 ( .A(n401), .B(G92GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U459 ( .A(n405), .B(n404), .Z(n410) );
  XOR2_X1 U460 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n407) );
  XNOR2_X1 U461 ( .A(G197GAT), .B(KEYINPUT90), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n445) );
  XNOR2_X1 U463 ( .A(n408), .B(n445), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n511) );
  NAND2_X1 U465 ( .A1(n541), .A2(n511), .ZN(n412) );
  XOR2_X1 U466 ( .A(G148GAT), .B(KEYINPUT2), .Z(n414) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n444) );
  XOR2_X1 U469 ( .A(G85GAT), .B(n444), .Z(n417) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(n415), .ZN(n416) );
  XNOR2_X1 U471 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n432) );
  XOR2_X1 U473 ( .A(KEYINPUT4), .B(G155GAT), .Z(n421) );
  XNOR2_X1 U474 ( .A(G127GAT), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U476 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n423) );
  XNOR2_X1 U477 ( .A(KEYINPUT6), .B(G57GAT), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U479 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n427) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT94), .B(n428), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U485 ( .A(n432), .B(n431), .Z(n469) );
  XOR2_X1 U486 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n434) );
  XNOR2_X1 U487 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n440) );
  XOR2_X1 U489 ( .A(n436), .B(n435), .Z(n438) );
  XNOR2_X1 U490 ( .A(G218GAT), .B(G106GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n449) );
  XOR2_X1 U493 ( .A(KEYINPUT23), .B(G211GAT), .Z(n442) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U496 ( .A(n443), .B(G204GAT), .Z(n447) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n463) );
  NAND2_X1 U500 ( .A1(n469), .A2(n463), .ZN(n450) );
  OR2_X1 U501 ( .A1(n570), .A2(n450), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n453) );
  NAND2_X1 U504 ( .A1(n521), .A2(n453), .ZN(n559) );
  NOR2_X1 U505 ( .A1(n533), .A2(n559), .ZN(n456) );
  XNOR2_X1 U506 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n454) );
  INV_X1 U507 ( .A(n469), .ZN(n571) );
  XNOR2_X1 U508 ( .A(n511), .B(KEYINPUT27), .ZN(n465) );
  AND2_X1 U509 ( .A1(n465), .A2(n571), .ZN(n539) );
  XNOR2_X1 U510 ( .A(n463), .B(KEYINPUT66), .ZN(n457) );
  XOR2_X1 U511 ( .A(n457), .B(KEYINPUT28), .Z(n515) );
  INV_X1 U512 ( .A(n515), .ZN(n458) );
  NAND2_X1 U513 ( .A1(n539), .A2(n458), .ZN(n523) );
  NOR2_X1 U514 ( .A1(n521), .A2(n523), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT98), .B(n459), .Z(n471) );
  NAND2_X1 U516 ( .A1(n511), .A2(n521), .ZN(n460) );
  NAND2_X1 U517 ( .A1(n460), .A2(n463), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n461), .B(KEYINPUT25), .ZN(n462) );
  XNOR2_X1 U519 ( .A(n462), .B(KEYINPUT99), .ZN(n467) );
  NOR2_X1 U520 ( .A1(n463), .A2(n521), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n464), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U522 ( .A1(n465), .A2(n572), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n483) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n473) );
  NAND2_X1 U527 ( .A1(n548), .A2(n533), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n473), .B(n472), .ZN(n474) );
  NAND2_X1 U529 ( .A1(n483), .A2(n474), .ZN(n475) );
  XNOR2_X1 U530 ( .A(n475), .B(KEYINPUT100), .ZN(n498) );
  NAND2_X1 U531 ( .A1(n542), .A2(n578), .ZN(n486) );
  NOR2_X1 U532 ( .A1(n498), .A2(n486), .ZN(n481) );
  NAND2_X1 U533 ( .A1(n571), .A2(n481), .ZN(n476) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U536 ( .A1(n481), .A2(n511), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U538 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U539 ( .A1(n481), .A2(n521), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U541 ( .A1(n515), .A2(n481), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n581), .A2(n483), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n484), .A2(n584), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(KEYINPUT37), .ZN(n509) );
  NOR2_X1 U546 ( .A1(n509), .A2(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(n489), .Z(n496) );
  NAND2_X1 U550 ( .A1(n496), .A2(n571), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n496), .A2(n511), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n521), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NAND2_X1 U559 ( .A1(n515), .A2(n496), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n500) );
  NAND2_X1 U562 ( .A1(n574), .A2(n560), .ZN(n508) );
  NOR2_X1 U563 ( .A1(n498), .A2(n508), .ZN(n504) );
  NAND2_X1 U564 ( .A1(n504), .A2(n571), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n501), .Z(G1332GAT) );
  NAND2_X1 U567 ( .A1(n504), .A2(n511), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n502), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n504), .A2(n521), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n503), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n515), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n571), .A2(n516), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n516), .A2(n511), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n516), .A2(n521), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n513), .B(KEYINPUT106), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n518) );
  NAND2_X1 U585 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U588 ( .A1(n521), .A2(n541), .ZN(n522) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n532), .A2(n542), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT112), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U594 ( .A1(n532), .A2(n560), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n529) );
  NAND2_X1 U598 ( .A1(n532), .A2(n566), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(G1342GAT) );
  INV_X1 U601 ( .A(n532), .ZN(n534) );
  NOR2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n538) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n536) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT115), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  XOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT117), .Z(n544) );
  AND2_X1 U608 ( .A1(n539), .A2(n572), .ZN(n540) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n553) );
  INV_X1 U610 ( .A(n553), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U614 ( .A1(n549), .A2(n560), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n555), .Z(G1347GAT) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n574), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n556), .B(KEYINPUT123), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  INV_X1 U627 ( .A(n559), .ZN(n567) );
  AND2_X1 U628 ( .A1(n560), .A2(n567), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n562) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n561) );
  XNOR2_X1 U631 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(KEYINPUT124), .B(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT126), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(n569), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n574), .A2(n583), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n583), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

