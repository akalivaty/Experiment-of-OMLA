

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732;

  INV_X2 U371 ( .A(G953), .ZN(n723) );
  XNOR2_X2 U372 ( .A(n515), .B(n514), .ZN(n679) );
  NAND2_X1 U373 ( .A1(n360), .A2(KEYINPUT34), .ZN(n359) );
  AND2_X2 U374 ( .A1(n598), .A2(n597), .ZN(n703) );
  NAND2_X1 U375 ( .A1(n351), .A2(n347), .ZN(n722) );
  AND2_X1 U376 ( .A1(n364), .A2(n362), .ZN(n361) );
  AND2_X1 U377 ( .A1(n365), .A2(n520), .ZN(n364) );
  BUF_X1 U378 ( .A(n516), .Z(n531) );
  OR2_X1 U379 ( .A1(n571), .A2(n550), .ZN(n499) );
  OR2_X1 U380 ( .A1(n652), .A2(n554), .ZN(n556) );
  OR2_X1 U381 ( .A1(n652), .A2(n489), .ZN(n491) );
  XNOR2_X1 U382 ( .A(n472), .B(n471), .ZN(n493) );
  AND2_X1 U383 ( .A1(n358), .A2(n357), .ZN(n356) );
  XNOR2_X1 U384 ( .A(n368), .B(G101), .ZN(n445) );
  INV_X1 U385 ( .A(n722), .ZN(n350) );
  XNOR2_X1 U386 ( .A(n549), .B(KEYINPUT84), .ZN(n352) );
  OR2_X1 U387 ( .A1(n608), .A2(G902), .ZN(n456) );
  XNOR2_X1 U388 ( .A(KEYINPUT69), .B(G131), .ZN(n440) );
  NOR2_X1 U389 ( .A1(n731), .A2(n606), .ZN(n565) );
  AND2_X1 U390 ( .A1(n531), .A2(n517), .ZN(n363) );
  NAND2_X1 U391 ( .A1(n366), .A2(KEYINPUT34), .ZN(n365) );
  NAND2_X2 U392 ( .A1(n356), .A2(n353), .ZN(n557) );
  OR2_X1 U393 ( .A1(n599), .A2(n354), .ZN(n353) );
  NAND2_X1 U394 ( .A1(n355), .A2(n412), .ZN(n354) );
  XNOR2_X1 U395 ( .A(n445), .B(KEYINPUT71), .ZN(n371) );
  BUF_X1 U396 ( .A(n512), .Z(n644) );
  NAND2_X1 U397 ( .A1(n349), .A2(n348), .ZN(n598) );
  AND2_X1 U398 ( .A1(n603), .A2(G953), .ZN(n707) );
  XNOR2_X1 U399 ( .A(n508), .B(n507), .ZN(n511) );
  INV_X1 U400 ( .A(KEYINPUT32), .ZN(n507) );
  XNOR2_X1 U401 ( .A(n371), .B(n713), .ZN(n438) );
  XNOR2_X1 U402 ( .A(n557), .B(KEYINPUT1), .ZN(n512) );
  AND2_X1 U403 ( .A1(n592), .A2(n589), .ZN(n347) );
  OR2_X1 U404 ( .A1(n587), .A2(n586), .ZN(n348) );
  NAND2_X1 U405 ( .A1(n352), .A2(n350), .ZN(n349) );
  INV_X1 U406 ( .A(n594), .ZN(n351) );
  INV_X1 U407 ( .A(n444), .ZN(n355) );
  NAND2_X1 U408 ( .A1(n444), .A2(G902), .ZN(n357) );
  NAND2_X1 U409 ( .A1(n599), .A2(n444), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n443), .B(n454), .ZN(n599) );
  NAND2_X2 U411 ( .A1(n361), .A2(n359), .ZN(n367) );
  INV_X1 U412 ( .A(n679), .ZN(n360) );
  NAND2_X1 U413 ( .A1(n679), .A2(n363), .ZN(n362) );
  INV_X1 U414 ( .A(n531), .ZN(n366) );
  XNOR2_X2 U415 ( .A(n367), .B(n521), .ZN(n614) );
  XNOR2_X1 U416 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U417 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U418 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n457) );
  XNOR2_X1 U419 ( .A(n398), .B(n397), .ZN(n516) );
  XNOR2_X1 U420 ( .A(n386), .B(n385), .ZN(n487) );
  NOR2_X1 U421 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U422 ( .A(n435), .B(n434), .ZN(n539) );
  XNOR2_X2 U423 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n368) );
  XNOR2_X1 U424 ( .A(G107), .B(G104), .ZN(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT90), .B(G110), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n713) );
  XNOR2_X1 U427 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n373) );
  XNOR2_X1 U428 ( .A(KEYINPUT18), .B(KEYINPUT79), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n376) );
  NAND2_X1 U430 ( .A1(n723), .A2(G224), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n374), .B(KEYINPUT78), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X2 U433 ( .A(G143), .B(G128), .ZN(n409) );
  XNOR2_X1 U434 ( .A(G146), .B(G125), .ZN(n416) );
  XNOR2_X1 U435 ( .A(n409), .B(n416), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n382) );
  XNOR2_X1 U437 ( .A(G116), .B(G113), .ZN(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT3), .B(G119), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n446) );
  XNOR2_X1 U440 ( .A(KEYINPUT16), .B(G122), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n446), .B(n381), .ZN(n715) );
  XNOR2_X1 U442 ( .A(n382), .B(n715), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n438), .B(n383), .ZN(n686) );
  XNOR2_X1 U444 ( .A(KEYINPUT15), .B(G902), .ZN(n587) );
  NAND2_X1 U445 ( .A1(n686), .A2(n587), .ZN(n386) );
  INV_X1 U446 ( .A(G902), .ZN(n412) );
  INV_X1 U447 ( .A(G237), .ZN(n384) );
  NAND2_X1 U448 ( .A1(n412), .A2(n384), .ZN(n387) );
  NAND2_X1 U449 ( .A1(n387), .A2(G210), .ZN(n385) );
  INV_X1 U450 ( .A(n487), .ZN(n389) );
  AND2_X1 U451 ( .A1(n387), .A2(G214), .ZN(n489) );
  INV_X1 U452 ( .A(n489), .ZN(n388) );
  NAND2_X1 U453 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n390), .B(KEYINPUT19), .ZN(n566) );
  XOR2_X1 U455 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n392) );
  NAND2_X1 U456 ( .A1(G234), .A2(G237), .ZN(n391) );
  XNOR2_X1 U457 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U458 ( .A(KEYINPUT74), .B(n393), .ZN(n394) );
  NAND2_X1 U459 ( .A1(G952), .A2(n394), .ZN(n676) );
  OR2_X1 U460 ( .A1(n676), .A2(G953), .ZN(n480) );
  NAND2_X1 U461 ( .A1(G902), .A2(n394), .ZN(n476) );
  INV_X1 U462 ( .A(G898), .ZN(n710) );
  NAND2_X1 U463 ( .A1(G953), .A2(n710), .ZN(n717) );
  OR2_X1 U464 ( .A1(n476), .A2(n717), .ZN(n395) );
  NAND2_X1 U465 ( .A1(n480), .A2(n395), .ZN(n396) );
  NAND2_X1 U466 ( .A1(n566), .A2(n396), .ZN(n398) );
  XNOR2_X1 U467 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n397) );
  XOR2_X1 U468 ( .A(KEYINPUT7), .B(KEYINPUT104), .Z(n400) );
  XNOR2_X1 U469 ( .A(G116), .B(G122), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U471 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n402) );
  XNOR2_X1 U472 ( .A(G107), .B(KEYINPUT103), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U474 ( .A(n404), .B(n403), .Z(n408) );
  XOR2_X1 U475 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n406) );
  NAND2_X1 U476 ( .A1(G234), .A2(n723), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n459) );
  NAND2_X1 U478 ( .A1(G217), .A2(n459), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n408), .B(n407), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n409), .B(G134), .ZN(n442) );
  INV_X1 U481 ( .A(n442), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n701) );
  NAND2_X1 U483 ( .A1(n701), .A2(n412), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n413), .B(G478), .ZN(n501) );
  INV_X1 U485 ( .A(KEYINPUT10), .ZN(n414) );
  XNOR2_X1 U486 ( .A(n414), .B(G140), .ZN(n415) );
  XNOR2_X1 U487 ( .A(n416), .B(n415), .ZN(n721) );
  XOR2_X1 U488 ( .A(KEYINPUT11), .B(G122), .Z(n418) );
  XNOR2_X1 U489 ( .A(G143), .B(G113), .ZN(n417) );
  XNOR2_X1 U490 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n721), .B(n419), .ZN(n426) );
  XOR2_X1 U492 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n421) );
  NOR2_X1 U493 ( .A1(G953), .A2(G237), .ZN(n447) );
  NAND2_X1 U494 ( .A1(G214), .A2(n447), .ZN(n420) );
  XNOR2_X1 U495 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U496 ( .A(G104), .B(n422), .ZN(n424) );
  INV_X1 U497 ( .A(n440), .ZN(n423) );
  XOR2_X1 U498 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U499 ( .A(n426), .B(n425), .ZN(n693) );
  NOR2_X1 U500 ( .A1(G902), .A2(n693), .ZN(n428) );
  XNOR2_X1 U501 ( .A(KEYINPUT13), .B(G475), .ZN(n427) );
  XNOR2_X1 U502 ( .A(n428), .B(n427), .ZN(n500) );
  OR2_X1 U503 ( .A1(n501), .A2(n500), .ZN(n664) );
  NAND2_X1 U504 ( .A1(n587), .A2(G234), .ZN(n429) );
  XNOR2_X1 U505 ( .A(n429), .B(KEYINPUT20), .ZN(n467) );
  NAND2_X1 U506 ( .A1(n467), .A2(G221), .ZN(n432) );
  XOR2_X1 U507 ( .A(KEYINPUT97), .B(KEYINPUT21), .Z(n430) );
  XNOR2_X1 U508 ( .A(n430), .B(KEYINPUT96), .ZN(n431) );
  XNOR2_X1 U509 ( .A(n432), .B(n431), .ZN(n646) );
  NOR2_X1 U510 ( .A1(n664), .A2(n646), .ZN(n433) );
  NAND2_X1 U511 ( .A1(n516), .A2(n433), .ZN(n435) );
  XOR2_X1 U512 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n434) );
  NAND2_X1 U513 ( .A1(G227), .A2(n723), .ZN(n436) );
  XNOR2_X1 U514 ( .A(G140), .B(n436), .ZN(n437) );
  XNOR2_X1 U515 ( .A(n438), .B(n437), .ZN(n443) );
  XNOR2_X1 U516 ( .A(KEYINPUT4), .B(G137), .ZN(n439) );
  XNOR2_X1 U517 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U518 ( .A(n442), .B(n441), .ZN(n720) );
  XNOR2_X1 U519 ( .A(n720), .B(G146), .ZN(n454) );
  XOR2_X1 U520 ( .A(KEYINPUT70), .B(G469), .Z(n444) );
  XNOR2_X1 U521 ( .A(n445), .B(n446), .ZN(n452) );
  NAND2_X1 U522 ( .A1(n447), .A2(G210), .ZN(n448) );
  XNOR2_X1 U523 ( .A(n448), .B(KEYINPUT76), .ZN(n450) );
  XNOR2_X1 U524 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n449) );
  XNOR2_X1 U525 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U526 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U527 ( .A(n454), .B(n453), .ZN(n608) );
  XNOR2_X1 U528 ( .A(G472), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X2 U529 ( .A(n456), .B(n455), .ZN(n652) );
  INV_X1 U530 ( .A(n652), .ZN(n525) );
  XNOR2_X1 U531 ( .A(n457), .B(KEYINPUT23), .ZN(n458) );
  XOR2_X1 U532 ( .A(KEYINPUT93), .B(n458), .Z(n461) );
  NAND2_X1 U533 ( .A1(G221), .A2(n459), .ZN(n460) );
  XNOR2_X1 U534 ( .A(n461), .B(n460), .ZN(n466) );
  XOR2_X1 U535 ( .A(G110), .B(G119), .Z(n463) );
  XNOR2_X1 U536 ( .A(G137), .B(G128), .ZN(n462) );
  XNOR2_X1 U537 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U538 ( .A(n721), .B(n464), .ZN(n465) );
  XNOR2_X1 U539 ( .A(n466), .B(n465), .ZN(n704) );
  NOR2_X1 U540 ( .A1(G902), .A2(n704), .ZN(n472) );
  NAND2_X1 U541 ( .A1(n467), .A2(G217), .ZN(n470) );
  XNOR2_X1 U542 ( .A(KEYINPUT94), .B(KEYINPUT25), .ZN(n468) );
  XOR2_X1 U543 ( .A(n468), .B(KEYINPUT95), .Z(n469) );
  INV_X1 U544 ( .A(n493), .ZN(n473) );
  INV_X1 U545 ( .A(n473), .ZN(n535) );
  NOR2_X1 U546 ( .A1(n525), .A2(n535), .ZN(n474) );
  NAND2_X1 U547 ( .A1(n644), .A2(n474), .ZN(n475) );
  NOR2_X1 U548 ( .A1(n539), .A2(n475), .ZN(n510) );
  XOR2_X1 U549 ( .A(G110), .B(n510), .Z(G12) );
  XNOR2_X1 U550 ( .A(n652), .B(KEYINPUT6), .ZN(n536) );
  INV_X1 U551 ( .A(n501), .ZN(n519) );
  NAND2_X1 U552 ( .A1(n519), .A2(n500), .ZN(n631) );
  NOR2_X1 U553 ( .A1(G900), .A2(n476), .ZN(n477) );
  NAND2_X1 U554 ( .A1(G953), .A2(n477), .ZN(n479) );
  INV_X1 U555 ( .A(KEYINPUT111), .ZN(n478) );
  XNOR2_X1 U556 ( .A(n479), .B(n478), .ZN(n481) );
  AND2_X1 U557 ( .A1(n481), .A2(n480), .ZN(n494) );
  NOR2_X1 U558 ( .A1(n493), .A2(n494), .ZN(n552) );
  NAND2_X1 U559 ( .A1(n388), .A2(n552), .ZN(n482) );
  OR2_X1 U560 ( .A1(n646), .A2(n482), .ZN(n483) );
  NOR2_X1 U561 ( .A1(n631), .A2(n483), .ZN(n484) );
  NAND2_X1 U562 ( .A1(n536), .A2(n484), .ZN(n576) );
  XOR2_X1 U563 ( .A(KEYINPUT112), .B(n576), .Z(n485) );
  NAND2_X1 U564 ( .A1(n485), .A2(n644), .ZN(n486) );
  XNOR2_X1 U565 ( .A(n486), .B(KEYINPUT43), .ZN(n488) );
  BUF_X1 U566 ( .A(n487), .Z(n575) );
  NAND2_X1 U567 ( .A1(n488), .A2(n575), .ZN(n592) );
  XNOR2_X1 U568 ( .A(n592), .B(G140), .ZN(G42) );
  INV_X1 U569 ( .A(KEYINPUT30), .ZN(n490) );
  XNOR2_X1 U570 ( .A(n491), .B(n490), .ZN(n496) );
  INV_X1 U571 ( .A(n646), .ZN(n492) );
  NAND2_X1 U572 ( .A1(n493), .A2(n492), .ZN(n643) );
  OR2_X1 U573 ( .A1(n643), .A2(n557), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n526), .A2(n494), .ZN(n495) );
  AND2_X1 U575 ( .A1(n496), .A2(n495), .ZN(n497) );
  XNOR2_X1 U576 ( .A(n497), .B(KEYINPUT77), .ZN(n571) );
  XNOR2_X1 U577 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n498) );
  XNOR2_X1 U578 ( .A(n575), .B(n498), .ZN(n550) );
  XNOR2_X1 U579 ( .A(n499), .B(KEYINPUT39), .ZN(n561) );
  INV_X1 U580 ( .A(n500), .ZN(n518) );
  NAND2_X1 U581 ( .A1(n518), .A2(n501), .ZN(n502) );
  XNOR2_X1 U582 ( .A(n502), .B(KEYINPUT105), .ZN(n623) );
  NAND2_X1 U583 ( .A1(n561), .A2(n623), .ZN(n589) );
  XNOR2_X1 U584 ( .A(n589), .B(G134), .ZN(G36) );
  INV_X1 U585 ( .A(n539), .ZN(n506) );
  NOR2_X1 U586 ( .A1(n644), .A2(n535), .ZN(n503) );
  XOR2_X1 U587 ( .A(KEYINPUT108), .B(n503), .Z(n504) );
  NOR2_X1 U588 ( .A1(n504), .A2(n536), .ZN(n505) );
  NAND2_X1 U589 ( .A1(n506), .A2(n505), .ZN(n508) );
  XOR2_X1 U590 ( .A(G119), .B(KEYINPUT126), .Z(n509) );
  XNOR2_X1 U591 ( .A(n511), .B(n509), .ZN(G21) );
  NOR2_X1 U592 ( .A1(n511), .A2(n510), .ZN(n522) );
  OR2_X2 U593 ( .A1(n512), .A2(n643), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(KEYINPUT109), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n513), .A2(n536), .ZN(n515) );
  XNOR2_X1 U596 ( .A(KEYINPUT110), .B(KEYINPUT33), .ZN(n514) );
  INV_X1 U597 ( .A(KEYINPUT34), .ZN(n517) );
  OR2_X1 U598 ( .A1(n519), .A2(n518), .ZN(n572) );
  INV_X1 U599 ( .A(n572), .ZN(n520) );
  XNOR2_X1 U600 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n521) );
  NAND2_X1 U601 ( .A1(n522), .A2(n614), .ZN(n524) );
  INV_X1 U602 ( .A(KEYINPUT44), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n541), .A2(KEYINPUT72), .ZN(n523) );
  XNOR2_X1 U604 ( .A(n524), .B(n523), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U606 ( .A1(n531), .A2(n527), .ZN(n528) );
  XNOR2_X1 U607 ( .A(KEYINPUT100), .B(n528), .ZN(n618) );
  NOR2_X1 U608 ( .A1(n529), .A2(n652), .ZN(n530) );
  NAND2_X1 U609 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U610 ( .A(KEYINPUT31), .B(n532), .Z(n633) );
  NAND2_X1 U611 ( .A1(n618), .A2(n633), .ZN(n533) );
  INV_X1 U612 ( .A(n631), .ZN(n629) );
  OR2_X1 U613 ( .A1(n623), .A2(n629), .ZN(n665) );
  NAND2_X1 U614 ( .A1(n533), .A2(n665), .ZN(n534) );
  XNOR2_X1 U615 ( .A(n534), .B(KEYINPUT106), .ZN(n544) );
  NOR2_X1 U616 ( .A1(n536), .A2(n473), .ZN(n537) );
  NAND2_X1 U617 ( .A1(n537), .A2(n644), .ZN(n538) );
  NOR2_X1 U618 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U619 ( .A(KEYINPUT107), .B(n540), .Z(n730) );
  NOR2_X1 U620 ( .A1(n541), .A2(KEYINPUT72), .ZN(n542) );
  NOR2_X1 U621 ( .A1(n730), .A2(n542), .ZN(n543) );
  NAND2_X1 U622 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U623 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U624 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n547) );
  XNOR2_X1 U625 ( .A(n548), .B(n547), .ZN(n588) );
  NOR2_X1 U626 ( .A1(n588), .A2(n587), .ZN(n549) );
  INV_X1 U627 ( .A(n550), .ZN(n662) );
  NAND2_X1 U628 ( .A1(n662), .A2(n388), .ZN(n666) );
  NOR2_X1 U629 ( .A1(n664), .A2(n666), .ZN(n551) );
  XNOR2_X1 U630 ( .A(KEYINPUT41), .B(n551), .ZN(n678) );
  INV_X1 U631 ( .A(n552), .ZN(n553) );
  OR2_X1 U632 ( .A1(n646), .A2(n553), .ZN(n554) );
  XOR2_X1 U633 ( .A(KEYINPUT28), .B(KEYINPUT113), .Z(n555) );
  XNOR2_X1 U634 ( .A(n556), .B(n555), .ZN(n558) );
  OR2_X1 U635 ( .A1(n558), .A2(n557), .ZN(n568) );
  OR2_X1 U636 ( .A1(n678), .A2(n568), .ZN(n560) );
  INV_X1 U637 ( .A(KEYINPUT42), .ZN(n559) );
  XNOR2_X1 U638 ( .A(n560), .B(n559), .ZN(n731) );
  NAND2_X1 U639 ( .A1(n561), .A2(n629), .ZN(n564) );
  INV_X1 U640 ( .A(KEYINPUT114), .ZN(n562) );
  XNOR2_X1 U641 ( .A(n562), .B(KEYINPUT40), .ZN(n563) );
  XNOR2_X1 U642 ( .A(n564), .B(n563), .ZN(n606) );
  XNOR2_X1 U643 ( .A(n565), .B(KEYINPUT46), .ZN(n583) );
  INV_X1 U644 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U645 ( .A(n569), .B(KEYINPUT80), .ZN(n628) );
  NAND2_X1 U646 ( .A1(n628), .A2(n665), .ZN(n570) );
  XNOR2_X1 U647 ( .A(n570), .B(KEYINPUT47), .ZN(n581) );
  INV_X1 U648 ( .A(n571), .ZN(n574) );
  NOR2_X1 U649 ( .A1(n572), .A2(n575), .ZN(n573) );
  AND2_X1 U650 ( .A1(n574), .A2(n573), .ZN(n627) );
  XNOR2_X1 U651 ( .A(n627), .B(KEYINPUT83), .ZN(n579) );
  OR2_X1 U652 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n577), .B(KEYINPUT36), .ZN(n578) );
  OR2_X1 U654 ( .A1(n578), .A2(n644), .ZN(n637) );
  NAND2_X1 U655 ( .A1(n579), .A2(n637), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U657 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n585), .B(n584), .ZN(n594) );
  INV_X1 U659 ( .A(KEYINPUT2), .ZN(n586) );
  BUF_X1 U660 ( .A(n588), .Z(n638) );
  INV_X1 U661 ( .A(n638), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n589), .A2(KEYINPUT2), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT81), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  AND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n641) );
  INV_X1 U667 ( .A(n641), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n703), .A2(G469), .ZN(n602) );
  XOR2_X1 U669 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n600) );
  XNOR2_X1 U670 ( .A(n599), .B(n600), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n602), .B(n601), .ZN(n604) );
  INV_X1 U672 ( .A(G952), .ZN(n603) );
  NOR2_X2 U673 ( .A1(n604), .A2(n707), .ZN(n605) );
  XNOR2_X1 U674 ( .A(n605), .B(KEYINPUT124), .ZN(G54) );
  XOR2_X1 U675 ( .A(G131), .B(n606), .Z(G33) );
  NAND2_X1 U676 ( .A1(n703), .A2(G472), .ZN(n610) );
  XOR2_X1 U677 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X2 U680 ( .A1(n611), .A2(n707), .ZN(n613) );
  XNOR2_X1 U681 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n613), .B(n612), .ZN(G57) );
  XNOR2_X1 U683 ( .A(n614), .B(G122), .ZN(G24) );
  NOR2_X1 U684 ( .A1(n618), .A2(n631), .ZN(n615) );
  XOR2_X1 U685 ( .A(G104), .B(n615), .Z(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT118), .B(KEYINPUT27), .Z(n617) );
  XNOR2_X1 U687 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n622) );
  INV_X1 U689 ( .A(n623), .ZN(n634) );
  NOR2_X1 U690 ( .A1(n618), .A2(n634), .ZN(n620) );
  XNOR2_X1 U691 ( .A(G107), .B(KEYINPUT26), .ZN(n619) );
  XNOR2_X1 U692 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(G9) );
  XOR2_X1 U694 ( .A(KEYINPUT119), .B(KEYINPUT29), .Z(n625) );
  NAND2_X1 U695 ( .A1(n623), .A2(n628), .ZN(n624) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  XOR2_X1 U697 ( .A(G128), .B(n626), .Z(G30) );
  XOR2_X1 U698 ( .A(G143), .B(n627), .Z(G45) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U700 ( .A(G146), .B(n630), .ZN(G48) );
  NOR2_X1 U701 ( .A1(n631), .A2(n633), .ZN(n632) );
  XOR2_X1 U702 ( .A(G113), .B(n632), .Z(G15) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U704 ( .A(G116), .B(n635), .Z(G18) );
  XOR2_X1 U705 ( .A(G125), .B(KEYINPUT37), .Z(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(G27) );
  NOR2_X1 U707 ( .A1(n638), .A2(n722), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n639), .A2(KEYINPUT2), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(KEYINPUT82), .ZN(n642) );
  NOR2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n684) );
  XNOR2_X1 U711 ( .A(KEYINPUT51), .B(KEYINPUT122), .ZN(n660) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U713 ( .A(KEYINPUT50), .B(n645), .ZN(n650) );
  XOR2_X1 U714 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n648) );
  NAND2_X1 U715 ( .A1(n646), .A2(n473), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n656) );
  OR2_X1 U718 ( .A1(n656), .A2(KEYINPUT121), .ZN(n651) );
  NAND2_X1 U719 ( .A1(n651), .A2(n652), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n652), .A2(KEYINPUT121), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n529), .A2(n653), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n656), .A2(KEYINPUT121), .ZN(n657) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U726 ( .A1(n661), .A2(n678), .ZN(n673) );
  NOR2_X1 U727 ( .A1(n662), .A2(n388), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n664), .A2(n663), .ZN(n670) );
  INV_X1 U729 ( .A(n665), .ZN(n667) );
  NOR2_X1 U730 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U731 ( .A(KEYINPUT123), .B(n668), .Z(n669) );
  NOR2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n671), .A2(n360), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n674), .B(KEYINPUT52), .ZN(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U737 ( .A1(n677), .A2(G953), .ZN(n682) );
  INV_X1 U738 ( .A(n678), .ZN(n680) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U741 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n685), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U743 ( .A1(n703), .A2(G210), .ZN(n690) );
  XOR2_X1 U744 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n687) );
  XNOR2_X1 U745 ( .A(n687), .B(KEYINPUT87), .ZN(n688) );
  XNOR2_X1 U746 ( .A(n686), .B(n688), .ZN(n689) );
  XNOR2_X1 U747 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X2 U748 ( .A1(n691), .A2(n707), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n692), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U750 ( .A1(n703), .A2(G475), .ZN(n697) );
  XNOR2_X1 U751 ( .A(KEYINPUT125), .B(KEYINPUT88), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n693), .B(KEYINPUT59), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U754 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X2 U755 ( .A1(n698), .A2(n707), .ZN(n699) );
  XNOR2_X1 U756 ( .A(n699), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U757 ( .A1(n703), .A2(G478), .ZN(n700) );
  XOR2_X1 U758 ( .A(n701), .B(n700), .Z(n702) );
  NOR2_X1 U759 ( .A1(n707), .A2(n702), .ZN(G63) );
  NAND2_X1 U760 ( .A1(n703), .A2(G217), .ZN(n705) );
  XNOR2_X1 U761 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n707), .A2(n706), .ZN(G66) );
  NOR2_X1 U763 ( .A1(n638), .A2(G953), .ZN(n712) );
  NAND2_X1 U764 ( .A1(G953), .A2(G224), .ZN(n708) );
  XOR2_X1 U765 ( .A(KEYINPUT61), .B(n708), .Z(n709) );
  NOR2_X1 U766 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n719) );
  XOR2_X1 U768 ( .A(G101), .B(n713), .Z(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U770 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U771 ( .A(n719), .B(n718), .ZN(G69) );
  XOR2_X1 U772 ( .A(n720), .B(n721), .Z(n725) );
  XNOR2_X1 U773 ( .A(n722), .B(n725), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n729) );
  XNOR2_X1 U775 ( .A(n725), .B(G227), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U779 ( .A(n730), .B(G101), .Z(G3) );
  XNOR2_X1 U780 ( .A(G137), .B(KEYINPUT127), .ZN(n732) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G39) );
endmodule

