//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927;
  INV_X1    g000(.A(KEYINPUT24), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(G183gat), .A3(G190gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G183gat), .B(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(new_n202), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT23), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT25), .ZN(new_n212));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(KEYINPUT23), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n205), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n208), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n211), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n212), .B1(new_n205), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n216), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT66), .B(new_n212), .C1(new_n205), .C2(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(KEYINPUT68), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n228), .A2(KEYINPUT26), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n206), .B1(new_n228), .B2(KEYINPUT26), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n231), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G183gat), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G190gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(G190gat), .B1(new_n234), .B2(KEYINPUT67), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n240), .B1(new_n244), .B2(KEYINPUT28), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n226), .A2(new_n227), .B1(new_n232), .B2(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(G113gat), .A2(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(G113gat), .A2(G120gat), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G127gat), .A2(G134gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g051(.A1(G127gat), .A2(G134gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT70), .B1(new_n255), .B2(new_n250), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT71), .B(KEYINPUT1), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n249), .A2(new_n254), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n253), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n255), .B2(new_n250), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n247), .A2(new_n248), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n261), .C1(KEYINPUT1), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT72), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n246), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n270), .B(KEYINPUT64), .Z(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT34), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n273), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n281), .B2(KEYINPUT33), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT32), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n282), .A2(new_n284), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n276), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n282), .A2(new_n284), .ZN(new_n289));
  INV_X1    g088(.A(new_n276), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT79), .B(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT2), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(G155gat), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n299), .A2(new_n300), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n299), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n300), .A2(new_n302), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n296), .A2(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n263), .A3(new_n258), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT4), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n265), .A2(new_n309), .A3(new_n267), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n316));
  OAI21_X1  g115(.A(G162gat), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n304), .B1(new_n317), .B2(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT3), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  INV_X1    g121(.A(new_n296), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n322), .B(new_n319), .C1(new_n323), .C2(new_n304), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n324), .A3(new_n264), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n265), .A2(KEYINPUT4), .A3(new_n309), .A4(new_n267), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n310), .A2(new_n311), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n327), .A3(new_n325), .A4(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n319), .B1(new_n323), .B2(new_n304), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n264), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n310), .ZN(new_n334));
  INV_X1    g133(.A(new_n327), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n314), .A2(new_n328), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  AOI21_X1  g140(.A(KEYINPUT6), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(new_n341), .B2(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n314), .A2(new_n328), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n331), .A2(new_n336), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n341), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n224), .A2(new_n225), .ZN(new_n351));
  INV_X1    g150(.A(new_n216), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n227), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n232), .A2(new_n245), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT29), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G226gat), .A2(G233gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT74), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT75), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n359));
  INV_X1    g158(.A(new_n357), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n359), .B(new_n360), .C1(new_n246), .C2(KEYINPUT29), .ZN(new_n361));
  INV_X1    g160(.A(G211gat), .ZN(new_n362));
  INV_X1    g161(.A(G218gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G197gat), .ZN(new_n365));
  INV_X1    g164(.A(G204gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368));
  OAI22_X1  g167(.A1(KEYINPUT22), .A2(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G211gat), .B(G218gat), .Z(new_n370));
  OR2_X1    g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(KEYINPUT73), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n353), .A2(new_n354), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n357), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n361), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT76), .ZN(new_n380));
  XOR2_X1   g179(.A(G8gat), .B(G36gat), .Z(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT77), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n357), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n357), .B2(new_n355), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n376), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n358), .A2(new_n389), .A3(new_n361), .A4(new_n378), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n380), .A2(new_n385), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT30), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT30), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT78), .A3(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n379), .A2(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n388), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n384), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n309), .B1(new_n404), .B2(new_n322), .ZN(new_n405));
  INV_X1    g204(.A(new_n376), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n309), .B2(new_n322), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(G228gat), .B(G233gat), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n371), .B2(new_n373), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n332), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n411), .B(new_n412), .C1(new_n406), .C2(new_n407), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT31), .B(G50gat), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n409), .B2(new_n413), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n403), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n402), .A3(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n293), .A2(new_n350), .A3(new_n400), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT81), .B1(new_n337), .B2(new_n341), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n346), .A2(new_n427), .A3(new_n347), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n342), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(new_n348), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT35), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n293), .A2(new_n400), .A3(new_n423), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT36), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n286), .A2(new_n287), .A3(new_n276), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n290), .B1(new_n289), .B2(new_n285), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n288), .A2(KEYINPUT36), .A3(new_n291), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n422), .B1(new_n399), .B2(new_n349), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n428), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n313), .A2(new_n311), .ZN(new_n445));
  INV_X1    g244(.A(new_n312), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n325), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n447), .B2(new_n335), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n444), .A3(new_n335), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n334), .A2(new_n335), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n447), .A2(new_n444), .A3(new_n335), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n452), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(new_n341), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT40), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT40), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n456), .A3(new_n459), .A4(new_n341), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n443), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n422), .B1(new_n399), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT82), .B(KEYINPUT38), .ZN(new_n463));
  XOR2_X1   g262(.A(KEYINPUT83), .B(KEYINPUT37), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n380), .A2(new_n388), .A3(new_n390), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT37), .B1(new_n396), .B2(new_n397), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n384), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n468), .A2(KEYINPUT85), .A3(new_n384), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n384), .A2(new_n463), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n476), .B1(new_n387), .B2(new_n406), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n358), .A2(new_n361), .A3(new_n376), .A4(new_n386), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n429), .A2(new_n391), .A3(new_n348), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n430), .A2(new_n480), .A3(KEYINPUT84), .A4(new_n391), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n462), .B1(new_n473), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT86), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n462), .B(KEYINPUT86), .C1(new_n473), .C2(new_n485), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n442), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n434), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(G29gat), .A2(G36gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT14), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G29gat), .ZN(new_n495));
  INV_X1    g294(.A(G36gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G43gat), .B(G50gat), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n498), .A2(KEYINPUT15), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT88), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT87), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n493), .A2(new_n504), .B1(new_n495), .B2(new_n496), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT90), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT89), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n515), .B(G8gat), .C1(KEYINPUT89), .C2(new_n509), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n507), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT13), .Z(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n507), .B(KEYINPUT17), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT18), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G113gat), .B(G141gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(new_n365), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT11), .B(G169gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT12), .Z(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n520), .A4(new_n526), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT91), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n529), .A2(new_n539), .A3(new_n535), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n529), .A2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n491), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT98), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554));
  AND2_X1   g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT99), .B(G85gat), .Z(new_n556));
  OAI221_X1 g355(.A(new_n553), .B1(new_n554), .B2(new_n555), .C1(G92gat), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G99gat), .B(G106gat), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT100), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT100), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n564), .A3(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n524), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n566), .A2(new_n507), .B1(KEYINPUT41), .B2(new_n546), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n239), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n239), .B1(new_n568), .B2(new_n569), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n363), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n572), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(G218gat), .A3(new_n570), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(new_n575), .A3(new_n576), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n549), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n549), .A3(new_n581), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G57gat), .B(G64gat), .Z(new_n586));
  INV_X1    g385(.A(G71gat), .ZN(new_n587));
  INV_X1    g386(.A(G78gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n586), .B1(KEYINPUT9), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G127gat), .B(G155gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT92), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n518), .B1(new_n594), .B2(new_n593), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT93), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n604));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n585), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G230gat), .ZN(new_n610));
  INV_X1    g409(.A(G233gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n562), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n615), .A2(new_n561), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n561), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n593), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n592), .B1(new_n563), .B2(new_n565), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n566), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n612), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n624), .B(new_n625), .Z(new_n626));
  INV_X1    g425(.A(new_n612), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n618), .A2(new_n619), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n623), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630));
  INV_X1    g429(.A(new_n626), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n628), .A2(new_n627), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(KEYINPUT102), .B(new_n631), .C1(new_n622), .C2(new_n632), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n609), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n545), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n349), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g440(.A1(new_n545), .A2(new_n399), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT16), .B(G8gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n648), .B1(new_n645), .B2(new_n512), .ZN(new_n649));
  MUX2_X1   g448(.A(new_n648), .B(new_n649), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g449(.A(G15gat), .B1(new_n639), .B2(new_n293), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT104), .ZN(new_n652));
  INV_X1    g451(.A(new_n440), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(G15gat), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n639), .B2(new_n654), .ZN(G1326gat));
  NOR2_X1   g454(.A1(new_n638), .A2(new_n423), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT43), .B(G22gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT105), .B(KEYINPUT106), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  NAND2_X1  g459(.A1(new_n488), .A2(new_n489), .ZN(new_n661));
  INV_X1    g460(.A(new_n442), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT107), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n664));
  AOI211_X1 g463(.A(new_n664), .B(new_n442), .C1(new_n488), .C2(new_n489), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n433), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n585), .A2(KEYINPUT44), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(KEYINPUT108), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n584), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n582), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n434), .B2(new_n490), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT44), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT108), .B1(new_n666), .B2(new_n667), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n636), .A2(new_n608), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n544), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(new_n349), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G29gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n491), .A2(new_n670), .A3(new_n678), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G29gat), .A3(new_n350), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1328gat));
  OAI211_X1 g483(.A(new_n399), .B(new_n678), .C1(new_n673), .C2(new_n674), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n496), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n686), .B2(new_n685), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n670), .A2(new_n676), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n643), .A2(new_n496), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1329gat));
  NOR3_X1   g494(.A1(new_n681), .A2(G43gat), .A3(new_n292), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n675), .A2(new_n653), .A3(new_n678), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G43gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g498(.A(new_n422), .B(new_n678), .C1(new_n673), .C2(new_n674), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G50gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n423), .A2(G50gat), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT113), .Z(new_n703));
  AND2_X1   g502(.A1(new_n689), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n545), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(KEYINPUT48), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n701), .A2(KEYINPUT112), .B1(new_n545), .B2(new_n704), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n700), .A2(new_n709), .A3(G50gat), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n707), .B(KEYINPUT48), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n701), .A2(KEYINPUT112), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n710), .A3(new_n705), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT114), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n706), .B1(new_n711), .B2(new_n715), .ZN(G1331gat));
  INV_X1    g515(.A(new_n666), .ZN(new_n717));
  INV_X1    g516(.A(new_n544), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n585), .A2(new_n718), .A3(new_n608), .A4(new_n636), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n717), .A2(KEYINPUT115), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT115), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n350), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n400), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n722), .B2(new_n440), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n293), .A2(new_n587), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n722), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g532(.A1(new_n722), .A2(new_n423), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(new_n588), .ZN(G1335gat));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n607), .ZN(new_n736));
  INV_X1    g535(.A(new_n636), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n675), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n349), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n556), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n717), .A2(new_n585), .A3(new_n736), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n636), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n350), .A2(new_n556), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(G1336gat));
  INV_X1    g545(.A(G92gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n737), .A2(new_n400), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n743), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n675), .A2(new_n399), .A3(new_n738), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g552(.A1(new_n744), .A2(G99gat), .A3(new_n292), .ZN(new_n754));
  INV_X1    g553(.A(G99gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n739), .B2(new_n653), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n754), .A2(new_n756), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n675), .A2(new_n422), .A3(new_n738), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G106gat), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n423), .A2(G106gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n744), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n519), .A2(new_n522), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT116), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n525), .A2(new_n526), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n520), .B2(new_n765), .ZN(new_n766));
  AOI22_X1  g565(.A1(new_n538), .A2(new_n540), .B1(new_n533), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n620), .A2(new_n612), .A3(new_n621), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT54), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n626), .B1(new_n622), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n769), .A2(KEYINPUT55), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n629), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT55), .B1(new_n769), .B2(new_n771), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n670), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n544), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n533), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n541), .A2(new_n635), .A3(new_n634), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n585), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n608), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n609), .A2(new_n544), .A3(new_n636), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n422), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n292), .A2(new_n399), .A3(new_n350), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n544), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n636), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n608), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g593(.A1(new_n787), .A2(new_n585), .ZN(new_n795));
  INV_X1    g594(.A(G134gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n797), .A2(KEYINPUT56), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n800), .A2(new_n801), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n798), .B(new_n799), .C1(new_n803), .C2(new_n804), .ZN(G1343gat));
  NOR3_X1   g604(.A1(new_n653), .A2(new_n350), .A3(new_n399), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n423), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n783), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n779), .A2(KEYINPUT118), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n636), .A2(new_n812), .A3(new_n767), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n813), .A3(new_n777), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n585), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n608), .B1(new_n815), .B2(new_n776), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n810), .B1(new_n816), .B2(KEYINPUT119), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n779), .A2(KEYINPUT118), .B1(new_n775), .B2(new_n544), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n670), .B1(new_n818), .B2(new_n813), .ZN(new_n819));
  AND4_X1   g618(.A1(new_n584), .A2(new_n583), .A3(new_n767), .A4(new_n775), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n607), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n809), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n808), .B1(new_n784), .B2(new_n423), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n807), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n297), .B1(new_n826), .B2(new_n544), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT120), .B1(new_n784), .B2(new_n350), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n349), .C1(new_n782), .C2(new_n783), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n653), .A2(new_n399), .A3(new_n423), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n832), .A2(G141gat), .A3(new_n718), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT58), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n809), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n783), .B1(new_n821), .B2(new_n822), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n782), .A2(new_n783), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT57), .B1(new_n839), .B2(new_n422), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n544), .B(new_n806), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT121), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n843), .A3(new_n544), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n842), .A2(new_n844), .A3(G141gat), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n833), .A2(KEYINPUT58), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(G1344gat));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n636), .A3(new_n830), .A4(new_n831), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT59), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n298), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n826), .A2(new_n851), .A3(new_n636), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n422), .B1(new_n816), .B2(new_n783), .ZN(new_n853));
  AOI22_X1  g652(.A1(new_n839), .A2(new_n809), .B1(new_n853), .B2(new_n808), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n806), .A2(new_n636), .ZN(new_n855));
  OAI211_X1 g654(.A(KEYINPUT59), .B(G148gat), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n850), .A2(new_n852), .A3(new_n856), .A4(KEYINPUT122), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1345gat));
  AOI21_X1  g660(.A(new_n294), .B1(new_n826), .B2(new_n608), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863));
  INV_X1    g662(.A(new_n294), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n832), .A2(new_n864), .A3(new_n607), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n863), .B1(new_n862), .B2(new_n865), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1346gat));
  AND2_X1   g667(.A1(new_n826), .A2(new_n670), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n670), .A2(new_n295), .ZN(new_n870));
  OAI22_X1  g669(.A1(new_n869), .A2(new_n295), .B1(new_n832), .B2(new_n870), .ZN(G1347gat));
  NOR3_X1   g670(.A1(new_n400), .A2(new_n292), .A3(new_n422), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n839), .A2(new_n350), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n874), .A2(new_n220), .A3(new_n221), .A4(new_n544), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT124), .Z(new_n876));
  NAND2_X1  g675(.A1(new_n399), .A2(new_n350), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n292), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n785), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879), .B2(new_n718), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(G1348gat));
  AOI21_X1  g680(.A(G176gat), .B1(new_n874), .B2(new_n636), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n785), .A2(G176gat), .A3(new_n636), .A4(new_n878), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT126), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n882), .A2(new_n883), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(G1349gat));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n608), .A2(new_n238), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n873), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n873), .B2(new_n891), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G183gat), .B1(new_n879), .B2(new_n607), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT60), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n239), .A3(new_n670), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n785), .A2(new_n670), .A3(new_n878), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(G190gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n902), .B2(G190gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(G1351gat));
  INV_X1    g706(.A(new_n854), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n653), .A2(new_n877), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(new_n365), .A3(new_n718), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n839), .A2(new_n350), .A3(new_n422), .A4(new_n440), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n400), .ZN(new_n913));
  AOI21_X1  g712(.A(G197gat), .B1(new_n913), .B2(new_n544), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n911), .A2(new_n914), .ZN(G1352gat));
  OAI21_X1  g714(.A(G204gat), .B1(new_n910), .B2(new_n737), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n748), .A2(new_n366), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT62), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OR3_X1    g717(.A1(new_n912), .A2(KEYINPUT62), .A3(new_n917), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(G1353gat));
  NAND3_X1  g719(.A1(new_n913), .A2(new_n362), .A3(new_n608), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n908), .A2(new_n608), .A3(new_n909), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n922), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT63), .B1(new_n922), .B2(G211gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n910), .B2(new_n585), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n913), .A2(new_n363), .A3(new_n670), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1355gat));
endmodule


