

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U551 ( .A1(n781), .A2(n795), .ZN(n520) );
  NOR2_X1 U552 ( .A1(n986), .A2(n688), .ZN(n690) );
  NAND2_X1 U553 ( .A1(n782), .A2(n520), .ZN(n783) );
  NOR2_X1 U554 ( .A1(n643), .A2(G651), .ZN(n638) );
  NAND2_X1 U555 ( .A1(G2104), .A2(G101), .ZN(n521) );
  NOR2_X1 U556 ( .A1(G2105), .A2(n521), .ZN(n522) );
  XNOR2_X1 U557 ( .A(KEYINPUT66), .B(n522), .ZN(n523) );
  XNOR2_X1 U558 ( .A(n523), .B(KEYINPUT23), .ZN(n527) );
  XNOR2_X1 U559 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n525) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U561 ( .A(n525), .B(n524), .ZN(n875) );
  NAND2_X1 U562 ( .A1(G137), .A2(n875), .ZN(n526) );
  NAND2_X1 U563 ( .A1(n527), .A2(n526), .ZN(n532) );
  INV_X1 U564 ( .A(G2104), .ZN(n546) );
  INV_X1 U565 ( .A(G2105), .ZN(n528) );
  NOR2_X1 U566 ( .A1(n546), .A2(n528), .ZN(n870) );
  NAND2_X1 U567 ( .A1(G113), .A2(n870), .ZN(n530) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n528), .ZN(n871) );
  NAND2_X1 U569 ( .A1(G125), .A2(n871), .ZN(n529) );
  NAND2_X1 U570 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U571 ( .A1(n532), .A2(n531), .ZN(n534) );
  INV_X1 U572 ( .A(KEYINPUT65), .ZN(n533) );
  XNOR2_X1 U573 ( .A(n534), .B(n533), .ZN(n680) );
  BUF_X1 U574 ( .A(n680), .Z(G160) );
  INV_X1 U575 ( .A(G651), .ZN(n538) );
  NOR2_X1 U576 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n535), .Z(n642) );
  NAND2_X1 U578 ( .A1(G64), .A2(n642), .ZN(n537) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n643) );
  NAND2_X1 U580 ( .A1(G52), .A2(n638), .ZN(n536) );
  NAND2_X1 U581 ( .A1(n537), .A2(n536), .ZN(n544) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n632) );
  NAND2_X1 U583 ( .A1(G90), .A2(n632), .ZN(n541) );
  OR2_X1 U584 ( .A1(n538), .A2(n643), .ZN(n539) );
  XOR2_X1 U585 ( .A(KEYINPUT68), .B(n539), .Z(n631) );
  NAND2_X1 U586 ( .A1(G77), .A2(n631), .ZN(n540) );
  NAND2_X1 U587 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U588 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U589 ( .A1(n544), .A2(n543), .ZN(G171) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U591 ( .A1(G135), .A2(n875), .ZN(n545) );
  XNOR2_X1 U592 ( .A(n545), .B(KEYINPUT74), .ZN(n553) );
  NOR2_X1 U593 ( .A1(G2105), .A2(n546), .ZN(n878) );
  NAND2_X1 U594 ( .A1(G99), .A2(n878), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G111), .A2(n870), .ZN(n547) );
  NAND2_X1 U596 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U597 ( .A1(n871), .A2(G123), .ZN(n549) );
  XOR2_X1 U598 ( .A(KEYINPUT18), .B(n549), .Z(n550) );
  NOR2_X1 U599 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n553), .A2(n552), .ZN(n917) );
  XNOR2_X1 U601 ( .A(G2096), .B(n917), .ZN(n554) );
  OR2_X1 U602 ( .A1(G2100), .A2(n554), .ZN(G156) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G132), .ZN(G219) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  NAND2_X1 U606 ( .A1(G88), .A2(n632), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G75), .A2(n631), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U609 ( .A1(G62), .A2(n642), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G50), .A2(n638), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U612 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U613 ( .A(KEYINPUT78), .B(n561), .Z(G303) );
  XOR2_X1 U614 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n563) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U616 ( .A(n563), .B(n562), .ZN(G223) );
  INV_X1 U617 ( .A(G223), .ZN(n823) );
  NAND2_X1 U618 ( .A1(n823), .A2(G567), .ZN(n564) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U620 ( .A1(n632), .A2(G81), .ZN(n565) );
  XNOR2_X1 U621 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G68), .A2(n631), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(n568), .ZN(n575) );
  XOR2_X1 U625 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n570) );
  NAND2_X1 U626 ( .A1(G56), .A2(n642), .ZN(n569) );
  XNOR2_X1 U627 ( .A(n570), .B(n569), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G43), .A2(n638), .ZN(n571) );
  XNOR2_X1 U629 ( .A(KEYINPUT73), .B(n571), .ZN(n572) );
  NOR2_X1 U630 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U631 ( .A1(n575), .A2(n574), .ZN(n986) );
  INV_X1 U632 ( .A(G860), .ZN(n605) );
  OR2_X1 U633 ( .A1(n986), .A2(n605), .ZN(G153) );
  INV_X1 U634 ( .A(G171), .ZN(G301) );
  NAND2_X1 U635 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U636 ( .A1(G92), .A2(n632), .ZN(n577) );
  NAND2_X1 U637 ( .A1(G79), .A2(n631), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G66), .A2(n642), .ZN(n579) );
  NAND2_X1 U640 ( .A1(G54), .A2(n638), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT15), .B(n582), .Z(n968) );
  OR2_X1 U644 ( .A1(n968), .A2(G868), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U646 ( .A1(n632), .A2(G89), .ZN(n585) );
  XNOR2_X1 U647 ( .A(n585), .B(KEYINPUT4), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G76), .A2(n631), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U650 ( .A(n588), .B(KEYINPUT5), .ZN(n593) );
  NAND2_X1 U651 ( .A1(G63), .A2(n642), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G51), .A2(n638), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT6), .B(n591), .Z(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U656 ( .A(n594), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U657 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U658 ( .A1(G91), .A2(n632), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G78), .A2(n631), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(KEYINPUT70), .B(n597), .Z(n601) );
  NAND2_X1 U662 ( .A1(G65), .A2(n642), .ZN(n599) );
  NAND2_X1 U663 ( .A1(G53), .A2(n638), .ZN(n598) );
  AND2_X1 U664 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U665 ( .A1(n601), .A2(n600), .ZN(G299) );
  INV_X1 U666 ( .A(G868), .ZN(n602) );
  NOR2_X1 U667 ( .A1(G286), .A2(n602), .ZN(n604) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U669 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n606), .A2(n968), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n986), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n968), .A2(G868), .ZN(n608) );
  NOR2_X1 U675 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U676 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U677 ( .A1(n968), .A2(G559), .ZN(n653) );
  XNOR2_X1 U678 ( .A(n986), .B(n653), .ZN(n611) );
  NOR2_X1 U679 ( .A1(G860), .A2(n611), .ZN(n613) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n613), .B(n612), .ZN(n620) );
  NAND2_X1 U682 ( .A1(G67), .A2(n642), .ZN(n615) );
  NAND2_X1 U683 ( .A1(G55), .A2(n638), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G93), .A2(n632), .ZN(n617) );
  NAND2_X1 U686 ( .A1(G80), .A2(n631), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n656) );
  XOR2_X1 U689 ( .A(n620), .B(n656), .Z(G145) );
  NAND2_X1 U690 ( .A1(G86), .A2(n632), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G61), .A2(n642), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n631), .A2(G73), .ZN(n623) );
  XNOR2_X1 U694 ( .A(n623), .B(KEYINPUT77), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT2), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n638), .A2(G48), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(G305) );
  NAND2_X1 U699 ( .A1(G60), .A2(n642), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G47), .A2(n638), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n636) );
  NAND2_X1 U702 ( .A1(G72), .A2(n631), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n632), .A2(G85), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT69), .ZN(G290) );
  NAND2_X1 U707 ( .A1(G49), .A2(n638), .ZN(n640) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U711 ( .A1(n643), .A2(G87), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n645), .A2(n644), .ZN(G288) );
  XNOR2_X1 U713 ( .A(n656), .B(G290), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n646), .B(G288), .ZN(n647) );
  XNOR2_X1 U715 ( .A(KEYINPUT19), .B(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n986), .B(KEYINPUT79), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(G305), .B(n650), .ZN(n652) );
  INV_X1 U719 ( .A(G299), .ZN(n978) );
  XNOR2_X1 U720 ( .A(n978), .B(G303), .ZN(n651) );
  XNOR2_X1 U721 ( .A(n652), .B(n651), .ZN(n896) );
  XNOR2_X1 U722 ( .A(KEYINPUT80), .B(n653), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n896), .B(n654), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(G868), .ZN(n658) );
  OR2_X1 U725 ( .A1(G868), .A2(n656), .ZN(n657) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U727 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U728 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U729 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U732 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U733 ( .A1(G220), .A2(G219), .ZN(n663) );
  XNOR2_X1 U734 ( .A(KEYINPUT22), .B(n663), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G96), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n665), .A2(G218), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT81), .ZN(n828) );
  NAND2_X1 U738 ( .A1(G2106), .A2(n828), .ZN(n670) );
  NAND2_X1 U739 ( .A1(G120), .A2(G108), .ZN(n667) );
  NOR2_X1 U740 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U741 ( .A1(G69), .A2(n668), .ZN(n827) );
  NAND2_X1 U742 ( .A1(G567), .A2(n827), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT82), .B(n671), .Z(G319) );
  INV_X1 U745 ( .A(G319), .ZN(n673) );
  NAND2_X1 U746 ( .A1(G661), .A2(G483), .ZN(n672) );
  NOR2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n826) );
  NAND2_X1 U748 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U749 ( .A1(G138), .A2(n875), .ZN(n675) );
  NAND2_X1 U750 ( .A1(G102), .A2(n878), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U752 ( .A1(G114), .A2(n870), .ZN(n677) );
  NAND2_X1 U753 ( .A1(G126), .A2(n871), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U755 ( .A1(n679), .A2(n678), .ZN(G164) );
  NOR2_X1 U756 ( .A1(G164), .A2(G1384), .ZN(n765) );
  AND2_X1 U757 ( .A1(n680), .A2(G40), .ZN(n763) );
  NAND2_X2 U758 ( .A1(n765), .A2(n763), .ZN(n723) );
  NAND2_X1 U759 ( .A1(G1961), .A2(n723), .ZN(n682) );
  INV_X1 U760 ( .A(n723), .ZN(n697) );
  XOR2_X1 U761 ( .A(G2078), .B(KEYINPUT25), .Z(n953) );
  NAND2_X1 U762 ( .A1(n697), .A2(n953), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n682), .A2(n681), .ZN(n710) );
  OR2_X1 U764 ( .A1(G301), .A2(n710), .ZN(n709) );
  INV_X1 U765 ( .A(n723), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G1996), .A2(n683), .ZN(n684) );
  XNOR2_X1 U767 ( .A(n684), .B(KEYINPUT26), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G1341), .A2(n723), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U770 ( .A(KEYINPUT91), .B(n687), .Z(n688) );
  NOR2_X1 U771 ( .A1(n690), .A2(n968), .ZN(n689) );
  XOR2_X1 U772 ( .A(n689), .B(KEYINPUT92), .Z(n696) );
  NAND2_X1 U773 ( .A1(n690), .A2(n968), .ZN(n694) );
  NOR2_X1 U774 ( .A1(n697), .A2(G1348), .ZN(n692) );
  NOR2_X1 U775 ( .A1(G2067), .A2(n723), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n702) );
  NAND2_X1 U779 ( .A1(n697), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U780 ( .A(n698), .B(KEYINPUT27), .ZN(n700) );
  AND2_X1 U781 ( .A1(G1956), .A2(n723), .ZN(n699) );
  NOR2_X1 U782 ( .A1(n700), .A2(n699), .ZN(n703) );
  NAND2_X1 U783 ( .A1(n978), .A2(n703), .ZN(n701) );
  NAND2_X1 U784 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U785 ( .A1(n978), .A2(n703), .ZN(n704) );
  XOR2_X1 U786 ( .A(n704), .B(KEYINPUT28), .Z(n705) );
  NAND2_X1 U787 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U788 ( .A(n707), .B(KEYINPUT29), .Z(n708) );
  NAND2_X1 U789 ( .A1(n709), .A2(n708), .ZN(n721) );
  NAND2_X1 U790 ( .A1(G301), .A2(n710), .ZN(n711) );
  XNOR2_X1 U791 ( .A(n711), .B(KEYINPUT95), .ZN(n718) );
  NAND2_X1 U792 ( .A1(G8), .A2(n723), .ZN(n795) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n795), .ZN(n734) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n723), .ZN(n731) );
  NOR2_X1 U795 ( .A1(n734), .A2(n731), .ZN(n712) );
  XOR2_X1 U796 ( .A(KEYINPUT93), .B(n712), .Z(n713) );
  NAND2_X1 U797 ( .A1(n713), .A2(G8), .ZN(n714) );
  XNOR2_X1 U798 ( .A(n714), .B(KEYINPUT30), .ZN(n715) );
  XNOR2_X1 U799 ( .A(KEYINPUT94), .B(n715), .ZN(n716) );
  NOR2_X1 U800 ( .A1(n716), .A2(G168), .ZN(n717) );
  NOR2_X1 U801 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U802 ( .A(KEYINPUT31), .B(n719), .Z(n720) );
  NAND2_X1 U803 ( .A1(n721), .A2(n720), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G286), .A2(n732), .ZN(n728) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n795), .ZN(n722) );
  XNOR2_X1 U806 ( .A(n722), .B(KEYINPUT96), .ZN(n725) );
  NOR2_X1 U807 ( .A1(n723), .A2(G2090), .ZN(n724) );
  NOR2_X1 U808 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U809 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U810 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U811 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U812 ( .A(n730), .B(KEYINPUT32), .ZN(n785) );
  NAND2_X1 U813 ( .A1(G8), .A2(n731), .ZN(n736) );
  INV_X1 U814 ( .A(n732), .ZN(n733) );
  NOR2_X1 U815 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U816 ( .A1(n736), .A2(n735), .ZN(n786) );
  INV_X1 U817 ( .A(n795), .ZN(n737) );
  NAND2_X1 U818 ( .A1(G1976), .A2(G288), .ZN(n972) );
  AND2_X1 U819 ( .A1(n737), .A2(n972), .ZN(n739) );
  AND2_X1 U820 ( .A1(n786), .A2(n739), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n785), .A2(n738), .ZN(n744) );
  INV_X1 U822 ( .A(n739), .ZN(n742) );
  NOR2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U824 ( .A1(G303), .A2(G1971), .ZN(n740) );
  NOR2_X1 U825 ( .A1(n971), .A2(n740), .ZN(n741) );
  OR2_X1 U826 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U828 ( .A(n745), .B(KEYINPUT64), .ZN(n746) );
  NOR2_X1 U829 ( .A1(KEYINPUT33), .A2(n746), .ZN(n784) );
  XOR2_X1 U830 ( .A(G1981), .B(G305), .Z(n964) );
  NAND2_X1 U831 ( .A1(G131), .A2(n875), .ZN(n748) );
  NAND2_X1 U832 ( .A1(G95), .A2(n878), .ZN(n747) );
  NAND2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G107), .A2(n870), .ZN(n750) );
  NAND2_X1 U835 ( .A1(G119), .A2(n871), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n751) );
  OR2_X1 U837 ( .A1(n752), .A2(n751), .ZN(n883) );
  NAND2_X1 U838 ( .A1(G1991), .A2(n883), .ZN(n753) );
  XOR2_X1 U839 ( .A(KEYINPUT87), .B(n753), .Z(n762) );
  NAND2_X1 U840 ( .A1(G141), .A2(n875), .ZN(n755) );
  NAND2_X1 U841 ( .A1(G117), .A2(n870), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n878), .A2(G105), .ZN(n756) );
  XOR2_X1 U844 ( .A(KEYINPUT38), .B(n756), .Z(n757) );
  NOR2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n760) );
  NAND2_X1 U846 ( .A1(n871), .A2(G129), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n866) );
  NAND2_X1 U848 ( .A1(G1996), .A2(n866), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n916) );
  INV_X1 U850 ( .A(n763), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n816) );
  NAND2_X1 U852 ( .A1(n916), .A2(n816), .ZN(n766) );
  XOR2_X1 U853 ( .A(KEYINPUT88), .B(n766), .Z(n807) );
  INV_X1 U854 ( .A(n807), .ZN(n780) );
  XOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .Z(n767) );
  XNOR2_X1 U856 ( .A(KEYINPUT83), .B(n767), .ZN(n814) );
  NAND2_X1 U857 ( .A1(G116), .A2(n870), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G128), .A2(n871), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n771) );
  XOR2_X1 U860 ( .A(KEYINPUT35), .B(KEYINPUT86), .Z(n770) );
  XNOR2_X1 U861 ( .A(n771), .B(n770), .ZN(n778) );
  XNOR2_X1 U862 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n772), .B(KEYINPUT34), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G140), .A2(n875), .ZN(n774) );
  NAND2_X1 U865 ( .A1(G104), .A2(n878), .ZN(n773) );
  NAND2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U867 ( .A(n776), .B(n775), .Z(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n779), .ZN(n890) );
  NOR2_X1 U870 ( .A1(n814), .A2(n890), .ZN(n936) );
  NAND2_X1 U871 ( .A1(n816), .A2(n936), .ZN(n811) );
  AND2_X1 U872 ( .A1(n780), .A2(n811), .ZN(n799) );
  AND2_X1 U873 ( .A1(n964), .A2(n799), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n971), .A2(KEYINPUT33), .ZN(n781) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n801) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n789) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n790), .A2(n795), .ZN(n797) );
  XNOR2_X1 U881 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n791), .B(KEYINPUT89), .ZN(n793) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XNOR2_X1 U884 ( .A(n793), .B(n792), .ZN(n794) );
  OR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n803) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U890 ( .A1(n982), .A2(n816), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n819) );
  XOR2_X1 U892 ( .A(KEYINPUT39), .B(KEYINPUT98), .Z(n804) );
  XNOR2_X1 U893 ( .A(KEYINPUT97), .B(n804), .ZN(n810) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n866), .ZN(n923) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n883), .ZN(n920) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n920), .A2(n805), .ZN(n806) );
  NOR2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n923), .A2(n808), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n810), .B(n809), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT99), .B(n813), .Z(n815) );
  NAND2_X1 U903 ( .A1(n814), .A2(n890), .ZN(n933) );
  NAND2_X1 U904 ( .A1(n815), .A2(n933), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n822) );
  XOR2_X1 U907 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n820) );
  XNOR2_X1 U908 ( .A(KEYINPUT40), .B(n820), .ZN(n821) );
  XNOR2_X1 U909 ( .A(n822), .B(n821), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U912 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n826), .A2(n825), .ZN(G188) );
  XNOR2_X1 U915 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  NOR2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U920 ( .A(G325), .ZN(G261) );
  XOR2_X1 U921 ( .A(G2474), .B(G1981), .Z(n830) );
  XNOR2_X1 U922 ( .A(G1966), .B(G1961), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U924 ( .A(n831), .B(KEYINPUT103), .Z(n833) );
  XNOR2_X1 U925 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U927 ( .A(G1976), .B(G1971), .Z(n835) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1956), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U930 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U931 ( .A(KEYINPUT104), .B(KEYINPUT41), .ZN(n838) );
  XNOR2_X1 U932 ( .A(n839), .B(n838), .ZN(G229) );
  XOR2_X1 U933 ( .A(G2100), .B(G2096), .Z(n841) );
  XNOR2_X1 U934 ( .A(KEYINPUT42), .B(G2678), .ZN(n840) );
  XNOR2_X1 U935 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2090), .Z(n843) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n842) );
  XNOR2_X1 U938 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U939 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U941 ( .A(n847), .B(n846), .ZN(G227) );
  NAND2_X1 U942 ( .A1(G124), .A2(n871), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT105), .B(n848), .Z(n849) );
  XNOR2_X1 U944 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U945 ( .A1(G136), .A2(n875), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U947 ( .A1(G100), .A2(n878), .ZN(n853) );
  NAND2_X1 U948 ( .A1(G112), .A2(n870), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U951 ( .A(KEYINPUT106), .B(n856), .ZN(G162) );
  NAND2_X1 U952 ( .A1(G118), .A2(n870), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G130), .A2(n871), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U955 ( .A1(n878), .A2(G106), .ZN(n859) );
  XOR2_X1 U956 ( .A(KEYINPUT107), .B(n859), .Z(n861) );
  NAND2_X1 U957 ( .A1(n875), .A2(G142), .ZN(n860) );
  NAND2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U959 ( .A(n862), .B(KEYINPUT45), .Z(n863) );
  NOR2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n865), .B(n917), .ZN(n869) );
  XNOR2_X1 U962 ( .A(G164), .B(n866), .ZN(n867) );
  XNOR2_X1 U963 ( .A(n867), .B(G162), .ZN(n868) );
  XOR2_X1 U964 ( .A(n869), .B(n868), .Z(n889) );
  NAND2_X1 U965 ( .A1(G115), .A2(n870), .ZN(n873) );
  NAND2_X1 U966 ( .A1(G127), .A2(n871), .ZN(n872) );
  NAND2_X1 U967 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U968 ( .A(n874), .B(KEYINPUT47), .ZN(n877) );
  NAND2_X1 U969 ( .A1(G139), .A2(n875), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G103), .A2(n878), .ZN(n879) );
  XNOR2_X1 U972 ( .A(KEYINPUT109), .B(n879), .ZN(n880) );
  NOR2_X1 U973 ( .A1(n881), .A2(n880), .ZN(n927) );
  XOR2_X1 U974 ( .A(KEYINPUT108), .B(KEYINPUT46), .Z(n882) );
  XNOR2_X1 U975 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U976 ( .A(n884), .B(KEYINPUT48), .Z(n886) );
  XNOR2_X1 U977 ( .A(G160), .B(KEYINPUT110), .ZN(n885) );
  XNOR2_X1 U978 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U979 ( .A(n927), .B(n887), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n889), .B(n888), .ZN(n891) );
  XNOR2_X1 U981 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U982 ( .A1(G37), .A2(n892), .ZN(G395) );
  XOR2_X1 U983 ( .A(KEYINPUT111), .B(G286), .Z(n894) );
  XNOR2_X1 U984 ( .A(G171), .B(n968), .ZN(n893) );
  XNOR2_X1 U985 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U986 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U987 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U988 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n899) );
  NOR2_X1 U989 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n911) );
  XOR2_X1 U991 ( .A(G2451), .B(G2443), .Z(n901) );
  XNOR2_X1 U992 ( .A(G2427), .B(G2454), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U994 ( .A(n902), .B(G2446), .Z(n904) );
  XNOR2_X1 U995 ( .A(G1348), .B(G1341), .ZN(n903) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U997 ( .A(G2435), .B(KEYINPUT102), .Z(n906) );
  XNOR2_X1 U998 ( .A(G2430), .B(G2438), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1000 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n909), .ZN(n914) );
  NAND2_X1 U1002 ( .A1(n914), .A2(G319), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G69), .ZN(G235) );
  INV_X1 U1008 ( .A(n914), .ZN(G401) );
  XNOR2_X1 U1009 ( .A(KEYINPUT52), .B(KEYINPUT115), .ZN(n938) );
  XOR2_X1 U1010 ( .A(G160), .B(G2084), .Z(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G2090), .B(KEYINPUT114), .Z(n921) );
  XNOR2_X1 U1015 ( .A(G162), .B(n921), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1017 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1019 ( .A(G2072), .B(n927), .Z(n929) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n928) );
  NOR2_X1 U1021 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1022 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1024 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1025 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(n938), .B(n937), .ZN(n939) );
  OR2_X1 U1027 ( .A1(KEYINPUT55), .A2(n939), .ZN(n940) );
  NAND2_X1 U1028 ( .A1(G29), .A2(n940), .ZN(n1024) );
  XOR2_X1 U1029 ( .A(G2084), .B(G34), .Z(n941) );
  XNOR2_X1 U1030 ( .A(KEYINPUT54), .B(n941), .ZN(n944) );
  XOR2_X1 U1031 ( .A(G2090), .B(KEYINPUT116), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G35), .B(n942), .ZN(n943) );
  NAND2_X1 U1033 ( .A1(n944), .A2(n943), .ZN(n959) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1035 ( .A(G1991), .B(G25), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1037 ( .A(G2072), .B(G33), .Z(n947) );
  NAND2_X1 U1038 ( .A1(n947), .A2(G28), .ZN(n950) );
  XOR2_X1 U1039 ( .A(KEYINPUT117), .B(G1996), .Z(n948) );
  XNOR2_X1 U1040 ( .A(G32), .B(n948), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G27), .B(n953), .ZN(n954) );
  NOR2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n956), .ZN(n957) );
  XNOR2_X1 U1046 ( .A(KEYINPUT118), .B(n957), .ZN(n958) );
  NOR2_X1 U1047 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1048 ( .A(KEYINPUT55), .B(n960), .Z(n961) );
  NOR2_X1 U1049 ( .A1(G29), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1050 ( .A(KEYINPUT119), .B(n962), .ZN(n963) );
  NAND2_X1 U1051 ( .A1(n963), .A2(G11), .ZN(n1022) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n966), .B(KEYINPUT120), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(KEYINPUT57), .B(n967), .ZN(n990) );
  XOR2_X1 U1057 ( .A(G1348), .B(n968), .Z(n970) );
  XOR2_X1 U1058 ( .A(G171), .B(G1961), .Z(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n985) );
  INV_X1 U1060 ( .A(n971), .ZN(n973) );
  NAND2_X1 U1061 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1062 ( .A(KEYINPUT121), .B(n974), .Z(n976) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G303), .ZN(n975) );
  NOR2_X1 U1064 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1065 ( .A(KEYINPUT122), .B(n977), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(n978), .B(G1956), .ZN(n979) );
  NAND2_X1 U1067 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1068 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1069 ( .A(KEYINPUT123), .B(n983), .Z(n984) );
  NAND2_X1 U1070 ( .A1(n985), .A2(n984), .ZN(n988) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n986), .ZN(n987) );
  NOR2_X1 U1072 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1073 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1074 ( .A1(n992), .A2(n991), .ZN(n1020) );
  INV_X1 U1075 ( .A(G16), .ZN(n1018) );
  XNOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(n993), .B(G4), .ZN(n997) );
  XNOR2_X1 U1078 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1079 ( .A(G1956), .B(G20), .ZN(n994) );
  NOR2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1082 ( .A(KEYINPUT125), .B(G1981), .Z(n998) );
  XNOR2_X1 U1083 ( .A(G6), .B(n998), .ZN(n999) );
  NOR2_X1 U1084 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(n1001), .B(KEYINPUT60), .ZN(n1004) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n1002) );
  XNOR2_X1 U1087 ( .A(KEYINPUT126), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1088 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1005), .B(KEYINPUT127), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G1961), .B(KEYINPUT124), .Z(n1006) );
  XNOR2_X1 U1091 ( .A(G5), .B(n1006), .ZN(n1007) );
  NAND2_X1 U1092 ( .A1(n1008), .A2(n1007), .ZN(n1015) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1102 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1103 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1104 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
  INV_X1 U1107 ( .A(G303), .ZN(G166) );
endmodule

