//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NOR2_X1   g0014(.A1(G58), .A2(G68), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n216), .A2(G50), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  OAI22_X1  g0021(.A1(new_n213), .A2(new_n214), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G116), .ZN(new_n224));
  INV_X1    g0024(.A(G270), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G97), .ZN(new_n230));
  INV_X1    g0030(.A(G257), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n226), .B(new_n232), .C1(G58), .C2(G232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n209), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT1), .Z(new_n235));
  AOI211_X1 g0035(.A(new_n222), .B(new_n235), .C1(new_n214), .C2(new_n213), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n239), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n225), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n224), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(KEYINPUT74), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT10), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT73), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT8), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n208), .A2(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n257), .B(new_n259), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n219), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n256), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n269), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G1), .B2(new_n208), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n254), .B(KEYINPUT9), .C1(new_n270), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n267), .A2(new_n269), .ZN(new_n277));
  INV_X1    g0077(.A(new_n256), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT73), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(G222), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G77), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT68), .B1(new_n295), .B2(new_n219), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT68), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n220), .A2(new_n297), .A3(new_n294), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT67), .A4(new_n290), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n220), .A2(new_n294), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(new_n302), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G226), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n301), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G190), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(G200), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n270), .A2(KEYINPUT9), .A3(new_n275), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n252), .B(new_n253), .C1(new_n282), .C2(new_n314), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n316));
  AOI211_X1 g0116(.A(new_n256), .B(new_n274), .C1(new_n267), .C2(new_n269), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n254), .B1(new_n317), .B2(KEYINPUT9), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n279), .A2(KEYINPUT73), .A3(new_n280), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n252), .A2(new_n253), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT74), .A2(KEYINPUT10), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n316), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT70), .B(G179), .Z(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n317), .B1(new_n325), .B2(new_n310), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G169), .B2(new_n310), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n315), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT12), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n255), .B2(G68), .ZN(new_n330));
  INV_X1    g0130(.A(new_n255), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n228), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n330), .B(new_n332), .C1(new_n272), .C2(new_n228), .ZN(new_n333));
  XOR2_X1   g0133(.A(new_n333), .B(KEYINPUT75), .Z(new_n334));
  INV_X1    g0134(.A(new_n258), .ZN(new_n335));
  INV_X1    g0135(.A(G77), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n335), .A2(new_n273), .B1(new_n266), .B2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n208), .A2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n269), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT11), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n283), .A2(G226), .A3(new_n285), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n283), .A2(G232), .A3(G1698), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G97), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n304), .B1(new_n345), .B2(new_n299), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n307), .A2(G238), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G200), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(G190), .A3(new_n351), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(KEYINPUT76), .A3(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n349), .A2(G179), .A3(new_n351), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT14), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n352), .A2(KEYINPUT76), .A3(new_n360), .A4(G169), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n341), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n261), .A2(new_n228), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n215), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n258), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT77), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n287), .A2(new_n288), .A3(G20), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(KEYINPUT7), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT77), .B(new_n374), .C1(new_n283), .C2(G20), .ZN(new_n375));
  OR2_X1    g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NAND2_X1  g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n289), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n373), .A2(new_n375), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n370), .B1(new_n382), .B2(new_n228), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n374), .B1(new_n283), .B2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n378), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n369), .B1(new_n387), .B2(G68), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n271), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n265), .A2(new_n255), .ZN(new_n391));
  INV_X1    g0191(.A(new_n272), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n265), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(G226), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n394));
  OAI211_X1 g0194(.A(G223), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT79), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT79), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n394), .A2(new_n395), .A3(new_n399), .A4(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n299), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n307), .A2(G232), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n305), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G200), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n401), .A2(G190), .A3(new_n402), .A4(new_n305), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n390), .A2(new_n393), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n407));
  INV_X1    g0207(.A(new_n393), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n385), .B2(new_n389), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n409), .A2(new_n410), .A3(new_n404), .A4(new_n405), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n409), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n401), .A2(new_n325), .A3(new_n402), .A4(new_n305), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT18), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n409), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n412), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n283), .A2(G232), .A3(new_n285), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n283), .A2(G1698), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n423), .B1(new_n424), .B2(new_n283), .C1(new_n425), .C2(new_n229), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n299), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n307), .A2(G244), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n305), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n414), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n331), .A2(new_n336), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n392), .A2(G77), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G20), .A2(G77), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n433), .B1(new_n263), .B2(new_n335), .C1(new_n266), .C2(new_n434), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n435), .A2(KEYINPUT71), .A3(new_n269), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT71), .B1(new_n435), .B2(new_n269), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT72), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n429), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n325), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n430), .A2(KEYINPUT72), .A3(new_n438), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n438), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n429), .A2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(G190), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n429), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NOR4_X1   g0250(.A1(new_n328), .A2(new_n365), .A3(new_n422), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n207), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n255), .A2(new_n452), .A3(new_n219), .A4(new_n268), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n424), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n208), .A2(G107), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT23), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  XOR2_X1   g0258(.A(new_n458), .B(KEYINPUT86), .Z(new_n459));
  NAND3_X1  g0259(.A1(new_n283), .A2(new_n208), .A3(G87), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(KEYINPUT22), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n456), .B(new_n459), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n460), .B(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n456), .A4(new_n459), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n454), .B1(new_n468), .B2(new_n269), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n255), .A2(G107), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT25), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n283), .A2(G250), .A3(new_n285), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G294), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(new_n425), .C2(new_n231), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(new_n306), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n475), .A2(new_n299), .B1(G264), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n478), .A2(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G274), .A3(new_n477), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(G169), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n472), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n485), .A2(G200), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n486), .A2(G190), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n469), .A2(new_n492), .A3(new_n493), .A4(new_n471), .ZN(new_n494));
  INV_X1    g0294(.A(G200), .ZN(new_n495));
  INV_X1    g0295(.A(new_n484), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n283), .A2(G257), .A3(new_n285), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n283), .A2(G264), .A3(G1698), .ZN(new_n498));
  INV_X1    g0298(.A(G303), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n283), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n500), .B2(new_n299), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n481), .A2(G270), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G283), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n208), .C1(G33), .C2(new_n230), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n505), .B(new_n269), .C1(new_n208), .C2(G116), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n255), .B2(G116), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n453), .B2(new_n224), .ZN(new_n511));
  INV_X1    g0311(.A(new_n453), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n509), .A3(G116), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  OR3_X1    g0314(.A1(new_n503), .A2(new_n514), .A3(KEYINPUT85), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT85), .B1(new_n503), .B2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n501), .A2(new_n502), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n516), .C1(new_n448), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n517), .A3(G169), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT21), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n517), .A2(new_n489), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n514), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT21), .A4(G169), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n491), .A2(new_n494), .A3(new_n518), .A4(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n504), .A4(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n533), .A2(new_n534), .A3(new_n299), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n533), .B2(new_n299), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n480), .A2(new_n306), .A3(G257), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n484), .A2(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT81), .B1(new_n539), .B2(new_n495), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n255), .A2(G97), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n453), .B2(new_n230), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n258), .A2(G77), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n424), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n230), .A2(new_n424), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n545), .B1(new_n548), .B2(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G20), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n544), .B(new_n550), .C1(new_n382), .C2(new_n424), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n543), .B1(new_n551), .B2(new_n269), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n538), .B1(new_n533), .B2(new_n299), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n533), .A2(new_n299), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT80), .ZN(new_n556));
  INV_X1    g0356(.A(new_n538), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n533), .A2(new_n534), .A3(new_n299), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(G200), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n540), .A2(new_n552), .A3(new_n554), .A4(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n434), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n255), .ZN(new_n564));
  INV_X1    g0364(.A(G87), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n453), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n567), .A2(new_n208), .A3(G33), .A4(G97), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n547), .A2(new_n565), .B1(new_n344), .B2(new_n208), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(new_n567), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n208), .B(G68), .C1(new_n287), .C2(new_n288), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n283), .A2(KEYINPUT82), .A3(new_n208), .A4(G68), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI211_X1 g0375(.A(new_n564), .B(new_n566), .C1(new_n575), .C2(new_n269), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n577));
  OAI211_X1 g0377(.A(G238), .B(new_n285), .C1(new_n287), .C2(new_n288), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n457), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n299), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n306), .B(G250), .C1(G1), .C2(new_n476), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n477), .A2(G274), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n580), .A2(G190), .A3(new_n581), .A4(new_n582), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n576), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n575), .A2(new_n269), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n512), .A2(new_n563), .ZN(new_n588));
  INV_X1    g0388(.A(new_n564), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n414), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n580), .A2(new_n325), .A3(new_n581), .A4(new_n582), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n553), .A2(G169), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n539), .B2(new_n325), .ZN(new_n596));
  INV_X1    g0396(.A(new_n552), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n562), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT83), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n562), .A2(KEYINPUT83), .A3(new_n598), .A4(new_n594), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n527), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n451), .A2(new_n603), .ZN(G372));
  OR2_X1    g0404(.A1(new_n356), .A2(new_n445), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n362), .A2(new_n363), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(new_n407), .B2(new_n411), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n419), .B2(new_n421), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n409), .A2(new_n417), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT18), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT7), .B1(new_n289), .B2(new_n208), .ZN(new_n612));
  INV_X1    g0412(.A(new_n378), .ZN(new_n613));
  OAI21_X1  g0413(.A(G68), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n269), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n384), .B2(new_n383), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n416), .B(new_n415), .C1(new_n617), .C2(new_n408), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n420), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(new_n619), .A3(KEYINPUT90), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n323), .B(new_n315), .C1(new_n607), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n327), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n623), .B(KEYINPUT91), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n594), .A2(new_n596), .A3(KEYINPUT26), .A4(new_n597), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n556), .A2(new_n325), .A3(new_n557), .A4(new_n558), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n555), .A2(new_n557), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n414), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(new_n552), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n594), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(KEYINPUT88), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n628), .A2(new_n636), .A3(new_n630), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n552), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n584), .A2(KEYINPUT87), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT87), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n583), .A2(new_n640), .A3(G200), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n639), .A2(new_n585), .A3(new_n576), .A4(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n593), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT26), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n562), .A2(new_n494), .A3(new_n598), .A4(new_n643), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n487), .B1(new_n469), .B2(new_n471), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n525), .B1(new_n647), .B2(new_n490), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n593), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n451), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n624), .A2(new_n651), .ZN(G369));
  NOR2_X1   g0452(.A1(new_n210), .A2(G20), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n207), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n514), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n526), .B1(new_n518), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n661), .B(new_n663), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n491), .ZN(new_n666));
  INV_X1    g0466(.A(new_n659), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n494), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n469), .B2(new_n471), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n491), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n526), .A2(new_n659), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n671), .A2(new_n675), .B1(new_n666), .B2(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(G399));
  NOR2_X1   g0477(.A1(new_n211), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G1), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n547), .A2(new_n565), .A3(new_n224), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n680), .A2(new_n681), .B1(new_n218), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n601), .A2(new_n602), .ZN(new_n684));
  INV_X1    g0484(.A(new_n527), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n667), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT31), .ZN(new_n687));
  INV_X1    g0487(.A(new_n583), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n559), .A2(new_n485), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(KEYINPUT93), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n559), .A2(new_n691), .A3(new_n485), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n690), .A2(new_n325), .A3(new_n517), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n629), .A2(new_n583), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n522), .A2(new_n694), .A3(KEYINPUT30), .A4(new_n482), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n482), .A2(new_n501), .A3(G179), .A4(new_n502), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n688), .A2(new_n553), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  AOI211_X1 g0500(.A(new_n687), .B(new_n667), .C1(new_n693), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n689), .A2(KEYINPUT93), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n583), .A3(new_n517), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n692), .A2(new_n325), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n705), .B2(new_n659), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n686), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT94), .B1(new_n708), .B2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT94), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  AOI211_X1 g0511(.A(new_n710), .B(new_n711), .C1(new_n686), .C2(new_n707), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n491), .A2(new_n526), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n562), .A2(new_n598), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n494), .A2(new_n643), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n714), .A2(new_n715), .A3(new_n716), .A4(KEYINPUT95), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n646), .B2(new_n648), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n632), .A2(new_n721), .A3(new_n594), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n638), .A2(new_n643), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT26), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n720), .A2(new_n593), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n667), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n650), .A2(new_n667), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n713), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n683), .B1(new_n732), .B2(G1), .ZN(G364));
  OR2_X1    g0533(.A1(new_n664), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n653), .A2(G45), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n679), .A2(G1), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n665), .A3(new_n736), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT96), .Z(new_n738));
  AOI21_X1  g0538(.A(new_n219), .B1(G20), .B2(new_n414), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n208), .A2(new_n448), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n324), .A2(new_n495), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G322), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n324), .A2(G20), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  OAI21_X1  g0547(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT101), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n495), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n740), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n499), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n208), .A2(G190), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT99), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n489), .A2(new_n495), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT100), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(new_n750), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G329), .A2(new_n758), .B1(new_n760), .B2(G283), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n324), .A2(new_n495), .A3(new_n753), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n744), .A2(new_n448), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n283), .B1(new_n765), .B2(G326), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n766), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n749), .A2(new_n752), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G159), .ZN(new_n773));
  OR3_X1    g0573(.A1(new_n757), .A2(KEYINPUT32), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT32), .B1(new_n757), .B2(new_n773), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n565), .C2(new_n751), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n283), .B1(new_n261), .B2(new_n741), .C1(new_n769), .C2(new_n230), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n760), .A2(G107), .B1(new_n765), .B2(G50), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n336), .B2(new_n763), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n746), .A2(new_n228), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n739), .B1(new_n772), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n211), .A2(new_n289), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G355), .B1(new_n224), .B2(new_n211), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n247), .A2(G45), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n218), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n211), .A2(new_n283), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT98), .Z(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n739), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n736), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n794), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n782), .B(new_n796), .C1(new_n664), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n738), .A2(new_n798), .ZN(G396));
  INV_X1    g0599(.A(new_n765), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n800), .A2(new_n499), .B1(new_n770), .B2(new_n741), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n759), .A2(new_n565), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n763), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G116), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n758), .A2(G311), .B1(new_n745), .B2(G283), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n289), .B1(new_n751), .B2(new_n424), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n768), .B2(G97), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n803), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n765), .A2(G137), .B1(new_n804), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G143), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n741), .C1(new_n812), .C2(new_n746), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G132), .A2(new_n758), .B1(new_n760), .B2(G68), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n283), .B1(new_n273), .B2(new_n751), .C1(new_n769), .C2(new_n261), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n739), .A2(new_n792), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(new_n739), .B1(new_n336), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n736), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n446), .A2(new_n667), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n445), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(new_n445), .B2(new_n449), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n820), .B(new_n821), .C1(new_n793), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT104), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n823), .A2(new_n824), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT102), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n728), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(KEYINPUT103), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n667), .B(new_n825), .C1(new_n645), .C2(new_n649), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n728), .B2(new_n829), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(KEYINPUT103), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n827), .B1(new_n835), .B2(new_n713), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(KEYINPUT104), .C1(new_n709), .C2(new_n712), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n713), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n826), .B1(new_n839), .B2(new_n821), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n705), .A2(new_n659), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(KEYINPUT109), .A3(new_n687), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n687), .A2(KEYINPUT109), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n705), .A2(new_n659), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n686), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n341), .A2(new_n667), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n365), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n364), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n828), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n609), .A2(new_n412), .A3(new_n620), .ZN(new_n851));
  INV_X1    g0651(.A(new_n657), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n617), .B2(new_n408), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n618), .A2(new_n406), .A3(new_n853), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT108), .B1(new_n856), .B2(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT107), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT37), .B1(new_n618), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n610), .A2(KEYINPUT107), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n860), .A2(new_n406), .A3(new_n861), .A4(new_n853), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n856), .A2(KEYINPUT108), .A3(KEYINPUT37), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n855), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n408), .B1(new_n866), .B2(new_n389), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n657), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n422), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n406), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n867), .B1(new_n417), .B2(new_n657), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n869), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n845), .B(new_n850), .C1(new_n865), .C2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n364), .A2(new_n848), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n846), .B(new_n356), .C1(new_n362), .C2(new_n363), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n825), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n844), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n603), .B2(new_n667), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(new_n842), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n869), .A2(new_n873), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT40), .B1(new_n885), .B2(new_n874), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n876), .A2(KEYINPUT40), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n451), .A2(new_n845), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n887), .B(new_n888), .Z(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(G330), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n877), .A2(new_n878), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n445), .A2(new_n659), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n832), .A2(KEYINPUT105), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT105), .B1(new_n832), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT106), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n885), .A2(new_n874), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n900), .B(new_n892), .C1(new_n895), .C2(new_n896), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  INV_X1    g0703(.A(new_n863), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n904), .A2(new_n857), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n905), .A2(new_n862), .B1(new_n851), .B2(new_n854), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n903), .B(new_n874), .C1(new_n906), .C2(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT38), .B1(new_n869), .B2(new_n873), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT39), .B1(new_n875), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n606), .A2(new_n659), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n910), .A2(new_n911), .B1(new_n621), .B2(new_n657), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n890), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n727), .A2(new_n730), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n451), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(new_n624), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n914), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n207), .B2(new_n653), .ZN(new_n919));
  OAI211_X1 g0719(.A(G20), .B(new_n220), .C1(new_n549), .C2(KEYINPUT35), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n224), .B(new_n920), .C1(KEYINPUT35), .C2(new_n549), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT36), .Z(new_n922));
  NOR3_X1   g0722(.A1(new_n218), .A2(new_n336), .A3(new_n366), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n228), .A2(G50), .ZN(new_n924));
  OAI211_X1 g0724(.A(G1), .B(new_n210), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n919), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI21_X1  g0726(.A(new_n715), .B1(new_n552), .B2(new_n667), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n638), .A2(new_n659), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n598), .B1(new_n929), .B2(new_n491), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n667), .ZN(new_n931));
  INV_X1    g0731(.A(new_n672), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n928), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n675), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT110), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT110), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n934), .A2(KEYINPUT42), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n576), .A2(new_n667), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n643), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n593), .B2(new_n945), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT43), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT111), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n940), .A2(new_n949), .A3(new_n942), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n944), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n944), .B2(new_n950), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n674), .A2(new_n929), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n735), .A2(G1), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n933), .A2(new_n676), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT45), .Z(new_n959));
  NOR2_X1   g0759(.A1(new_n933), .A2(new_n676), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT44), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n959), .A2(new_n674), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n674), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n672), .B(new_n675), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n665), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n731), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n731), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n678), .B(KEYINPUT41), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n957), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n954), .B1(new_n951), .B2(new_n953), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n955), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n768), .A2(G68), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n758), .A2(G137), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n745), .A2(G159), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n765), .A2(G143), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G50), .A2(new_n804), .B1(new_n742), .B2(G150), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n261), .B2(new_n751), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n759), .A2(new_n336), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n978), .A2(new_n980), .A3(new_n289), .A4(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G283), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n289), .B1(new_n983), .B2(new_n763), .C1(new_n757), .C2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n745), .A2(G294), .B1(new_n742), .B2(G303), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n230), .B2(new_n759), .C1(new_n762), .C2(new_n800), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(G107), .C2(new_n768), .ZN(new_n988));
  INV_X1    g0788(.A(new_n751), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n982), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  AOI21_X1  g0793(.A(new_n736), .B1(new_n993), .B2(new_n739), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n795), .B1(new_n212), .B2(new_n434), .C1(new_n243), .C2(new_n789), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n797), .C2(new_n947), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n973), .A2(new_n996), .ZN(G387));
  AOI22_X1  g0797(.A1(new_n745), .A2(G311), .B1(new_n742), .B2(G317), .ZN(new_n998));
  XOR2_X1   g0798(.A(KEYINPUT113), .B(G322), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n765), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(new_n499), .C2(new_n763), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(G283), .B2(new_n768), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n770), .B2(new_n751), .C1(new_n1003), .C2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT49), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n283), .B1(new_n760), .B2(G116), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1007), .B(new_n1010), .C1(G326), .C2(new_n758), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n769), .A2(new_n434), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n283), .C1(new_n230), .C2(new_n759), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n757), .A2(new_n812), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n800), .A2(new_n773), .B1(new_n273), .B2(new_n741), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n989), .A2(G77), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n763), .B2(new_n228), .C1(new_n746), .C2(new_n265), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n739), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n263), .A2(G50), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(G45), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n228), .B2(new_n336), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n681), .B(KEYINPUT112), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(KEYINPUT50), .C2(new_n1022), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n788), .B(new_n1027), .C1(new_n240), .C2(new_n476), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n783), .A2(new_n681), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G107), .C2(new_n212), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n795), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1020), .A2(new_n821), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT115), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n932), .B2(new_n797), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n967), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n679), .B1(new_n731), .B2(new_n966), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1034), .B(new_n1037), .C1(new_n957), .C2(new_n966), .ZN(G393));
  NAND2_X1  g0838(.A1(new_n929), .A2(new_n794), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n795), .B1(new_n230), .B2(new_n212), .C1(new_n250), .C2(new_n789), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n768), .A2(G116), .B1(new_n804), .B2(G294), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n746), .B2(new_n499), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT116), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n765), .A2(G317), .B1(new_n742), .B2(G311), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n283), .B1(new_n989), .B2(G283), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n758), .A2(new_n999), .B1(new_n760), .B2(G107), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n746), .A2(new_n273), .B1(new_n811), .B2(new_n757), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n769), .A2(new_n336), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n264), .C2(new_n804), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n289), .B(new_n802), .C1(G68), .C2(new_n989), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n765), .A2(G150), .B1(new_n742), .B2(G159), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT51), .Z(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1048), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n736), .B1(new_n1056), .B2(new_n739), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1039), .A2(new_n1040), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n964), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n1035), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n964), .A2(new_n967), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n678), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT117), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1058), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n957), .B2(new_n1059), .ZN(G390));
  NAND2_X1  g0867(.A1(new_n845), .A2(new_n850), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1068), .A2(new_n711), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n911), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n910), .B1(new_n897), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n874), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n1071), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n894), .B1(new_n726), .B2(new_n828), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n892), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1070), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n865), .A2(new_n875), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n911), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n724), .A2(new_n593), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n719), .B2(new_n717), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n659), .B1(new_n1081), .B2(new_n722), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n893), .B1(new_n1082), .B2(new_n825), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1083), .B2(new_n891), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n713), .A2(new_n879), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n832), .A2(new_n894), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT105), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n832), .A2(KEYINPUT105), .A3(new_n894), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n911), .B1(new_n1090), .B2(new_n892), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1084), .B(new_n1085), .C1(new_n1091), .C2(new_n910), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n829), .A2(new_n845), .A3(G330), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n891), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n1083), .C1(new_n713), .C2(new_n879), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n825), .B1(new_n709), .B2(new_n712), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1069), .B1(new_n1097), .B2(new_n891), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1090), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n451), .A2(new_n845), .A3(G330), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n916), .A2(new_n624), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n678), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT118), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1093), .A2(new_n957), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n289), .B1(new_n758), .B2(G125), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n273), .B2(new_n759), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT120), .Z(new_n1113));
  NAND2_X1  g0913(.A1(new_n765), .A2(G128), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n763), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n989), .A2(G150), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n745), .A2(G137), .B1(KEYINPUT53), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n769), .B2(new_n773), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1117), .B(new_n1120), .C1(G132), .C2(new_n742), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1113), .B(new_n1121), .C1(KEYINPUT53), .C2(new_n1118), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n763), .A2(new_n230), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n746), .A2(new_n424), .B1(new_n224), .B2(new_n741), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1050), .A2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n758), .A2(G294), .B1(new_n765), .B2(G283), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n289), .B1(new_n759), .B2(new_n228), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(G87), .B2(new_n989), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1122), .B1(new_n1123), .B2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1130), .A2(new_n739), .B1(new_n265), .B2(new_n819), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n821), .B(new_n1131), .C1(new_n910), .C2(new_n793), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1109), .A2(new_n1110), .A3(new_n1132), .ZN(G378));
  OAI21_X1  g0933(.A(new_n1102), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(KEYINPUT57), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT122), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT56), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n317), .A2(new_n657), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n328), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT55), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1138), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n315), .A2(new_n323), .A3(new_n327), .A4(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT55), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(KEYINPUT56), .A3(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1145), .A2(new_n1149), .A3(KEYINPUT121), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n887), .B2(new_n711), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1145), .A2(new_n1149), .A3(KEYINPUT121), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT40), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n882), .B2(new_n1073), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n875), .B2(new_n908), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n1068), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1152), .B(G330), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1136), .B1(new_n913), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n913), .A2(new_n1158), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n902), .A2(new_n1151), .A3(new_n912), .A4(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1162), .B2(new_n1136), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n678), .B1(new_n1135), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT123), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1134), .A2(new_n1162), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT57), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT123), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n678), .C1(new_n1135), .C2(new_n1163), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1162), .A2(new_n956), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1145), .A2(new_n1149), .A3(new_n792), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n819), .A2(new_n273), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n765), .A2(G125), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n742), .A2(G128), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n751), .C2(new_n1116), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n804), .A2(G137), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n769), .B2(new_n812), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G132), .C2(new_n745), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT59), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G41), .B1(new_n758), .B2(G124), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G33), .B1(new_n760), .B2(G159), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n273), .B1(new_n287), .B2(G41), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n974), .B(new_n289), .C1(new_n224), .C2(new_n800), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n746), .A2(new_n230), .B1(new_n983), .B2(new_n757), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n759), .A2(new_n261), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n742), .A2(G107), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n804), .A2(new_n563), .ZN(new_n1189));
  INV_X1    g0989(.A(G41), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1017), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT58), .Z(new_n1193));
  NAND3_X1  g0993(.A1(new_n1183), .A2(new_n1184), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n736), .B1(new_n1194), .B2(new_n739), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1172), .A2(new_n1173), .A3(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1171), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1170), .A2(new_n1197), .ZN(G375));
  OR2_X1    g0998(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n969), .A3(new_n1103), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n283), .B(new_n981), .C1(G97), .C2(new_n989), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n758), .A2(G303), .B1(new_n765), .B2(G294), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n745), .A2(G116), .B1(new_n742), .B2(G283), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1013), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n763), .A2(new_n424), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n758), .A2(G128), .B1(G150), .B2(new_n804), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n261), .B2(new_n759), .C1(new_n746), .C2(new_n1116), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n768), .A2(G50), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n765), .A2(G132), .B1(new_n742), .B2(G137), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n989), .A2(G159), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n283), .A4(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n1204), .A2(new_n1205), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1212), .A2(new_n739), .B1(new_n228), .B2(new_n819), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n821), .B(new_n1213), .C1(new_n892), .C2(new_n793), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1100), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1214), .B1(new_n1215), .B2(new_n957), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1200), .A2(new_n1217), .ZN(G381));
  NOR2_X1   g1018(.A1(G375), .A2(G378), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G387), .A2(G381), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(G393), .A2(G396), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(G390), .A2(G384), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1223), .ZN(G407));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n658), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(G407), .A2(G213), .A3(new_n1225), .ZN(G409));
  NAND3_X1  g1026(.A1(new_n1170), .A2(G378), .A3(new_n1197), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1166), .A2(new_n969), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n1196), .C1(new_n957), .C2(new_n1163), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1229), .A2(new_n1110), .A3(new_n1109), .A4(new_n1132), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT124), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n658), .A2(G213), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(G384), .B(KEYINPUT125), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1199), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1102), .B2(new_n1100), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n679), .B1(new_n1199), .B2(new_n1236), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1216), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1235), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1227), .A2(new_n1230), .A3(KEYINPUT124), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1233), .A2(new_n1234), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT126), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1231), .A2(new_n1246), .A3(new_n1234), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1252), .A2(new_n1249), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G393), .A2(G396), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1059), .A2(new_n957), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1255), .B(new_n1058), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G387), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1222), .B(new_n1254), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(G387), .A2(new_n1256), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1259), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G390), .A2(new_n996), .A3(new_n973), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1221), .B1(new_n1262), .B2(KEYINPUT127), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1260), .A2(new_n1257), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1254), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1253), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1233), .A2(new_n1234), .A3(new_n1247), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1245), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1241), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1269), .B2(new_n1241), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1248), .A2(new_n1275), .A3(new_n1249), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1251), .A2(new_n1267), .A3(new_n1274), .A4(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1252), .B2(KEYINPUT62), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1278), .B(new_n1280), .C1(KEYINPUT62), .C2(new_n1248), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1266), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(G405));
  NAND2_X1  g1083(.A1(new_n1266), .A2(new_n1246), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1261), .B(new_n1265), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G375), .B(G378), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1286), .B(new_n1288), .ZN(G402));
endmodule


