

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742;

  XNOR2_X2 U375 ( .A(n550), .B(n549), .ZN(n742) );
  XNOR2_X1 U376 ( .A(n497), .B(n450), .ZN(n456) );
  XNOR2_X2 U377 ( .A(n438), .B(KEYINPUT67), .ZN(n509) );
  XNOR2_X2 U378 ( .A(G131), .B(KEYINPUT68), .ZN(n438) );
  XNOR2_X2 U379 ( .A(n396), .B(KEYINPUT35), .ZN(n738) );
  NOR2_X1 U380 ( .A1(n587), .A2(n574), .ZN(n566) );
  INV_X1 U381 ( .A(n591), .ZN(n365) );
  INV_X2 U382 ( .A(G953), .ZN(n730) );
  XNOR2_X1 U383 ( .A(n519), .B(n372), .ZN(n644) );
  XNOR2_X1 U384 ( .A(n439), .B(KEYINPUT40), .ZN(n741) );
  NAND2_X1 U385 ( .A1(n644), .A2(n648), .ZN(n660) );
  NAND2_X1 U386 ( .A1(n675), .A2(n674), .ZN(n587) );
  NOR2_X1 U387 ( .A1(n547), .A2(n546), .ZN(n658) );
  XNOR2_X1 U388 ( .A(G104), .B(G122), .ZN(n371) );
  AND2_X1 U389 ( .A1(n407), .A2(n406), .ZN(n405) );
  NOR2_X1 U390 ( .A1(n366), .A2(n373), .ZN(n417) );
  NAND2_X1 U391 ( .A1(n495), .A2(n494), .ZN(n532) );
  NAND2_X1 U392 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U393 ( .A(n591), .B(n536), .ZN(n574) );
  XNOR2_X1 U394 ( .A(n384), .B(n479), .ZN(n669) );
  XNOR2_X1 U395 ( .A(n467), .B(G469), .ZN(n535) );
  XNOR2_X1 U396 ( .A(n420), .B(n419), .ZN(n546) );
  NOR2_X1 U397 ( .A1(n707), .A2(G902), .ZN(n467) );
  XNOR2_X1 U398 ( .A(n466), .B(n441), .ZN(n707) );
  XNOR2_X1 U399 ( .A(n454), .B(n453), .ZN(n718) );
  XNOR2_X1 U400 ( .A(n401), .B(n400), .ZN(n453) );
  INV_X1 U401 ( .A(n371), .ZN(n510) );
  XNOR2_X1 U402 ( .A(n435), .B(G128), .ZN(n497) );
  BUF_X1 U403 ( .A(n599), .Z(n353) );
  INV_X1 U404 ( .A(n584), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n375), .B(n597), .ZN(n599) );
  XNOR2_X1 U406 ( .A(n535), .B(n534), .ZN(n675) );
  XNOR2_X2 U407 ( .A(n398), .B(n456), .ZN(n727) );
  XNOR2_X1 U408 ( .A(n368), .B(G146), .ZN(n471) );
  INV_X1 U409 ( .A(G125), .ZN(n368) );
  INV_X1 U410 ( .A(G143), .ZN(n435) );
  INV_X1 U411 ( .A(KEYINPUT83), .ZN(n427) );
  XNOR2_X1 U412 ( .A(n509), .B(n436), .ZN(n398) );
  XNOR2_X1 U413 ( .A(n437), .B(G134), .ZN(n436) );
  INV_X1 U414 ( .A(G137), .ZN(n437) );
  XOR2_X1 U415 ( .A(n556), .B(KEYINPUT38), .Z(n657) );
  XNOR2_X1 U416 ( .A(n517), .B(G475), .ZN(n419) );
  OR2_X1 U417 ( .A1(n621), .A2(G902), .ZN(n420) );
  XNOR2_X1 U418 ( .A(n551), .B(KEYINPUT46), .ZN(n366) );
  NOR2_X1 U419 ( .A1(n738), .A2(KEYINPUT65), .ZN(n582) );
  XNOR2_X1 U420 ( .A(KEYINPUT75), .B(KEYINPUT74), .ZN(n446) );
  XOR2_X1 U421 ( .A(G116), .B(KEYINPUT5), .Z(n447) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n450) );
  XNOR2_X1 U423 ( .A(n471), .B(n409), .ZN(n408) );
  XNOR2_X1 U424 ( .A(n457), .B(KEYINPUT17), .ZN(n409) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n415) );
  AND2_X1 U426 ( .A1(n669), .A2(n521), .ZN(n538) );
  NOR2_X1 U427 ( .A1(n520), .A2(n668), .ZN(n521) );
  NAND2_X1 U428 ( .A1(n365), .A2(n553), .ZN(n431) );
  INV_X1 U429 ( .A(KEYINPUT100), .ZN(n377) );
  NOR2_X1 U430 ( .A1(n669), .A2(n668), .ZN(n674) );
  XNOR2_X1 U431 ( .A(G116), .B(G107), .ZN(n498) );
  XNOR2_X1 U432 ( .A(n442), .B(n444), .ZN(n400) );
  INV_X1 U433 ( .A(KEYINPUT69), .ZN(n444) );
  XNOR2_X1 U434 ( .A(n478), .B(n477), .ZN(n615) );
  XNOR2_X1 U435 ( .A(n476), .B(n440), .ZN(n477) );
  XNOR2_X1 U436 ( .A(n394), .B(n393), .ZN(n496) );
  XNOR2_X1 U437 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n393) );
  XNOR2_X1 U438 ( .A(n395), .B(KEYINPUT66), .ZN(n394) );
  NAND2_X1 U439 ( .A1(n730), .A2(G234), .ZN(n395) );
  XNOR2_X1 U440 ( .A(G134), .B(G122), .ZN(n500) );
  XNOR2_X1 U441 ( .A(n502), .B(n503), .ZN(n379) );
  AND2_X1 U442 ( .A1(n383), .A2(n423), .ZN(n380) );
  NOR2_X1 U443 ( .A1(n598), .A2(n427), .ZN(n426) );
  AND2_X1 U444 ( .A1(n392), .A2(n391), .ZN(n387) );
  NAND2_X1 U445 ( .A1(n532), .A2(n363), .ZN(n392) );
  INV_X1 U446 ( .A(KEYINPUT96), .ZN(n418) );
  XNOR2_X1 U447 ( .A(n506), .B(n378), .ZN(n547) );
  INV_X1 U448 ( .A(G478), .ZN(n378) );
  INV_X1 U449 ( .A(KEYINPUT77), .ZN(n410) );
  AND2_X1 U450 ( .A1(n642), .A2(n414), .ZN(n413) );
  XNOR2_X1 U451 ( .A(G137), .B(G128), .ZN(n473) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n482) );
  OR2_X1 U453 ( .A1(G237), .A2(G902), .ZN(n492) );
  XNOR2_X1 U454 ( .A(n466), .B(n449), .ZN(n490) );
  XNOR2_X1 U455 ( .A(n448), .B(n360), .ZN(n399) );
  NAND2_X1 U456 ( .A1(n598), .A2(n427), .ZN(n424) );
  XNOR2_X1 U457 ( .A(G902), .B(KEYINPUT15), .ZN(n598) );
  XNOR2_X1 U458 ( .A(G101), .B(G104), .ZN(n460) );
  XOR2_X1 U459 ( .A(G140), .B(G107), .Z(n461) );
  XNOR2_X1 U460 ( .A(n718), .B(n428), .ZN(n607) );
  XNOR2_X1 U461 ( .A(n455), .B(KEYINPUT18), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n456), .B(n408), .ZN(n458) );
  AND2_X1 U463 ( .A1(n653), .A2(n433), .ZN(n432) );
  INV_X1 U464 ( .A(n652), .ZN(n433) );
  XNOR2_X1 U465 ( .A(n369), .B(KEYINPUT41), .ZN(n686) );
  NOR2_X1 U466 ( .A1(n615), .A2(G902), .ZN(n384) );
  XNOR2_X1 U467 ( .A(n431), .B(KEYINPUT30), .ZN(n430) );
  INV_X1 U468 ( .A(KEYINPUT104), .ZN(n381) );
  XNOR2_X1 U469 ( .A(n571), .B(n377), .ZN(n376) );
  NAND2_X1 U470 ( .A1(n674), .A2(n523), .ZN(n589) );
  XNOR2_X1 U471 ( .A(n379), .B(n501), .ZN(n504) );
  NAND2_X1 U472 ( .A1(n385), .A2(n387), .ZN(n439) );
  AND2_X1 U473 ( .A1(n386), .A2(n388), .ZN(n385) );
  INV_X1 U474 ( .A(n568), .ZN(n569) );
  AND2_X1 U475 ( .A1(n548), .A2(n564), .ZN(n642) );
  INV_X1 U476 ( .A(KEYINPUT98), .ZN(n372) );
  NOR2_X1 U477 ( .A1(n518), .A2(n547), .ZN(n519) );
  XNOR2_X1 U478 ( .A(n709), .B(n708), .ZN(n710) );
  AND2_X1 U479 ( .A1(n543), .A2(n651), .ZN(n355) );
  XOR2_X1 U480 ( .A(KEYINPUT12), .B(KEYINPUT94), .Z(n356) );
  AND2_X1 U481 ( .A1(G210), .A2(n492), .ZN(n357) );
  XOR2_X1 U482 ( .A(n660), .B(KEYINPUT79), .Z(n358) );
  XNOR2_X1 U483 ( .A(KEYINPUT72), .B(n544), .ZN(n359) );
  AND2_X1 U484 ( .A1(n511), .A2(G210), .ZN(n360) );
  XNOR2_X1 U485 ( .A(n453), .B(n399), .ZN(n449) );
  AND2_X1 U486 ( .A1(n425), .A2(n424), .ZN(n361) );
  NAND2_X1 U487 ( .A1(n531), .A2(KEYINPUT47), .ZN(n362) );
  INV_X1 U488 ( .A(n644), .ZN(n388) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n363) );
  OR2_X1 U490 ( .A1(n598), .A2(n698), .ZN(n364) );
  XNOR2_X2 U491 ( .A(n491), .B(G472), .ZN(n591) );
  AND2_X2 U492 ( .A1(n367), .A2(n364), .ZN(n600) );
  NAND2_X1 U493 ( .A1(n380), .A2(n361), .ZN(n367) );
  NAND2_X1 U494 ( .A1(n661), .A2(n658), .ZN(n369) );
  NAND2_X1 U495 ( .A1(n434), .A2(n432), .ZN(n729) );
  XNOR2_X1 U496 ( .A(n443), .B(n445), .ZN(n401) );
  NAND2_X1 U497 ( .A1(n526), .A2(n553), .ZN(n539) );
  BUF_X1 U498 ( .A(n353), .Z(n370) );
  NAND2_X1 U499 ( .A1(n412), .A2(KEYINPUT2), .ZN(n411) );
  NOR2_X1 U500 ( .A1(n490), .A2(G902), .ZN(n491) );
  NOR2_X1 U501 ( .A1(n654), .A2(n590), .ZN(n567) );
  INV_X1 U502 ( .A(n729), .ZN(n383) );
  NOR2_X1 U503 ( .A1(n644), .A2(n574), .ZN(n537) );
  NOR2_X1 U504 ( .A1(n579), .A2(n365), .ZN(n580) );
  NAND2_X1 U505 ( .A1(n355), .A2(n362), .ZN(n373) );
  XNOR2_X1 U506 ( .A(n546), .B(n418), .ZN(n518) );
  XNOR2_X1 U507 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X2 U508 ( .A(n727), .B(G146), .ZN(n466) );
  XNOR2_X2 U509 ( .A(n374), .B(n410), .ZN(n702) );
  NOR2_X2 U510 ( .A1(n411), .A2(n729), .ZN(n374) );
  NAND2_X1 U511 ( .A1(n402), .A2(n405), .ZN(n375) );
  NOR2_X1 U512 ( .A1(n590), .A2(n376), .ZN(n573) );
  XNOR2_X1 U513 ( .A(n382), .B(n381), .ZN(n548) );
  NAND2_X1 U514 ( .A1(n525), .A2(n524), .ZN(n382) );
  NAND2_X1 U515 ( .A1(n390), .A2(n389), .ZN(n386) );
  NAND2_X1 U516 ( .A1(n387), .A2(n386), .ZN(n545) );
  NOR2_X1 U517 ( .A1(n657), .A2(n363), .ZN(n389) );
  INV_X1 U518 ( .A(n532), .ZN(n390) );
  NAND2_X1 U519 ( .A1(n657), .A2(n363), .ZN(n391) );
  NAND2_X1 U520 ( .A1(n397), .A2(n569), .ZN(n396) );
  XNOR2_X1 U521 ( .A(n567), .B(KEYINPUT34), .ZN(n397) );
  XNOR2_X1 U522 ( .A(n404), .B(n403), .ZN(n402) );
  INV_X1 U523 ( .A(KEYINPUT44), .ZN(n403) );
  NAND2_X1 U524 ( .A1(n421), .A2(n582), .ZN(n404) );
  NOR2_X1 U525 ( .A1(n595), .A2(n596), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n583), .A2(n421), .ZN(n407) );
  XNOR2_X1 U527 ( .A(n458), .B(n429), .ZN(n428) );
  NOR2_X1 U528 ( .A1(n430), .A2(n520), .ZN(n494) );
  NAND2_X1 U529 ( .A1(n359), .A2(n417), .ZN(n416) );
  NOR2_X1 U530 ( .A1(n739), .A2(n636), .ZN(n421) );
  INV_X1 U531 ( .A(n599), .ZN(n412) );
  XNOR2_X1 U532 ( .A(n416), .B(n415), .ZN(n434) );
  NOR2_X4 U533 ( .A1(n600), .A2(n702), .ZN(n712) );
  NAND2_X1 U534 ( .A1(n413), .A2(n358), .ZN(n544) );
  INV_X1 U535 ( .A(KEYINPUT47), .ZN(n414) );
  NAND2_X1 U536 ( .A1(n422), .A2(n576), .ZN(n578) );
  AND2_X1 U537 ( .A1(n422), .A2(n584), .ZN(n585) );
  NOR2_X2 U538 ( .A1(n579), .A2(n575), .ZN(n422) );
  NAND2_X1 U539 ( .A1(n412), .A2(n426), .ZN(n423) );
  NAND2_X1 U540 ( .A1(n353), .A2(n427), .ZN(n425) );
  INV_X1 U541 ( .A(n526), .ZN(n556) );
  NAND2_X1 U542 ( .A1(n539), .A2(KEYINPUT19), .ZN(n530) );
  XNOR2_X2 U543 ( .A(n459), .B(n357), .ZN(n526) );
  XNOR2_X1 U544 ( .A(n573), .B(n572), .ZN(n579) );
  XNOR2_X1 U545 ( .A(n475), .B(KEYINPUT24), .ZN(n440) );
  XOR2_X1 U546 ( .A(n465), .B(n464), .Z(n441) );
  XNOR2_X1 U547 ( .A(n513), .B(n512), .ZN(n514) );
  INV_X1 U548 ( .A(KEYINPUT6), .ZN(n536) );
  XNOR2_X1 U549 ( .A(KEYINPUT22), .B(KEYINPUT71), .ZN(n572) );
  INV_X1 U550 ( .A(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U551 ( .A(n707), .B(n706), .ZN(n708) );
  INV_X1 U552 ( .A(KEYINPUT60), .ZN(n626) );
  XOR2_X1 U553 ( .A(G119), .B(G101), .Z(n443) );
  XNOR2_X1 U554 ( .A(KEYINPUT89), .B(KEYINPUT70), .ZN(n442) );
  XNOR2_X1 U555 ( .A(G113), .B(KEYINPUT3), .ZN(n445) );
  XNOR2_X1 U556 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U557 ( .A1(G953), .A2(G237), .ZN(n511) );
  XOR2_X1 U558 ( .A(n490), .B(KEYINPUT62), .Z(n602) );
  XOR2_X2 U559 ( .A(G110), .B(KEYINPUT76), .Z(n463) );
  XOR2_X1 U560 ( .A(KEYINPUT16), .B(n463), .Z(n452) );
  XOR2_X1 U561 ( .A(n510), .B(n498), .Z(n451) );
  XNOR2_X1 U562 ( .A(n452), .B(n451), .ZN(n454) );
  NAND2_X1 U563 ( .A1(G224), .A2(n730), .ZN(n455) );
  INV_X1 U564 ( .A(KEYINPUT90), .ZN(n457) );
  NAND2_X1 U565 ( .A1(n607), .A2(n598), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U567 ( .A(n463), .B(n462), .Z(n465) );
  NAND2_X1 U568 ( .A1(G227), .A2(n730), .ZN(n464) );
  INV_X1 U569 ( .A(n535), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n470) );
  NAND2_X1 U571 ( .A1(n598), .A2(G234), .ZN(n468) );
  XNOR2_X1 U572 ( .A(n468), .B(KEYINPUT20), .ZN(n480) );
  NAND2_X1 U573 ( .A1(n480), .A2(G217), .ZN(n469) );
  XNOR2_X1 U574 ( .A(n470), .B(n469), .ZN(n479) );
  XNOR2_X1 U575 ( .A(n471), .B(KEYINPUT10), .ZN(n472) );
  XNOR2_X1 U576 ( .A(n472), .B(G140), .ZN(n726) );
  XNOR2_X1 U577 ( .A(n726), .B(KEYINPUT23), .ZN(n478) );
  NAND2_X1 U578 ( .A1(G221), .A2(n496), .ZN(n476) );
  XOR2_X1 U579 ( .A(G110), .B(G119), .Z(n474) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U581 ( .A1(G221), .A2(n480), .ZN(n481) );
  XOR2_X1 U582 ( .A(KEYINPUT21), .B(n481), .Z(n570) );
  INV_X1 U583 ( .A(n570), .ZN(n668) );
  XOR2_X1 U584 ( .A(KEYINPUT102), .B(n589), .Z(n495) );
  XOR2_X1 U585 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n483) );
  XNOR2_X1 U586 ( .A(n483), .B(n482), .ZN(n485) );
  NAND2_X1 U587 ( .A1(n485), .A2(G952), .ZN(n484) );
  XOR2_X1 U588 ( .A(KEYINPUT92), .B(n484), .Z(n691) );
  NAND2_X1 U589 ( .A1(n730), .A2(n691), .ZN(n561) );
  INV_X1 U590 ( .A(n561), .ZN(n489) );
  NAND2_X1 U591 ( .A1(G902), .A2(n485), .ZN(n558) );
  NOR2_X1 U592 ( .A1(G900), .A2(n558), .ZN(n486) );
  NAND2_X1 U593 ( .A1(G953), .A2(n486), .ZN(n487) );
  XNOR2_X1 U594 ( .A(KEYINPUT101), .B(n487), .ZN(n488) );
  NOR2_X1 U595 ( .A1(n489), .A2(n488), .ZN(n520) );
  NAND2_X1 U596 ( .A1(n492), .A2(G214), .ZN(n493) );
  XNOR2_X1 U597 ( .A(KEYINPUT91), .B(n493), .ZN(n656) );
  NAND2_X1 U598 ( .A1(G217), .A2(n496), .ZN(n505) );
  XNOR2_X1 U599 ( .A(KEYINPUT97), .B(KEYINPUT7), .ZN(n503) );
  XNOR2_X1 U600 ( .A(n497), .B(KEYINPUT9), .ZN(n502) );
  INV_X1 U601 ( .A(n498), .ZN(n499) );
  XOR2_X1 U602 ( .A(n500), .B(n499), .Z(n501) );
  XNOR2_X1 U603 ( .A(n505), .B(n504), .ZN(n711) );
  NOR2_X1 U604 ( .A1(n711), .A2(G902), .ZN(n506) );
  XNOR2_X1 U605 ( .A(G143), .B(G113), .ZN(n507) );
  XNOR2_X1 U606 ( .A(n356), .B(n507), .ZN(n508) );
  XOR2_X1 U607 ( .A(n509), .B(n508), .Z(n515) );
  XNOR2_X1 U608 ( .A(n510), .B(KEYINPUT11), .ZN(n513) );
  NAND2_X1 U609 ( .A1(G214), .A2(n511), .ZN(n512) );
  XNOR2_X1 U610 ( .A(n726), .B(n516), .ZN(n621) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(KEYINPUT95), .ZN(n517) );
  NAND2_X1 U612 ( .A1(n547), .A2(n518), .ZN(n648) );
  NOR2_X1 U613 ( .A1(n545), .A2(n648), .ZN(n652) );
  AND2_X1 U614 ( .A1(n365), .A2(n538), .ZN(n522) );
  XNOR2_X1 U615 ( .A(n522), .B(KEYINPUT28), .ZN(n525) );
  XOR2_X1 U616 ( .A(n523), .B(KEYINPUT103), .Z(n524) );
  INV_X1 U617 ( .A(n656), .ZN(n553) );
  INV_X1 U618 ( .A(KEYINPUT19), .ZN(n527) );
  AND2_X1 U619 ( .A1(n527), .A2(n553), .ZN(n528) );
  NAND2_X1 U620 ( .A1(n526), .A2(n528), .ZN(n529) );
  NAND2_X1 U621 ( .A1(n530), .A2(n529), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n660), .A2(n642), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n547), .A2(n546), .ZN(n568) );
  NOR2_X1 U624 ( .A1(n532), .A2(n568), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n526), .A2(n533), .ZN(n641) );
  XNOR2_X1 U626 ( .A(KEYINPUT80), .B(n641), .ZN(n543) );
  NAND2_X1 U627 ( .A1(n538), .A2(n537), .ZN(n552) );
  NOR2_X1 U628 ( .A1(n552), .A2(n539), .ZN(n541) );
  XNOR2_X1 U629 ( .A(KEYINPUT106), .B(KEYINPUT36), .ZN(n540) );
  XNOR2_X1 U630 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n354), .A2(n542), .ZN(n651) );
  XOR2_X1 U632 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n550) );
  NOR2_X1 U633 ( .A1(n656), .A2(n657), .ZN(n661) );
  NAND2_X1 U634 ( .A1(n686), .A2(n548), .ZN(n549) );
  NAND2_X1 U635 ( .A1(n741), .A2(n742), .ZN(n551) );
  NOR2_X1 U636 ( .A1(n354), .A2(n552), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U638 ( .A(n555), .B(KEYINPUT43), .ZN(n557) );
  NAND2_X1 U639 ( .A1(n557), .A2(n556), .ZN(n653) );
  INV_X1 U640 ( .A(n558), .ZN(n559) );
  NOR2_X1 U641 ( .A1(G898), .A2(n730), .ZN(n717) );
  NAND2_X1 U642 ( .A1(n559), .A2(n717), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U644 ( .A(KEYINPUT93), .B(n562), .Z(n563) );
  XNOR2_X2 U645 ( .A(n565), .B(KEYINPUT0), .ZN(n590) );
  XNOR2_X1 U646 ( .A(n566), .B(KEYINPUT33), .ZN(n654) );
  AND2_X1 U647 ( .A1(n570), .A2(n658), .ZN(n571) );
  INV_X1 U648 ( .A(n574), .ZN(n575) );
  AND2_X1 U649 ( .A1(n675), .A2(n669), .ZN(n576) );
  INV_X1 U650 ( .A(KEYINPUT32), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n578), .B(n577), .ZN(n739) );
  INV_X1 U652 ( .A(n669), .ZN(n586) );
  INV_X1 U653 ( .A(n675), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n584), .A2(n580), .ZN(n581) );
  NOR2_X1 U655 ( .A1(n586), .A2(n581), .ZN(n636) );
  AND2_X1 U656 ( .A1(n738), .A2(KEYINPUT65), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n628) );
  INV_X1 U658 ( .A(n628), .ZN(n596) );
  OR2_X1 U659 ( .A1(n591), .A2(n587), .ZN(n681) );
  NOR2_X1 U660 ( .A1(n590), .A2(n681), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT31), .B(n588), .ZN(n647) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n632) );
  NAND2_X1 U664 ( .A1(n647), .A2(n632), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n593), .A2(n358), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT99), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n597) );
  INV_X1 U668 ( .A(KEYINPUT2), .ZN(n698) );
  NAND2_X1 U669 ( .A1(n712), .A2(G472), .ZN(n601) );
  XNOR2_X1 U670 ( .A(n602), .B(n601), .ZN(n604) );
  NOR2_X1 U671 ( .A1(G952), .A2(n730), .ZN(n603) );
  XNOR2_X1 U672 ( .A(KEYINPUT88), .B(n603), .ZN(n715) );
  INV_X1 U673 ( .A(n715), .ZN(n624) );
  NAND2_X1 U674 ( .A1(n604), .A2(n624), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT63), .B(KEYINPUT107), .Z(n605) );
  XNOR2_X1 U676 ( .A(n606), .B(n605), .ZN(G57) );
  NAND2_X1 U677 ( .A1(G210), .A2(n712), .ZN(n611) );
  XNOR2_X1 U678 ( .A(KEYINPUT55), .B(KEYINPUT87), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT54), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n612), .A2(n624), .ZN(n614) );
  XNOR2_X1 U683 ( .A(KEYINPUT56), .B(KEYINPUT85), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n614), .B(n613), .ZN(G51) );
  NAND2_X1 U685 ( .A1(G217), .A2(n712), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT123), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n618), .A2(n624), .ZN(n620) );
  INV_X1 U689 ( .A(KEYINPUT124), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(n619), .ZN(G66) );
  NAND2_X1 U691 ( .A1(G475), .A2(n712), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT59), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U695 ( .A(n627), .B(n626), .ZN(G60) );
  XNOR2_X1 U696 ( .A(G101), .B(KEYINPUT108), .ZN(n629) );
  XNOR2_X1 U697 ( .A(n629), .B(n628), .ZN(G3) );
  NOR2_X1 U698 ( .A1(n644), .A2(n632), .ZN(n631) );
  XNOR2_X1 U699 ( .A(G104), .B(KEYINPUT109), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(G6) );
  NOR2_X1 U701 ( .A1(n648), .A2(n632), .ZN(n634) );
  XNOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U704 ( .A(G107), .B(n635), .ZN(G9) );
  XOR2_X1 U705 ( .A(G110), .B(n636), .Z(G12) );
  XOR2_X1 U706 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n639) );
  INV_X1 U707 ( .A(n648), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n642), .A2(n637), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U710 ( .A(G128), .B(n640), .ZN(G30) );
  XNOR2_X1 U711 ( .A(G143), .B(n641), .ZN(G45) );
  NAND2_X1 U712 ( .A1(n388), .A2(n642), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(G146), .ZN(G48) );
  NOR2_X1 U714 ( .A1(n644), .A2(n647), .ZN(n646) );
  XNOR2_X1 U715 ( .A(G113), .B(KEYINPUT111), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G15) );
  NOR2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U718 ( .A(G116), .B(n649), .Z(G18) );
  XOR2_X1 U719 ( .A(G125), .B(KEYINPUT37), .Z(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(G27) );
  XOR2_X1 U721 ( .A(G134), .B(n652), .Z(G36) );
  XNOR2_X1 U722 ( .A(G140), .B(n653), .ZN(G42) );
  INV_X1 U723 ( .A(n654), .ZN(n666) );
  NAND2_X1 U724 ( .A1(n686), .A2(n666), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(KEYINPUT120), .ZN(n694) );
  NAND2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U729 ( .A(KEYINPUT118), .B(n662), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U731 ( .A(KEYINPUT119), .B(n665), .Z(n667) );
  NAND2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n689) );
  XOR2_X1 U733 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n684) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT49), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(KEYINPUT112), .ZN(n672) );
  NOR2_X1 U737 ( .A1(n365), .A2(n672), .ZN(n673) );
  XOR2_X1 U738 ( .A(KEYINPUT113), .B(n673), .Z(n680) );
  XOR2_X1 U739 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n677) );
  OR2_X1 U740 ( .A1(n354), .A2(n674), .ZN(n676) );
  XNOR2_X1 U741 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U742 ( .A(KEYINPUT114), .B(n678), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U744 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n685), .Z(n687) );
  NAND2_X1 U747 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(KEYINPUT52), .ZN(n692) );
  NAND2_X1 U750 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n695), .B(KEYINPUT121), .ZN(n696) );
  NAND2_X1 U753 ( .A1(n696), .A2(n730), .ZN(n704) );
  NAND2_X1 U754 ( .A1(n698), .A2(n370), .ZN(n697) );
  XNOR2_X1 U755 ( .A(n697), .B(KEYINPUT82), .ZN(n700) );
  NAND2_X1 U756 ( .A1(n698), .A2(n729), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U758 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U759 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U760 ( .A(KEYINPUT53), .B(n705), .ZN(G75) );
  NAND2_X1 U761 ( .A1(n712), .A2(G469), .ZN(n709) );
  XOR2_X1 U762 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  NOR2_X1 U763 ( .A1(n710), .A2(n715), .ZN(G54) );
  XNOR2_X1 U764 ( .A(n711), .B(KEYINPUT122), .ZN(n714) );
  NAND2_X1 U765 ( .A1(G478), .A2(n712), .ZN(n713) );
  XNOR2_X1 U766 ( .A(n714), .B(n713), .ZN(n716) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(G63) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n725) );
  NOR2_X1 U769 ( .A1(G953), .A2(n370), .ZN(n719) );
  XNOR2_X1 U770 ( .A(n719), .B(KEYINPUT125), .ZN(n723) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U773 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n725), .B(n724), .ZN(G69) );
  XOR2_X1 U776 ( .A(n726), .B(n727), .Z(n728) );
  XNOR2_X1 U777 ( .A(KEYINPUT126), .B(n728), .ZN(n732) );
  XNOR2_X1 U778 ( .A(n729), .B(n732), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U780 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U782 ( .A1(G953), .A2(n734), .ZN(n735) );
  XOR2_X1 U783 ( .A(KEYINPUT127), .B(n735), .Z(n736) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(G72) );
  XOR2_X1 U785 ( .A(n738), .B(G122), .Z(G24) );
  BUF_X1 U786 ( .A(n739), .Z(n740) );
  XOR2_X1 U787 ( .A(G119), .B(n740), .Z(G21) );
  XNOR2_X1 U788 ( .A(G131), .B(n741), .ZN(G33) );
  XNOR2_X1 U789 ( .A(n742), .B(G137), .ZN(G39) );
endmodule

