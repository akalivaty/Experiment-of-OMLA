//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT84), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n206), .B(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G36gat), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n213), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n214));
  OR3_X1    g013(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT15), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  XNOR2_X1  g015(.A(G43gat), .B(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(new_n218), .B2(new_n219), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n209), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G229gat), .A2(G233gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT18), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n209), .B(new_n221), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n227), .B(KEYINPUT13), .Z(new_n232));
  AOI22_X1  g031(.A1(new_n228), .A2(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT85), .B1(new_n228), .B2(new_n229), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT12), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n230), .B(new_n233), .C1(new_n235), .C2(new_n240), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(G57gat), .A2(G64gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(G57gat), .A2(G64gat), .ZN(new_n247));
  AND2_X1   g046(.A1(G71gat), .A2(G78gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n246), .B(new_n247), .C1(new_n248), .C2(KEYINPUT9), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT86), .B1(G71gat), .B2(G78gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(G71gat), .A2(G78gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n249), .B(new_n250), .C1(new_n248), .C2(new_n252), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT21), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G231gat), .A2(G233gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G127gat), .B(G155gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT20), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G183gat), .B(G211gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n209), .B1(new_n258), .B2(new_n257), .ZN(new_n267));
  XOR2_X1   g066(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G99gat), .A2(G106gat), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(KEYINPUT8), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G99gat), .B(G106gat), .Z(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(KEYINPUT88), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT88), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n282), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n287), .C1(new_n223), .C2(new_n225), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n283), .ZN(new_n289));
  NAND2_X1  g088(.A1(G232gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n289), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n294), .B(KEYINPUT89), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n291), .A2(KEYINPUT41), .ZN(new_n298));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(KEYINPUT90), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n273), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n284), .A2(new_n286), .B1(new_n254), .B2(new_n255), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n306), .B1(new_n289), .B2(new_n257), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT91), .B1(new_n307), .B2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT91), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n256), .B1(new_n287), .B2(new_n283), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n310), .C1(new_n311), .C2(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n256), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G230gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT92), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n307), .A2(new_n317), .ZN(new_n320));
  XNOR2_X1  g119(.A(G120gat), .B(G148gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G176gat), .B(G204gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n314), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n308), .B2(new_n312), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n320), .B1(new_n326), .B2(new_n317), .ZN(new_n327));
  INV_X1    g126(.A(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n305), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n333), .B(new_n334), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(G169gat), .ZN(new_n340));
  OR2_X1    g139(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT23), .ZN(new_n345));
  INV_X1    g144(.A(G169gat), .ZN(new_n346));
  INV_X1    g145(.A(G176gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  AND2_X1   g151(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(G190gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n338), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n338), .B1(new_n356), .B2(KEYINPUT23), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT65), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT65), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n361), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n352), .A2(new_n351), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT27), .B(G183gat), .ZN(new_n368));
  INV_X1    g167(.A(G190gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT26), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT26), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n344), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n371), .B(new_n351), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n368), .A2(new_n367), .A3(new_n369), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n355), .A2(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n337), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n368), .A2(new_n369), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT28), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n348), .A2(new_n372), .A3(new_n344), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n371), .A2(new_n351), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n381), .A2(new_n377), .A3(new_n382), .A4(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n387), .A2(new_n340), .B1(new_n348), .B2(new_n345), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n359), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT25), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n349), .A2(new_n357), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n364), .B2(new_n363), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n384), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n337), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G204gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G197gat), .ZN(new_n397));
  INV_X1    g196(.A(G197gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G204gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n402));
  OAI21_X1  g201(.A(G218gat), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT68), .B(KEYINPUT22), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G211gat), .B(G218gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n405), .B(new_n408), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n379), .A2(KEYINPUT72), .A3(new_n395), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT71), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n378), .B2(new_n337), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n393), .A2(KEYINPUT71), .A3(new_n394), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n343), .A3(new_n349), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(new_n338), .B1(new_n358), .B2(new_n365), .ZN(new_n416));
  INV_X1    g215(.A(new_n377), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n417), .A2(new_n370), .A3(new_n375), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n412), .A2(new_n413), .B1(new_n337), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n410), .B1(new_n420), .B2(new_n409), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n379), .A2(new_n409), .A3(new_n395), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n336), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n378), .A2(new_n411), .A3(new_n337), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT71), .B1(new_n393), .B2(new_n394), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n379), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n406), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n405), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n422), .A2(new_n423), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n410), .A4(new_n335), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n422), .ZN(new_n436));
  AOI22_X1  g235(.A1(KEYINPUT72), .A2(new_n436), .B1(new_n428), .B2(new_n431), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n433), .A4(new_n335), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G148gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(G141gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(G148gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT2), .ZN(new_n448));
  INV_X1    g247(.A(G155gat), .ZN(new_n449));
  INV_X1    g248(.A(G162gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(G141gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G148gat), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT2), .B1(new_n442), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n449), .A3(new_n450), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n452), .A3(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n447), .A2(new_n454), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  INV_X1    g262(.A(G134gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G127gat), .ZN(new_n465));
  INV_X1    g264(.A(G127gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G134gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G113gat), .B(G120gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n469), .B2(KEYINPUT1), .ZN(new_n470));
  INV_X1    g269(.A(G120gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G113gat), .ZN(new_n472));
  INV_X1    g271(.A(G113gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G120gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G127gat), .B(G134gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT1), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n462), .A2(new_n463), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(G148gat), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n442), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n459), .A2(new_n452), .A3(new_n460), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n442), .A2(new_n456), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n448), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n484), .A2(new_n453), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n470), .A2(new_n478), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT4), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n461), .A2(new_n457), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n483), .A2(new_n442), .B1(new_n452), .B2(new_n451), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT3), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n487), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n444), .A2(new_n445), .A3(new_n441), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n453), .B1(new_n497), .B2(new_n443), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT3), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n500), .A3(new_n479), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT75), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n491), .A2(new_n492), .A3(new_n501), .A4(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n463), .B1(new_n462), .B2(new_n479), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n501), .A2(new_n492), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n462), .B(new_n489), .ZN(new_n512));
  INV_X1    g311(.A(new_n492), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G1gat), .B(G29gat), .Z(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G85gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n515), .B1(new_n505), .B2(new_n510), .ZN(new_n525));
  INV_X1    g324(.A(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n522), .B(new_n515), .C1(new_n505), .C2(new_n510), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n440), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT78), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n397), .A2(new_n399), .ZN(new_n535));
  INV_X1    g334(.A(G218gat), .ZN(new_n536));
  OR2_X1    g335(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(KEYINPUT69), .A2(G211gat), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT22), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT68), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT68), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT22), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n535), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n430), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n405), .A2(new_n408), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n414), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n488), .B1(new_n548), .B2(new_n499), .ZN(new_n549));
  NAND2_X1  g348(.A1(G228gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n488), .B2(new_n499), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n409), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n414), .B1(new_n405), .B2(new_n407), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n545), .A2(new_n406), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n499), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n500), .A2(new_n414), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n558), .A2(new_n462), .B1(new_n559), .B2(new_n431), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n560), .A2(KEYINPUT79), .A3(new_n551), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT29), .B1(new_n545), .B2(new_n406), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n405), .A2(new_n407), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT3), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n565), .A2(new_n488), .B1(new_n552), .B2(new_n409), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n566), .B2(new_n550), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n555), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(G22gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G78gat), .B(G106gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G50gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G22gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(new_n555), .C1(new_n561), .C2(new_n567), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n569), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT79), .B1(new_n560), .B2(new_n551), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(new_n562), .A3(new_n550), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n554), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT81), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT80), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n575), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT81), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n584), .A3(G22gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n574), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n581), .A2(new_n583), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n577), .B1(new_n587), .B2(new_n572), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n440), .A2(new_n532), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n534), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n572), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n576), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n432), .A2(new_n433), .A3(new_n410), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n336), .B1(new_n594), .B2(KEYINPUT37), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n437), .B2(new_n433), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT38), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n529), .A2(new_n530), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n517), .A2(new_n524), .A3(new_n522), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n379), .A2(new_n395), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n431), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n603), .B(KEYINPUT82), .C1(new_n428), .C2(new_n431), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n409), .B1(new_n379), .B2(new_n395), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT82), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n596), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT38), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n336), .C1(KEYINPUT37), .C2(new_n594), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n598), .A2(new_n601), .A3(new_n609), .A4(new_n434), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n512), .B2(new_n492), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n501), .A2(new_n506), .A3(new_n507), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n513), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n615), .B(new_n522), .C1(KEYINPUT39), .C2(new_n614), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n527), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n617), .B2(new_n616), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n439), .A3(new_n435), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n593), .A2(new_n610), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n479), .B1(new_n416), .B2(new_n418), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n384), .B(new_n489), .C1(new_n390), .C2(new_n392), .ZN(new_n623));
  INV_X1    g422(.A(G227gat), .ZN(new_n624));
  INV_X1    g423(.A(G233gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT67), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT34), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G15gat), .B(G43gat), .Z(new_n631));
  XNOR2_X1  g430(.A(G71gat), .B(G99gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n627), .B1(new_n622), .B2(new_n623), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT66), .B(KEYINPUT33), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT32), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n623), .ZN(new_n641));
  AOI221_X4 g440(.A(new_n638), .B1(new_n636), .B2(new_n633), .C1(new_n641), .C2(new_n626), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n630), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n626), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT32), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n635), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n633), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n637), .A2(new_n639), .ZN(new_n648));
  INV_X1    g447(.A(new_n630), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n628), .A2(new_n629), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n643), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n651), .B1(new_n643), .B2(new_n650), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n643), .A2(new_n650), .ZN(new_n657));
  INV_X1    g456(.A(new_n651), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT36), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n591), .A2(new_n621), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT35), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n534), .A2(new_n590), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n653), .A2(new_n654), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n588), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n659), .A2(new_n652), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n593), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n440), .A2(new_n532), .A3(new_n663), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n662), .B1(new_n667), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT83), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT83), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n674), .B(new_n662), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n245), .B(new_n332), .C1(new_n673), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n601), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT93), .B(G1gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT95), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n680), .B(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n440), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n676), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n683), .B1(new_n686), .B2(new_n681), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n686), .A2(KEYINPUT94), .B1(new_n681), .B2(G8gat), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n686), .A2(KEYINPUT94), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(G1325gat));
  INV_X1    g489(.A(G15gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n691), .A3(new_n668), .ZN(new_n692));
  INV_X1    g491(.A(new_n661), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n676), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(new_n691), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n588), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT96), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n304), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n673), .B2(new_n675), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n272), .A2(new_n245), .A3(new_n330), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(G29gat), .A3(new_n532), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT45), .Z(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n672), .A2(new_n706), .A3(new_n304), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n669), .A2(new_n670), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n440), .A2(new_n589), .A3(new_n532), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n589), .B1(new_n440), .B2(new_n532), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT35), .B1(new_n711), .B2(new_n669), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n674), .B1(new_n713), .B2(new_n662), .ZN(new_n714));
  INV_X1    g513(.A(new_n675), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n304), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n707), .B1(new_n716), .B2(KEYINPUT44), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n702), .B(KEYINPUT97), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n532), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n721), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n440), .A2(G36gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n701), .A2(new_n702), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT98), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(new_n684), .A3(new_n719), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n723), .A2(new_n726), .B1(new_n727), .B2(G36gat), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n726), .A2(KEYINPUT99), .A3(new_n723), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT99), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT98), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n725), .B(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(KEYINPUT46), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n728), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT100), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n728), .B(KEYINPUT100), .C1(new_n729), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1329gat));
  INV_X1    g537(.A(new_n720), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n693), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G43gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n703), .A2(G43gat), .A3(new_n665), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT102), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n746));
  INV_X1    g545(.A(new_n744), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n746), .B(new_n747), .C1(new_n740), .C2(G43gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n742), .B(KEYINPUT101), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n740), .B2(G43gat), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n745), .A2(new_n748), .B1(KEYINPUT47), .B2(new_n750), .ZN(G1330gat));
  NAND3_X1  g550(.A1(new_n739), .A2(G50gat), .A3(new_n588), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n703), .A2(new_n593), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(G50gat), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g554(.A1(new_n672), .A2(new_n245), .A3(new_n305), .A4(new_n330), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n601), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n684), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  XNOR2_X1  g561(.A(new_n665), .B(KEYINPUT103), .ZN(new_n763));
  AOI21_X1  g562(.A(G71gat), .B1(new_n756), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n693), .A2(G71gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g566(.A1(new_n756), .A2(new_n588), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT104), .B(G78gat), .Z(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n272), .A2(new_n244), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n672), .A2(new_n304), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n331), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n275), .A3(new_n601), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n771), .A2(new_n330), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n717), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n779), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n673), .A2(new_n675), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n706), .B1(new_n782), .B2(new_n304), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT105), .B(new_n781), .C1(new_n783), .C2(new_n707), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n601), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n777), .B1(new_n786), .B2(new_n275), .ZN(G1336gat));
  AND3_X1   g586(.A1(new_n776), .A2(new_n276), .A3(new_n684), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT107), .B(KEYINPUT52), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n718), .A2(new_n781), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n791), .B2(new_n440), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n780), .A2(new_n684), .A3(new_n784), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(G92gat), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n794), .B2(G92gat), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(new_n788), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(G1337gat));
  INV_X1    g599(.A(G99gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n776), .A2(new_n801), .A3(new_n668), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n785), .A2(new_n693), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n801), .ZN(G1338gat));
  OAI21_X1  g603(.A(G106gat), .B1(new_n791), .B2(new_n593), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n593), .A2(G106gat), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n776), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n785), .A2(new_n588), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n809), .A2(G106gat), .B1(new_n776), .B2(new_n806), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  NAND3_X1  g611(.A1(new_n305), .A2(new_n245), .A3(new_n331), .ZN(new_n813));
  XOR2_X1   g612(.A(KEYINPUT108), .B(KEYINPUT54), .Z(new_n814));
  NAND3_X1  g613(.A1(new_n315), .A2(new_n318), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n326), .B2(new_n317), .ZN(new_n816));
  AOI211_X1 g615(.A(new_n318), .B(new_n325), .C1(new_n308), .C2(new_n312), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n815), .B(new_n328), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n326), .A2(new_n317), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n319), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n326), .A2(new_n317), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n323), .B1(new_n823), .B2(new_n814), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n824), .A3(KEYINPUT55), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(new_n324), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n227), .B1(new_n222), .B2(new_n226), .ZN(new_n827));
  OAI22_X1  g626(.A1(new_n827), .A2(KEYINPUT109), .B1(new_n231), .B2(new_n232), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n239), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT110), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n230), .A2(new_n233), .A3(new_n240), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n239), .C1(new_n828), .C2(new_n829), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n826), .A2(new_n700), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n244), .A3(new_n825), .A4(new_n324), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n831), .A2(new_n330), .A3(new_n832), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n304), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(KEYINPUT111), .A3(new_n838), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n813), .B1(new_n843), .B2(new_n272), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n601), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n666), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n440), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n473), .A3(new_n244), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n844), .A2(new_n593), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT112), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n840), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n700), .A3(new_n842), .ZN(new_n856));
  INV_X1    g655(.A(new_n836), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n272), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n813), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n854), .B(new_n593), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n684), .A2(new_n532), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n668), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(new_n245), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(G113gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n864), .B2(G113gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(G1340gat));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n471), .A3(new_n330), .ZN(new_n869));
  OAI21_X1  g668(.A(G120gat), .B1(new_n863), .B2(new_n331), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n863), .B2(new_n273), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n272), .A2(new_n466), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n848), .B2(new_n873), .ZN(G1342gat));
  NOR4_X1   g673(.A1(new_n846), .A2(G134gat), .A3(new_n684), .A4(new_n700), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n863), .B2(new_n700), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n661), .A2(new_n862), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT115), .Z(new_n883));
  AOI21_X1  g682(.A(new_n304), .B1(new_n837), .B2(new_n838), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n273), .B1(new_n836), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n593), .B1(new_n813), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT116), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n844), .B2(new_n588), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n244), .B(new_n883), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n445), .B2(new_n444), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n845), .A2(new_n588), .A3(new_n661), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n684), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n455), .A3(new_n244), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n880), .B(new_n881), .C1(new_n891), .C2(new_n894), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n879), .A2(new_n891), .A3(KEYINPUT58), .A4(new_n894), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n441), .A3(new_n330), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n888), .A2(new_n889), .ZN(new_n899));
  INV_X1    g698(.A(new_n883), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT59), .B(new_n441), .C1(new_n901), .C2(new_n330), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n844), .A2(KEYINPUT57), .A3(new_n588), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n844), .A2(new_n905), .A3(KEYINPUT57), .A4(new_n588), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n330), .A3(new_n883), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n903), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n898), .B1(new_n902), .B2(new_n911), .ZN(G1345gat));
  AOI21_X1  g711(.A(G155gat), .B1(new_n893), .B2(new_n272), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n272), .A2(G155gat), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT119), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n901), .B2(new_n915), .ZN(G1346gat));
  AOI21_X1  g715(.A(new_n450), .B1(new_n901), .B2(new_n304), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n892), .A2(G162gat), .A3(new_n684), .A4(new_n700), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  AND2_X1   g718(.A1(new_n844), .A2(new_n532), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n684), .A3(new_n666), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(G169gat), .B1(new_n922), .B2(new_n244), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n601), .A2(new_n440), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n763), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n853), .B2(new_n860), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n245), .A2(new_n346), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  AOI21_X1  g727(.A(G176gat), .B1(new_n922), .B2(new_n330), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n331), .A2(new_n387), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n926), .B2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(new_n925), .ZN(new_n932));
  INV_X1    g731(.A(new_n860), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n854), .B1(new_n844), .B2(new_n593), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n272), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n861), .A2(KEYINPUT120), .A3(new_n272), .A4(new_n932), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(G183gat), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n272), .A2(new_n368), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g740(.A1(KEYINPUT121), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G183gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n935), .B2(new_n936), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n945), .A2(new_n938), .B1(new_n922), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(KEYINPUT121), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT60), .B1(new_n946), .B2(KEYINPUT122), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n922), .A2(new_n369), .A3(new_n304), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n926), .A2(new_n304), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  AND4_X1   g751(.A1(KEYINPUT123), .A2(new_n951), .A3(new_n952), .A4(G190gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n369), .B1(new_n954), .B2(KEYINPUT61), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n951), .A2(new_n955), .B1(KEYINPUT123), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n950), .B1(new_n953), .B2(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n909), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n907), .A2(KEYINPUT124), .A3(new_n908), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n661), .A2(new_n924), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n963), .A2(new_n398), .A3(new_n245), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n693), .A2(new_n593), .A3(new_n440), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n920), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n244), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n964), .A2(new_n968), .ZN(G1352gat));
  NAND4_X1  g768(.A1(new_n959), .A2(new_n330), .A3(new_n960), .A4(new_n962), .ZN(new_n970));
  XOR2_X1   g769(.A(KEYINPUT125), .B(G204gat), .Z(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n920), .A2(new_n330), .A3(new_n965), .A4(new_n971), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT62), .Z(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n973), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1353gat));
  NAND3_X1  g779(.A1(new_n909), .A2(new_n272), .A3(new_n962), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(G211gat), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  NAND4_X1  g782(.A1(new_n967), .A2(new_n537), .A3(new_n538), .A4(new_n272), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1354gat));
  OAI21_X1  g784(.A(new_n536), .B1(new_n966), .B2(new_n700), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n304), .A2(G218gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n963), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


