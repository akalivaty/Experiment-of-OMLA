//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XOR2_X1   g020(.A(KEYINPUT64), .B(KEYINPUT1), .Z(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n461), .A2(new_n463), .A3(G137), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(KEYINPUT66), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n472), .B1(G2105), .B2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n461), .A2(new_n463), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n477), .A2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(KEYINPUT68), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n487), .A2(new_n461), .A3(new_n463), .A4(new_n464), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .A3(new_n464), .A4(new_n487), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n461), .A2(new_n463), .A3(G126), .A4(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n497), .A3(G2104), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n493), .B2(new_n498), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n490), .B(new_n492), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT69), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n503), .A2(new_n510), .B1(new_n511), .B2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT72), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT70), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n522), .A2(new_n525), .A3(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n512), .A2(G89), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n509), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n518), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n526), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(new_n512), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n503), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G171));
  INV_X1    g115(.A(new_n536), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n541), .A2(G81), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n503), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  AOI22_X1  g128(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n503), .B1(new_n555), .B2(new_n536), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT75), .A2(G53), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n522), .A2(new_n525), .A3(G543), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n505), .B1(new_n512), .B2(KEYINPUT70), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n561), .A2(new_n562), .A3(new_n522), .A4(new_n558), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n560), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n564), .B1(new_n560), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n557), .B1(new_n565), .B2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  XNOR2_X1  g143(.A(new_n532), .B(KEYINPUT77), .ZN(G286));
  NAND3_X1  g144(.A1(new_n509), .A2(G87), .A3(new_n512), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n522), .A2(new_n525), .A3(G49), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n503), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n509), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n513), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n503), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT78), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n541), .A2(G85), .B1(new_n526), .B2(G47), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(new_n506), .A2(new_n508), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n587), .A2(G92), .A3(new_n588), .A4(new_n512), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .A4(new_n512), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n561), .A2(G54), .A3(new_n522), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n503), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT79), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n587), .A2(new_n588), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n526), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n591), .A2(new_n592), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(G868), .B1(new_n597), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g182(.A(new_n606), .B1(G868), .B2(G171), .ZN(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  NAND2_X1  g185(.A1(new_n597), .A2(new_n605), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  AOI21_X1  g188(.A(KEYINPUT80), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT80), .ZN(new_n615));
  AOI211_X1 g190(.A(new_n615), .B(G559), .C1(new_n597), .C2(new_n605), .ZN(new_n616));
  OAI21_X1  g191(.A(G868), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n619));
  XNOR2_X1  g194(.A(G323), .B(new_n619), .ZN(G282));
  NAND2_X1  g195(.A1(new_n478), .A2(G2104), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n623));
  AOI22_X1  g198(.A1(new_n622), .A2(new_n623), .B1(KEYINPUT82), .B2(G2100), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  OR3_X1    g200(.A1(new_n625), .A2(KEYINPUT82), .A3(G2100), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(KEYINPUT82), .B2(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n478), .A2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n480), .A2(G123), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n630), .A2(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n630), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n626), .A2(new_n627), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n641), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  AOI21_X1  g233(.A(KEYINPUT18), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(new_n661), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  INV_X1    g248(.A(new_n671), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  MUX2_X1   g251(.A(new_n676), .B(new_n675), .S(new_n668), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n682), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G23), .B(G288), .S(G16), .Z(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n580), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  NOR3_X1   g277(.A1(new_n694), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT34), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(G290), .A2(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n695), .A2(G24), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT88), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(G1986), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n478), .A2(G131), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n480), .A2(G119), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n464), .A2(G107), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n713), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT87), .B(G29), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G25), .B(new_n717), .S(new_n719), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n720), .B(new_n721), .Z(new_n722));
  AND3_X1   g297(.A1(new_n711), .A2(new_n712), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n703), .A2(new_n704), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n705), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT36), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n695), .A2(G20), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  INV_X1    g303(.A(G299), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n695), .ZN(new_n730));
  INV_X1    g305(.A(G1956), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G19), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n733), .A2(KEYINPUT90), .A3(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(new_n733), .B2(G16), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n734), .B(new_n735), .C1(new_n547), .C2(new_n695), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n719), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n719), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT29), .Z(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT100), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n718), .A2(G26), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT28), .Z(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT92), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G128), .B2(new_n480), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n478), .A2(G140), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT91), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n745), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT93), .B(G2067), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n742), .A2(new_n743), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n740), .A2(KEYINPUT100), .A3(new_n741), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT89), .B(G1348), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G4), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n611), .B2(G16), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n756), .B(new_n757), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n737), .B(new_n762), .C1(new_n759), .C2(new_n761), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT25), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G139), .B2(new_n478), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n464), .B2(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G33), .B(new_n768), .S(G29), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  INV_X1    g347(.A(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(KEYINPUT30), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n772), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n770), .B(new_n776), .C1(new_n635), .C2(new_n718), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n769), .A2(G2072), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n719), .A2(G27), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n719), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT24), .B(G34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n718), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT94), .Z(new_n787));
  INV_X1    g362(.A(G160), .ZN(new_n788));
  INV_X1    g363(.A(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n779), .B(new_n783), .C1(new_n784), .C2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT98), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G301), .B2(new_n695), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n695), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n695), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n792), .A2(new_n795), .B1(new_n797), .B2(G1966), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G1966), .B2(new_n797), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n789), .A2(G32), .ZN(new_n800));
  AOI22_X1  g375(.A1(G129), .A2(new_n480), .B1(new_n478), .B2(G141), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT95), .B(KEYINPUT26), .Z(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n466), .A2(G105), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT96), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n800), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT27), .B(G1996), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n790), .A2(new_n784), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n795), .A2(new_n792), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n791), .A2(new_n799), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT99), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n726), .A2(new_n732), .A3(new_n763), .A4(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  AOI22_X1  g393(.A1(new_n541), .A2(G93), .B1(new_n526), .B2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n821));
  OAI21_X1  g396(.A(G651), .B1(new_n820), .B2(KEYINPUT101), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n611), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT38), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n545), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n547), .A2(new_n823), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n830), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n826), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n828), .B1(new_n836), .B2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(G160), .B(G162), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n635), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n622), .B(new_n717), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n478), .A2(G142), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n480), .A2(G130), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n845));
  INV_X1    g420(.A(G118), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n844), .A2(new_n845), .B1(new_n846), .B2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(new_n844), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n842), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n841), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n807), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n807), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n752), .B(new_n768), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(new_n498), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n493), .A2(new_n498), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n859), .A2(KEYINPUT103), .A3(new_n490), .A4(new_n492), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n853), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n840), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(new_n840), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n869), .A3(new_n864), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n874), .A2(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n602), .A2(new_n604), .ZN(new_n876));
  XOR2_X1   g451(.A(G299), .B(new_n876), .Z(new_n877));
  INV_X1    g452(.A(KEYINPUT41), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT41), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n614), .A2(new_n616), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n833), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n833), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n883), .B1(new_n888), .B2(new_n887), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n875), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G290), .B(G305), .ZN(new_n893));
  XNOR2_X1  g468(.A(G166), .B(G288), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n895), .B1(KEYINPUT106), .B2(new_n874), .ZN(new_n896));
  INV_X1    g471(.A(new_n891), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n889), .C1(KEYINPUT106), .C2(new_n874), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n892), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n892), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n825), .A2(G868), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G295));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(G331));
  XOR2_X1   g479(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NOR2_X1   g481(.A1(G286), .A2(G301), .ZN(new_n907));
  NOR2_X1   g482(.A1(G171), .A2(G168), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n833), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n831), .B(new_n832), .C1(new_n907), .C2(new_n908), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n910), .A2(new_n877), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n885), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n895), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n885), .A2(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n910), .A2(new_n877), .A3(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n895), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n906), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n910), .A2(new_n922), .A3(new_n911), .A4(new_n877), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n911), .A2(new_n910), .B1(new_n884), .B2(new_n879), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n895), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n917), .A2(new_n915), .A3(new_n918), .ZN(new_n927));
  AND4_X1   g502(.A1(new_n906), .A2(new_n926), .A3(new_n927), .A4(new_n871), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n905), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n916), .A2(new_n906), .A3(new_n920), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n926), .A2(new_n871), .A3(new_n927), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n930), .B(KEYINPUT44), .C1(new_n931), .C2(new_n906), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(G397));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n861), .B2(G1384), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n475), .A2(G2105), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n470), .A2(new_n936), .A3(G40), .A4(new_n471), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n807), .A2(G1996), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n752), .B(G2067), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n807), .A2(G1996), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n717), .A2(new_n721), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n721), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G290), .B(G1986), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n937), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n855), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n501), .B2(new_n950), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n952), .A2(new_n953), .A3(G2084), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n855), .A2(new_n950), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n937), .B1(new_n955), .B2(new_n934), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n957));
  AOI21_X1  g532(.A(G1966), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT120), .B(G8), .C1(new_n954), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G8), .ZN(new_n960));
  NOR2_X1   g535(.A1(G168), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT51), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n957), .ZN(new_n964));
  INV_X1    g539(.A(G1966), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n501), .A2(new_n950), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(new_n784), .A3(new_n948), .A4(new_n951), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT120), .B1(new_n970), .B2(G8), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT121), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(G8), .B1(new_n954), .B2(new_n958), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT120), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT121), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n959), .A4(new_n962), .ZN(new_n977));
  OAI211_X1 g552(.A(KEYINPUT51), .B(G8), .C1(new_n970), .C2(new_n532), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n970), .A2(new_n961), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT109), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(G166), .B2(new_n960), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND4_X1  g562(.A1(G303), .A2(new_n987), .A3(KEYINPUT55), .A4(G8), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n937), .B1(new_n967), .B2(new_n934), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n860), .A4(new_n950), .ZN(new_n992));
  AOI21_X1  g567(.A(G1971), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n948), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n501), .A2(new_n949), .A3(new_n950), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n858), .A2(KEYINPUT67), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n490), .A2(new_n492), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n949), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n995), .B1(new_n997), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n993), .B1(new_n741), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n990), .B1(new_n1007), .B2(new_n960), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n948), .B(new_n951), .C1(new_n1003), .C2(new_n949), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  OAI211_X1 g585(.A(G8), .B(new_n989), .C1(new_n993), .C2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n967), .A2(new_n934), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1014), .A2(new_n948), .A3(new_n992), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1015), .A2(G1971), .B1(G2090), .B2(new_n1009), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(KEYINPUT110), .A3(G8), .A4(new_n989), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n574), .A2(new_n570), .A3(G1976), .A4(new_n571), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n955), .B2(new_n937), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT113), .B(G1976), .Z(new_n1025));
  INV_X1    g600(.A(new_n574), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n572), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(KEYINPUT114), .A3(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1024), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n577), .A2(new_n579), .A3(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(G1981), .B1(new_n577), .B2(new_n579), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(KEYINPUT49), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(new_n1034), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1023), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1043), .B(KEYINPUT52), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n955), .A2(new_n937), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n1020), .A3(G8), .A4(new_n1021), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1047), .B2(KEYINPUT52), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1033), .B(new_n1042), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1014), .A2(new_n782), .A3(new_n948), .A4(new_n992), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n964), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT123), .B(G1961), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n1009), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G171), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AND4_X1   g635(.A1(new_n1008), .A2(new_n1018), .A3(new_n1050), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n982), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n982), .B2(new_n1061), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G288), .A2(G1976), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1042), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1041), .B1(new_n1068), .B2(new_n1034), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1018), .B2(new_n1049), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1049), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n973), .A2(G286), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1008), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n973), .A2(new_n1074), .A3(G286), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1016), .A2(G8), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1071), .B(new_n1076), .C1(new_n989), .C2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1070), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n560), .A2(new_n563), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1080), .A2(new_n556), .A3(KEYINPUT57), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n991), .A2(new_n992), .A3(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1082), .B(new_n1084), .C1(new_n1006), .C2(G1956), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1006), .B2(G1956), .ZN(new_n1087));
  AND2_X1   g662(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1081), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n955), .A2(new_n937), .A3(G2067), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1009), .B2(new_n758), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n611), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1086), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n597), .A2(new_n605), .A3(KEYINPUT119), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT119), .B1(new_n597), .B2(new_n605), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1091), .B2(KEYINPUT60), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n758), .B1(new_n952), .B2(new_n953), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1090), .ZN(new_n1099));
  AND4_X1   g674(.A1(KEYINPUT60), .A2(new_n1096), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1095), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(new_n995), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1004), .B1(new_n1003), .B2(new_n949), .ZN(new_n1106));
  AND4_X1   g681(.A1(new_n1004), .A2(new_n501), .A3(new_n949), .A4(new_n950), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n731), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1082), .B1(new_n1109), .B2(new_n1084), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1104), .B1(new_n1110), .B2(new_n1086), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1089), .A2(KEYINPUT61), .A3(new_n1085), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1103), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1996), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1014), .A2(new_n1114), .A3(new_n948), .A4(new_n992), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n991), .A2(KEYINPUT116), .A3(new_n1114), .A4(new_n992), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(G1341), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1046), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n547), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1122), .B2(new_n547), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1113), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1094), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n473), .A2(new_n474), .ZN(new_n1131));
  OAI21_X1  g706(.A(G2105), .B1(new_n1131), .B2(KEYINPUT124), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(KEYINPUT124), .B2(new_n1131), .ZN(new_n1133));
  INV_X1    g708(.A(G40), .ZN(new_n1134));
  NOR4_X1   g709(.A1(new_n1133), .A2(new_n1134), .A3(new_n472), .A4(new_n1054), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1135), .A2(new_n992), .A3(new_n935), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1053), .A2(new_n1136), .A3(new_n1057), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G171), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(KEYINPUT54), .C1(G171), .C2(new_n1058), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1071), .A2(new_n1139), .A3(new_n1008), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n979), .A2(new_n981), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1053), .A2(new_n1136), .A3(G301), .A4(new_n1057), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1059), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1140), .A2(new_n1141), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1079), .B1(new_n1130), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n947), .B1(new_n1066), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n938), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1151), .A2(G1986), .A3(G290), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1153), .A2(KEYINPUT48), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1153), .A2(KEYINPUT48), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1154), .B(new_n1155), .C1(new_n938), .C2(new_n945), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n938), .B1(new_n940), .B2(new_n807), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT46), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1151), .B2(G1996), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n938), .A2(KEYINPUT46), .A3(new_n1114), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  XOR2_X1   g737(.A(new_n943), .B(KEYINPUT127), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n942), .A2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n752), .A2(G2067), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1151), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1156), .A2(new_n1162), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1150), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(new_n921), .A2(new_n928), .ZN(new_n1170));
  OAI21_X1  g744(.A(G319), .B1(new_n651), .B2(new_n652), .ZN(new_n1171));
  NOR2_X1   g745(.A1(G227), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n872), .A2(new_n690), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1170), .A2(new_n1173), .ZN(G308));
  AND2_X1   g748(.A1(new_n690), .A2(new_n1172), .ZN(new_n1175));
  OAI211_X1 g749(.A(new_n1175), .B(new_n872), .C1(new_n921), .C2(new_n928), .ZN(G225));
endmodule


