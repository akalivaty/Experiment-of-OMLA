

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761;

  AND2_X1 U368 ( .A1(n361), .A2(n431), .ZN(n651) );
  OR2_X1 U369 ( .A1(n645), .A2(G902), .ZN(n445) );
  XNOR2_X1 U370 ( .A(n482), .B(G134), .ZN(n505) );
  BUF_X1 U371 ( .A(G128), .Z(n345) );
  XNOR2_X1 U372 ( .A(n740), .B(n446), .ZN(n533) );
  XNOR2_X1 U373 ( .A(n447), .B(KEYINPUT4), .ZN(n507) );
  INV_X2 U374 ( .A(G953), .ZN(n752) );
  AND2_X2 U375 ( .A1(n425), .A2(n424), .ZN(n423) );
  AND2_X2 U376 ( .A1(n442), .A2(n441), .ZN(n387) );
  NOR2_X2 U377 ( .A1(n705), .A2(n704), .ZN(n546) );
  XNOR2_X2 U378 ( .A(n590), .B(KEYINPUT1), .ZN(n705) );
  AND2_X2 U379 ( .A1(n432), .A2(n367), .ZN(n429) );
  XNOR2_X1 U380 ( .A(n507), .B(KEYINPUT72), .ZN(n446) );
  XOR2_X1 U381 ( .A(n506), .B(n505), .Z(n749) );
  AND2_X2 U382 ( .A1(n637), .A2(KEYINPUT81), .ZN(n638) );
  XOR2_X2 U383 ( .A(n398), .B(KEYINPUT38), .Z(n697) );
  NOR2_X1 U384 ( .A1(n727), .A2(n550), .ZN(n390) );
  INV_X1 U385 ( .A(KEYINPUT33), .ZN(n346) );
  XNOR2_X1 U386 ( .A(n624), .B(n623), .ZN(n634) );
  NAND2_X1 U387 ( .A1(n538), .A2(n450), .ZN(n449) );
  XNOR2_X1 U388 ( .A(n358), .B(n503), .ZN(n361) );
  OR2_X1 U389 ( .A1(n550), .A2(n549), .ZN(n675) );
  XNOR2_X1 U390 ( .A(n347), .B(n346), .ZN(n727) );
  NAND2_X1 U391 ( .A1(n546), .A2(n610), .ZN(n347) );
  XNOR2_X1 U392 ( .A(n421), .B(n368), .ZN(n494) );
  INV_X1 U393 ( .A(n502), .ZN(n350) );
  XNOR2_X1 U394 ( .A(G146), .B(n749), .ZN(n535) );
  XNOR2_X1 U395 ( .A(n479), .B(G113), .ZN(n480) );
  XOR2_X1 U396 ( .A(n481), .B(KEYINPUT73), .Z(n369) );
  INV_X1 U397 ( .A(n374), .ZN(n348) );
  XOR2_X1 U398 ( .A(G137), .B(KEYINPUT68), .Z(n530) );
  XNOR2_X1 U399 ( .A(G140), .B(KEYINPUT10), .ZN(n452) );
  XNOR2_X2 U400 ( .A(G143), .B(G128), .ZN(n482) );
  XNOR2_X2 U401 ( .A(n349), .B(n348), .ZN(n395) );
  NAND2_X1 U402 ( .A1(n351), .A2(n350), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n613), .B(n352), .ZN(n351) );
  INV_X1 U404 ( .A(n373), .ZN(n352) );
  XNOR2_X2 U405 ( .A(n420), .B(KEYINPUT84), .ZN(n613) );
  XNOR2_X2 U406 ( .A(n353), .B(n480), .ZN(n362) );
  XNOR2_X2 U407 ( .A(n448), .B(G119), .ZN(n353) );
  INV_X2 U408 ( .A(n589), .ZN(n695) );
  NOR2_X1 U409 ( .A1(n734), .A2(n751), .ZN(n691) );
  AND2_X2 U410 ( .A1(n664), .A2(n649), .ZN(n354) );
  XNOR2_X2 U411 ( .A(n449), .B(KEYINPUT32), .ZN(n664) );
  NAND2_X1 U412 ( .A1(n387), .A2(n386), .ZN(n355) );
  NAND2_X1 U413 ( .A1(n387), .A2(n386), .ZN(n389) );
  NOR2_X2 U414 ( .A1(n734), .A2(n751), .ZN(n356) );
  NOR2_X1 U415 ( .A1(n734), .A2(n751), .ZN(n357) );
  BUF_X1 U416 ( .A(n504), .Z(n358) );
  NOR2_X1 U417 ( .A1(n360), .A2(n502), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n613), .B(n373), .ZN(n360) );
  NOR2_X2 U419 ( .A1(n638), .A2(n437), .ZN(n436) );
  XNOR2_X2 U420 ( .A(n562), .B(n561), .ZN(n734) );
  XNOR2_X2 U421 ( .A(n552), .B(n551), .ZN(n682) );
  OR2_X2 U422 ( .A1(n554), .A2(n553), .ZN(n552) );
  XNOR2_X1 U423 ( .A(n504), .B(n503), .ZN(n538) );
  NAND2_X1 U424 ( .A1(n362), .A2(n369), .ZN(n365) );
  NAND2_X1 U425 ( .A1(n363), .A2(n364), .ZN(n366) );
  NAND2_X1 U426 ( .A1(n366), .A2(n365), .ZN(n742) );
  INV_X1 U427 ( .A(n362), .ZN(n363) );
  INV_X1 U428 ( .A(n369), .ZN(n364) );
  INV_X1 U429 ( .A(n651), .ZN(n430) );
  INV_X1 U430 ( .A(KEYINPUT103), .ZN(n433) );
  NAND2_X1 U431 ( .A1(n389), .A2(n675), .ZN(n385) );
  NOR2_X1 U432 ( .A1(G953), .A2(G237), .ZN(n510) );
  XNOR2_X1 U433 ( .A(n390), .B(KEYINPUT34), .ZN(n541) );
  NAND2_X1 U434 ( .A1(n427), .A2(n556), .ZN(n424) );
  INV_X1 U435 ( .A(KEYINPUT83), .ZN(n388) );
  XNOR2_X1 U436 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n485) );
  NOR2_X1 U437 ( .A1(n501), .A2(n567), .ZN(n502) );
  XNOR2_X1 U438 ( .A(KEYINPUT16), .B(G122), .ZN(n481) );
  INV_X1 U439 ( .A(G107), .ZN(n489) );
  XOR2_X1 U440 ( .A(G104), .B(G110), .Z(n490) );
  XNOR2_X1 U441 ( .A(n517), .B(KEYINPUT71), .ZN(n403) );
  XNOR2_X1 U442 ( .A(G119), .B(KEYINPUT23), .ZN(n517) );
  XOR2_X1 U443 ( .A(G122), .B(KEYINPUT7), .Z(n469) );
  XNOR2_X1 U444 ( .A(n463), .B(n462), .ZN(n654) );
  XNOR2_X1 U445 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U446 ( .A(G469), .ZN(n444) );
  XNOR2_X1 U447 ( .A(KEYINPUT15), .B(G902), .ZN(n635) );
  XOR2_X1 U448 ( .A(KEYINPUT5), .B(KEYINPUT75), .Z(n512) );
  XNOR2_X1 U449 ( .A(KEYINPUT67), .B(G131), .ZN(n506) );
  XNOR2_X1 U450 ( .A(KEYINPUT98), .B(KEYINPUT11), .ZN(n453) );
  XOR2_X1 U451 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n454) );
  XNOR2_X1 U452 ( .A(G143), .B(G113), .ZN(n458) );
  XOR2_X1 U453 ( .A(G122), .B(G104), .Z(n459) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n495) );
  XOR2_X1 U455 ( .A(KEYINPUT89), .B(KEYINPUT14), .Z(n496) );
  INV_X1 U456 ( .A(G237), .ZN(n491) );
  XNOR2_X1 U457 ( .A(n399), .B(n533), .ZN(n656) );
  XNOR2_X1 U458 ( .A(n742), .B(n488), .ZN(n399) );
  NAND2_X1 U459 ( .A1(n493), .A2(G214), .ZN(n696) );
  AND2_X1 U460 ( .A1(n400), .A2(n580), .ZN(n581) );
  XNOR2_X1 U461 ( .A(n401), .B(n376), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n374), .B(KEYINPUT93), .ZN(n391) );
  XNOR2_X1 U463 ( .A(n402), .B(n372), .ZN(n524) );
  XNOR2_X1 U464 ( .A(n521), .B(n403), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n472), .B(n405), .ZN(n640) );
  XNOR2_X1 U466 ( .A(n473), .B(n471), .ZN(n405) );
  NOR2_X1 U467 ( .A1(n371), .A2(n610), .ZN(n450) );
  NAND2_X1 U468 ( .A1(n440), .A2(n439), .ZN(n386) );
  NOR2_X1 U469 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U470 ( .A1(n610), .A2(n555), .ZN(n431) );
  INV_X1 U471 ( .A(KEYINPUT60), .ZN(n407) );
  INV_X1 U472 ( .A(KEYINPUT56), .ZN(n410) );
  AND2_X1 U473 ( .A1(n430), .A2(KEYINPUT82), .ZN(n367) );
  XOR2_X1 U474 ( .A(n492), .B(KEYINPUT88), .Z(n368) );
  XOR2_X1 U475 ( .A(n478), .B(KEYINPUT104), .Z(n370) );
  NAND2_X1 U476 ( .A1(n576), .A2(n626), .ZN(n371) );
  XOR2_X1 U477 ( .A(n519), .B(n518), .Z(n372) );
  XOR2_X1 U478 ( .A(KEYINPUT64), .B(KEYINPUT19), .Z(n373) );
  XOR2_X1 U479 ( .A(KEYINPUT65), .B(KEYINPUT0), .Z(n374) );
  XOR2_X1 U480 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n375) );
  XOR2_X1 U481 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n376) );
  XOR2_X1 U482 ( .A(n645), .B(n644), .Z(n377) );
  XOR2_X1 U483 ( .A(n657), .B(n660), .Z(n378) );
  XNOR2_X1 U484 ( .A(KEYINPUT122), .B(n640), .ZN(n379) );
  XNOR2_X1 U485 ( .A(KEYINPUT62), .B(n662), .ZN(n380) );
  XOR2_X1 U486 ( .A(n654), .B(KEYINPUT59), .Z(n381) );
  NOR2_X1 U487 ( .A1(KEYINPUT81), .A2(n635), .ZN(n382) );
  NAND2_X1 U488 ( .A1(n636), .A2(KEYINPUT2), .ZN(n383) );
  INV_X1 U489 ( .A(n670), .ZN(n418) );
  XOR2_X1 U490 ( .A(KEYINPUT85), .B(KEYINPUT63), .Z(n384) );
  NAND2_X1 U491 ( .A1(n385), .A2(n589), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n354), .B(n388), .ZN(n558) );
  NOR2_X1 U493 ( .A1(n355), .A2(n686), .ZN(n687) );
  NOR2_X1 U494 ( .A1(n355), .A2(n674), .ZN(n652) );
  XNOR2_X1 U495 ( .A(n359), .B(n391), .ZN(n550) );
  NAND2_X1 U496 ( .A1(n432), .A2(n430), .ZN(n427) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n432) );
  BUF_X1 U498 ( .A(n742), .Z(n392) );
  XNOR2_X1 U499 ( .A(n534), .B(n535), .ZN(n645) );
  INV_X1 U500 ( .A(n710), .ZN(n393) );
  XNOR2_X2 U501 ( .A(n545), .B(n544), .ZN(n710) );
  INV_X1 U502 ( .A(n557), .ZN(n394) );
  BUF_X1 U503 ( .A(n693), .Z(n396) );
  NAND2_X1 U504 ( .A1(n354), .A2(n653), .ZN(n397) );
  BUF_X1 U505 ( .A(n494), .Z(n398) );
  NAND2_X1 U506 ( .A1(n612), .A2(n393), .ZN(n401) );
  NOR2_X2 U507 ( .A1(n577), .A2(n578), .ZN(n612) );
  NAND2_X1 U508 ( .A1(n656), .A2(n635), .ZN(n421) );
  NAND2_X1 U509 ( .A1(n404), .A2(n622), .ZN(n624) );
  NOR2_X1 U510 ( .A1(n621), .A2(n620), .ZN(n404) );
  OR2_X2 U511 ( .A1(n682), .A2(n679), .ZN(n589) );
  NAND2_X1 U512 ( .A1(n423), .A2(n406), .ZN(n426) );
  NAND2_X1 U513 ( .A1(n422), .A2(n429), .ZN(n406) );
  XNOR2_X1 U514 ( .A(n408), .B(n407), .ZN(G60) );
  NAND2_X1 U515 ( .A1(n414), .A2(n418), .ZN(n408) );
  XNOR2_X1 U516 ( .A(n409), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U517 ( .A1(n415), .A2(n418), .ZN(n409) );
  XNOR2_X1 U518 ( .A(n411), .B(n410), .ZN(G51) );
  NAND2_X1 U519 ( .A1(n416), .A2(n418), .ZN(n411) );
  XNOR2_X1 U520 ( .A(n412), .B(KEYINPUT123), .ZN(G63) );
  NAND2_X1 U521 ( .A1(n417), .A2(n418), .ZN(n412) );
  XNOR2_X1 U522 ( .A(n413), .B(n384), .ZN(G57) );
  NAND2_X1 U523 ( .A1(n419), .A2(n418), .ZN(n413) );
  NAND2_X1 U524 ( .A1(n438), .A2(n383), .ZN(n437) );
  XNOR2_X1 U525 ( .A(n655), .B(n381), .ZN(n414) );
  XNOR2_X1 U526 ( .A(n646), .B(n377), .ZN(n415) );
  XNOR2_X1 U527 ( .A(n661), .B(n378), .ZN(n416) );
  XNOR2_X1 U528 ( .A(n641), .B(n379), .ZN(n417) );
  XNOR2_X1 U529 ( .A(n663), .B(n380), .ZN(n419) );
  NAND2_X1 U530 ( .A1(n494), .A2(n696), .ZN(n420) );
  NAND2_X1 U531 ( .A1(n397), .A2(KEYINPUT44), .ZN(n422) );
  NAND2_X1 U532 ( .A1(n428), .A2(n443), .ZN(n425) );
  NAND2_X1 U533 ( .A1(n426), .A2(n560), .ZN(n562) );
  NAND2_X1 U534 ( .A1(n354), .A2(n653), .ZN(n428) );
  NOR2_X4 U535 ( .A1(n436), .A2(n693), .ZN(n665) );
  XNOR2_X2 U536 ( .A(n435), .B(n639), .ZN(n693) );
  NAND2_X1 U537 ( .A1(n691), .A2(KEYINPUT2), .ZN(n435) );
  NAND2_X1 U538 ( .A1(n357), .A2(n382), .ZN(n438) );
  NOR2_X1 U539 ( .A1(n715), .A2(n375), .ZN(n439) );
  INV_X1 U540 ( .A(n547), .ZN(n440) );
  NAND2_X1 U541 ( .A1(n715), .A2(n375), .ZN(n441) );
  NAND2_X1 U542 ( .A1(n547), .A2(n375), .ZN(n442) );
  AND2_X1 U543 ( .A1(n556), .A2(KEYINPUT44), .ZN(n443) );
  XNOR2_X2 U544 ( .A(n445), .B(n444), .ZN(n590) );
  XNOR2_X2 U545 ( .A(G101), .B(KEYINPUT66), .ZN(n447) );
  XNOR2_X2 U546 ( .A(G116), .B(KEYINPUT3), .ZN(n448) );
  XOR2_X1 U547 ( .A(n532), .B(n531), .Z(n451) );
  INV_X1 U548 ( .A(KEYINPUT78), .ZN(n601) );
  INV_X1 U549 ( .A(KEYINPUT79), .ZN(n608) );
  XNOR2_X1 U550 ( .A(n609), .B(n608), .ZN(n621) );
  XNOR2_X1 U551 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U552 ( .A(n451), .B(n533), .ZN(n534) );
  INV_X1 U553 ( .A(KEYINPUT35), .ZN(n542) );
  INV_X1 U554 ( .A(KEYINPUT107), .ZN(n598) );
  XNOR2_X1 U555 ( .A(n599), .B(n598), .ZN(n760) );
  XNOR2_X2 U556 ( .A(G146), .B(G125), .ZN(n483) );
  XOR2_X1 U557 ( .A(n452), .B(n483), .Z(n522) );
  XNOR2_X1 U558 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U559 ( .A(n522), .B(n455), .Z(n457) );
  NAND2_X1 U560 ( .A1(G214), .A2(n510), .ZN(n456) );
  XNOR2_X1 U561 ( .A(n457), .B(n456), .ZN(n463) );
  XOR2_X1 U562 ( .A(n459), .B(n458), .Z(n461) );
  XNOR2_X1 U563 ( .A(KEYINPUT12), .B(n506), .ZN(n460) );
  INV_X1 U564 ( .A(G902), .ZN(n525) );
  NAND2_X1 U565 ( .A1(n654), .A2(n525), .ZN(n465) );
  XNOR2_X1 U566 ( .A(KEYINPUT13), .B(G475), .ZN(n464) );
  XNOR2_X2 U567 ( .A(n465), .B(n464), .ZN(n592) );
  XOR2_X1 U568 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n467) );
  NAND2_X1 U569 ( .A1(G234), .A2(n752), .ZN(n466) );
  XNOR2_X1 U570 ( .A(n467), .B(n466), .ZN(n520) );
  NAND2_X1 U571 ( .A1(G217), .A2(n520), .ZN(n468) );
  XNOR2_X1 U572 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U573 ( .A(n470), .B(KEYINPUT9), .Z(n472) );
  XNOR2_X1 U574 ( .A(G116), .B(G107), .ZN(n471) );
  INV_X1 U575 ( .A(n505), .ZN(n473) );
  NAND2_X1 U576 ( .A1(n640), .A2(n525), .ZN(n475) );
  XOR2_X1 U577 ( .A(KEYINPUT101), .B(G478), .Z(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n553) );
  INV_X1 U579 ( .A(n553), .ZN(n591) );
  AND2_X1 U580 ( .A1(n592), .A2(n591), .ZN(n698) );
  NAND2_X1 U581 ( .A1(n635), .A2(G234), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n476), .B(KEYINPUT20), .ZN(n526) );
  NAND2_X1 U583 ( .A1(G221), .A2(n526), .ZN(n477) );
  XOR2_X1 U584 ( .A(KEYINPUT21), .B(n477), .Z(n707) );
  NAND2_X1 U585 ( .A1(n698), .A2(n707), .ZN(n478) );
  INV_X1 U586 ( .A(KEYINPUT70), .ZN(n479) );
  XNOR2_X1 U587 ( .A(n483), .B(n482), .ZN(n487) );
  NAND2_X1 U588 ( .A1(n752), .A2(G224), .ZN(n484) );
  XNOR2_X1 U589 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U590 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n490), .B(n489), .ZN(n740) );
  NAND2_X1 U592 ( .A1(n525), .A2(n491), .ZN(n493) );
  NAND2_X1 U593 ( .A1(n493), .A2(G210), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U595 ( .A(KEYINPUT74), .B(n497), .ZN(n500) );
  NAND2_X1 U596 ( .A1(n500), .A2(G902), .ZN(n498) );
  XOR2_X1 U597 ( .A(n498), .B(KEYINPUT91), .Z(n563) );
  XOR2_X1 U598 ( .A(G898), .B(KEYINPUT90), .Z(n737) );
  NAND2_X1 U599 ( .A1(G953), .A2(n737), .ZN(n744) );
  NOR2_X1 U600 ( .A1(n563), .A2(n744), .ZN(n499) );
  XNOR2_X1 U601 ( .A(n499), .B(KEYINPUT92), .ZN(n501) );
  NAND2_X1 U602 ( .A1(G952), .A2(n500), .ZN(n724) );
  NOR2_X1 U603 ( .A1(n724), .A2(G953), .ZN(n567) );
  NAND2_X1 U604 ( .A1(n395), .A2(n370), .ZN(n504) );
  INV_X1 U605 ( .A(KEYINPUT22), .ZN(n503) );
  XOR2_X1 U606 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n509) );
  XNOR2_X1 U607 ( .A(n507), .B(G137), .ZN(n508) );
  XNOR2_X1 U608 ( .A(n509), .B(n508), .ZN(n515) );
  NAND2_X1 U609 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U611 ( .A(n362), .B(n513), .ZN(n514) );
  XNOR2_X1 U612 ( .A(n535), .B(n516), .ZN(n662) );
  NAND2_X1 U613 ( .A1(n662), .A2(n525), .ZN(n545) );
  INV_X1 U614 ( .A(G472), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n710), .B(KEYINPUT6), .ZN(n610) );
  XOR2_X1 U616 ( .A(KEYINPUT24), .B(KEYINPUT77), .Z(n518) );
  XNOR2_X1 U617 ( .A(n345), .B(G110), .ZN(n519) );
  NAND2_X1 U618 ( .A1(n520), .A2(G221), .ZN(n521) );
  INV_X1 U619 ( .A(n522), .ZN(n523) );
  XNOR2_X1 U620 ( .A(n530), .B(n523), .ZN(n748) );
  XNOR2_X1 U621 ( .A(n524), .B(n748), .ZN(n667) );
  NAND2_X1 U622 ( .A1(n667), .A2(n525), .ZN(n529) );
  NAND2_X1 U623 ( .A1(n526), .A2(G217), .ZN(n527) );
  XNOR2_X1 U624 ( .A(n527), .B(KEYINPUT25), .ZN(n528) );
  XNOR2_X1 U625 ( .A(n529), .B(n528), .ZN(n576) );
  XOR2_X1 U626 ( .A(n530), .B(G140), .Z(n532) );
  NAND2_X1 U627 ( .A1(G227), .A2(n752), .ZN(n531) );
  INV_X1 U628 ( .A(n705), .ZN(n626) );
  AND2_X1 U629 ( .A1(n576), .A2(n705), .ZN(n536) );
  AND2_X1 U630 ( .A1(n710), .A2(n536), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n361), .A2(n537), .ZN(n649) );
  INV_X1 U632 ( .A(n707), .ZN(n539) );
  OR2_X1 U633 ( .A1(n576), .A2(n539), .ZN(n704) );
  NOR2_X1 U634 ( .A1(n592), .A2(n591), .ZN(n540) );
  NAND2_X1 U635 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X2 U636 ( .A(n543), .B(n542), .ZN(n653) );
  INV_X1 U637 ( .A(n395), .ZN(n547) );
  XOR2_X1 U638 ( .A(n545), .B(n544), .Z(n579) );
  NAND2_X1 U639 ( .A1(n393), .A2(n546), .ZN(n715) );
  NOR2_X1 U640 ( .A1(n704), .A2(n590), .ZN(n548) );
  NAND2_X1 U641 ( .A1(n710), .A2(n548), .ZN(n549) );
  XNOR2_X1 U642 ( .A(n592), .B(KEYINPUT100), .ZN(n554) );
  INV_X1 U643 ( .A(KEYINPUT102), .ZN(n551) );
  AND2_X1 U644 ( .A1(n554), .A2(n553), .ZN(n679) );
  INV_X1 U645 ( .A(n576), .ZN(n708) );
  NAND2_X1 U646 ( .A1(n708), .A2(n705), .ZN(n555) );
  INV_X1 U647 ( .A(KEYINPUT82), .ZN(n556) );
  INV_X1 U648 ( .A(n653), .ZN(n557) );
  NOR2_X1 U649 ( .A1(n557), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U651 ( .A(KEYINPUT45), .ZN(n561) );
  OR2_X1 U652 ( .A1(n752), .A2(n563), .ZN(n564) );
  NOR2_X1 U653 ( .A1(G900), .A2(n564), .ZN(n565) );
  XOR2_X1 U654 ( .A(KEYINPUT105), .B(n565), .Z(n566) );
  NOR2_X1 U655 ( .A1(n567), .A2(n566), .ZN(n578) );
  NAND2_X1 U656 ( .A1(n579), .A2(n696), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n568), .B(KEYINPUT30), .ZN(n569) );
  NOR2_X1 U658 ( .A1(n578), .A2(n569), .ZN(n571) );
  INV_X1 U659 ( .A(n704), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n571), .A2(n570), .ZN(n596) );
  NOR2_X1 U661 ( .A1(n596), .A2(n590), .ZN(n572) );
  NAND2_X1 U662 ( .A1(n572), .A2(n697), .ZN(n573) );
  XNOR2_X1 U663 ( .A(n573), .B(KEYINPUT39), .ZN(n631) );
  NAND2_X1 U664 ( .A1(n631), .A2(n682), .ZN(n575) );
  XOR2_X1 U665 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n574) );
  XNOR2_X1 U666 ( .A(n575), .B(n574), .ZN(n761) );
  NAND2_X1 U667 ( .A1(n576), .A2(n707), .ZN(n577) );
  INV_X1 U668 ( .A(n590), .ZN(n580) );
  XNOR2_X1 U669 ( .A(n581), .B(KEYINPUT109), .ZN(n603) );
  INV_X1 U670 ( .A(n697), .ZN(n583) );
  NAND2_X1 U671 ( .A1(n698), .A2(n696), .ZN(n582) );
  NOR2_X1 U672 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n584), .B(KEYINPUT41), .ZN(n726) );
  NOR2_X1 U674 ( .A1(n603), .A2(n726), .ZN(n587) );
  XOR2_X1 U675 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n585) );
  XNOR2_X1 U676 ( .A(n585), .B(KEYINPUT111), .ZN(n586) );
  XNOR2_X1 U677 ( .A(n587), .B(n586), .ZN(n648) );
  NOR2_X1 U678 ( .A1(n761), .A2(n648), .ZN(n588) );
  XNOR2_X1 U679 ( .A(n588), .B(KEYINPUT46), .ZN(n622) );
  NAND2_X1 U680 ( .A1(KEYINPUT47), .A2(n695), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n591), .A2(n590), .ZN(n594) );
  INV_X1 U682 ( .A(n592), .ZN(n593) );
  NAND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n597), .A2(n398), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n600), .A2(n760), .ZN(n602) );
  XNOR2_X1 U686 ( .A(n602), .B(n601), .ZN(n607) );
  INV_X1 U687 ( .A(n603), .ZN(n605) );
  INV_X1 U688 ( .A(n360), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n617), .A2(KEYINPUT47), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n609) );
  AND2_X1 U692 ( .A1(n682), .A2(n610), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n625) );
  BUF_X1 U694 ( .A(n613), .Z(n614) );
  NOR2_X1 U695 ( .A1(n625), .A2(n614), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT36), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n616), .A2(n626), .ZN(n690) );
  NOR2_X1 U698 ( .A1(n695), .A2(KEYINPUT47), .ZN(n618) );
  INV_X1 U699 ( .A(n617), .ZN(n683) );
  NAND2_X1 U700 ( .A1(n618), .A2(n683), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n690), .A2(n619), .ZN(n620) );
  XNOR2_X1 U702 ( .A(KEYINPUT69), .B(KEYINPUT48), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n696), .A2(n627), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  XOR2_X1 U706 ( .A(KEYINPUT106), .B(n629), .Z(n630) );
  NOR2_X1 U707 ( .A1(n630), .A2(n398), .ZN(n650) );
  NAND2_X1 U708 ( .A1(n631), .A2(n679), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT113), .ZN(n759) );
  NOR2_X1 U710 ( .A1(n650), .A2(n759), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n751) );
  INV_X1 U712 ( .A(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n356), .A2(n636), .ZN(n637) );
  INV_X1 U714 ( .A(KEYINPUT76), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n665), .A2(G478), .ZN(n641) );
  INV_X1 U716 ( .A(G952), .ZN(n642) );
  AND2_X1 U717 ( .A1(n642), .A2(G953), .ZN(n670) );
  NAND2_X1 U718 ( .A1(n665), .A2(G469), .ZN(n646) );
  XOR2_X1 U719 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n643) );
  XNOR2_X1 U720 ( .A(n643), .B(KEYINPUT58), .ZN(n644) );
  XOR2_X1 U721 ( .A(G137), .B(KEYINPUT126), .Z(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(G39) );
  XNOR2_X1 U723 ( .A(n649), .B(G110), .ZN(G12) );
  XOR2_X1 U724 ( .A(G140), .B(n650), .Z(G42) );
  XOR2_X1 U725 ( .A(G101), .B(n651), .Z(G3) );
  INV_X1 U726 ( .A(n679), .ZN(n674) );
  XOR2_X1 U727 ( .A(G116), .B(n652), .Z(G18) );
  XNOR2_X1 U728 ( .A(n394), .B(G122), .ZN(G24) );
  NAND2_X1 U729 ( .A1(n665), .A2(G475), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n665), .A2(G210), .ZN(n661) );
  BUF_X1 U731 ( .A(n656), .Z(n657) );
  XOR2_X1 U732 ( .A(KEYINPUT87), .B(KEYINPUT54), .Z(n659) );
  XNOR2_X1 U733 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n665), .A2(G472), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(G119), .ZN(G21) );
  BUF_X1 U737 ( .A(n665), .Z(n666) );
  NAND2_X1 U738 ( .A1(n666), .A2(G217), .ZN(n669) );
  XOR2_X1 U739 ( .A(KEYINPUT124), .B(n667), .Z(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n671) );
  NOR2_X1 U741 ( .A1(n671), .A2(n670), .ZN(G66) );
  INV_X1 U742 ( .A(n682), .ZN(n686) );
  NOR2_X1 U743 ( .A1(n675), .A2(n686), .ZN(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT114), .B(n672), .Z(n673) );
  XNOR2_X1 U745 ( .A(G104), .B(n673), .ZN(G6) );
  XOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n677) );
  NOR2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U748 ( .A(n677), .B(n676), .Z(n678) );
  XNOR2_X1 U749 ( .A(G107), .B(n678), .ZN(G9) );
  XOR2_X1 U750 ( .A(n345), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U751 ( .A1(n683), .A2(n679), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(G30) );
  XOR2_X1 U753 ( .A(G146), .B(KEYINPUT115), .Z(n685) );
  NAND2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n685), .B(n684), .ZN(G48) );
  XOR2_X1 U756 ( .A(KEYINPUT116), .B(n687), .Z(n688) );
  XNOR2_X1 U757 ( .A(G113), .B(n688), .ZN(G15) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n689) );
  XNOR2_X1 U759 ( .A(n690), .B(n689), .ZN(G27) );
  NOR2_X1 U760 ( .A1(n356), .A2(KEYINPUT2), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n396), .A2(n692), .ZN(n732) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n700) );
  INV_X1 U765 ( .A(n698), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U768 ( .A1(n703), .A2(n727), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U770 ( .A(n706), .B(KEYINPUT50), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n709), .B(KEYINPUT49), .ZN(n711) );
  NAND2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U774 ( .A(KEYINPUT117), .B(n712), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n717), .ZN(n718) );
  NOR2_X1 U778 ( .A1(n718), .A2(n726), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U780 ( .A(n721), .B(KEYINPUT118), .ZN(n722) );
  XNOR2_X1 U781 ( .A(KEYINPUT52), .B(n722), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U783 ( .A(KEYINPUT119), .B(n725), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U786 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U788 ( .A(KEYINPUT53), .B(n733), .ZN(G75) );
  NOR2_X1 U789 ( .A1(n734), .A2(G953), .ZN(n739) );
  NAND2_X1 U790 ( .A1(G953), .A2(G224), .ZN(n735) );
  XOR2_X1 U791 ( .A(KEYINPUT61), .B(n735), .Z(n736) );
  NOR2_X1 U792 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n747) );
  XOR2_X1 U794 ( .A(n740), .B(KEYINPUT125), .Z(n741) );
  XNOR2_X1 U795 ( .A(n392), .B(n741), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n743), .B(G101), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(G69) );
  XNOR2_X1 U799 ( .A(KEYINPUT4), .B(n748), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n749), .B(n750), .ZN(n754) );
  XNOR2_X1 U801 ( .A(n751), .B(n754), .ZN(n753) );
  NAND2_X1 U802 ( .A1(n753), .A2(n752), .ZN(n758) );
  XNOR2_X1 U803 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U805 ( .A1(G953), .A2(n756), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U807 ( .A(G134), .B(n759), .Z(G36) );
  XNOR2_X1 U808 ( .A(G143), .B(n760), .ZN(G45) );
  XOR2_X1 U809 ( .A(G131), .B(n761), .Z(G33) );
endmodule

