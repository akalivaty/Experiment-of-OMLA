//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT71), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT23), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  AND4_X1   g008(.A1(KEYINPUT25), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(KEYINPUT24), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n213), .B(new_n214), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n210), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  AND3_X1   g021(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G183gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n212), .B1(KEYINPUT65), .B2(KEYINPUT28), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n231), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G190gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n230), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT26), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n209), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G169gat), .A2(G176gat), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(KEYINPUT26), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(new_n215), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n237), .A2(new_n241), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n203), .B1(new_n229), .B2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT25), .A4(new_n209), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n223), .A2(new_n225), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n218), .A2(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(KEYINPUT64), .B2(new_n218), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n215), .A2(new_n218), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n213), .A3(new_n214), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n248), .B1(new_n254), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n249), .B1(new_n261), .B2(new_n203), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  XNOR2_X1  g062(.A(G211gat), .B(G218gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266));
  INV_X1    g065(.A(G218gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT69), .A2(G218gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT22), .B1(new_n270), .B2(G211gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n263), .B(new_n265), .C1(new_n271), .C2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n265), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  INV_X1    g074(.A(G211gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n268), .B2(new_n269), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n264), .B(new_n272), .C1(new_n277), .C2(KEYINPUT22), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n279), .B2(new_n263), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT72), .B1(new_n261), .B2(new_n203), .ZN(new_n282));
  INV_X1    g081(.A(new_n203), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT29), .B1(new_n229), .B2(new_n248), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(KEYINPUT72), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT37), .B(new_n281), .C1(new_n287), .C2(new_n280), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT37), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n283), .B1(new_n259), .B2(new_n260), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT72), .B1(new_n290), .B2(new_n249), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n285), .B2(new_n283), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n280), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n281), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n288), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT38), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n291), .A2(new_n280), .A3(new_n293), .ZN(new_n305));
  INV_X1    g104(.A(new_n280), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n289), .B1(new_n286), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT38), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n296), .A2(new_n302), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT82), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n301), .B1(new_n294), .B2(new_n295), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n308), .A3(new_n312), .A4(new_n302), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n304), .A2(new_n310), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT2), .ZN(new_n319));
  OR2_X1    g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G155gat), .B(G162gat), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(KEYINPUT75), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n322), .B2(KEYINPUT75), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G141gat), .B(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(G155gat), .B2(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT75), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n323), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n322), .A2(KEYINPUT75), .A3(new_n323), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(KEYINPUT3), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n335));
  INV_X1    g134(.A(G127gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G134gat), .ZN(new_n337));
  INV_X1    g136(.A(G134gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(G127gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n335), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(G127gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n336), .A2(G134gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT66), .ZN(new_n343));
  INV_X1    g142(.A(G113gat), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT1), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G113gat), .A2(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n340), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n341), .A2(new_n342), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n350), .A2(new_n335), .A3(new_n347), .A4(new_n346), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n326), .A2(new_n334), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n326), .A2(new_n334), .A3(new_n352), .A4(KEYINPUT76), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n316), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n332), .A2(new_n333), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n349), .A2(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT4), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n332), .A2(new_n333), .B1(new_n349), .B2(new_n351), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT78), .A3(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(new_n358), .A3(new_n369), .ZN(new_n370));
  AOI221_X4 g169(.A(new_n316), .B1(new_n366), .B2(new_n362), .C1(new_n355), .C2(new_n356), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n332), .A2(new_n333), .A3(new_n349), .A4(new_n351), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT77), .B1(new_n373), .B2(new_n316), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n375), .B(new_n315), .C1(new_n365), .C2(new_n372), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT5), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n359), .A2(new_n361), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n316), .B1(new_n384), .B2(new_n367), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n375), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n373), .A2(KEYINPUT77), .A3(new_n316), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n358), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n355), .A2(new_n356), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n366), .A2(new_n362), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n315), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n360), .B1(new_n359), .B2(new_n361), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(KEYINPUT78), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT5), .B1(new_n394), .B2(new_n364), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n388), .A2(new_n391), .B1(new_n395), .B2(new_n357), .ZN(new_n396));
  INV_X1    g195(.A(new_n382), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT6), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n388), .A2(new_n391), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n402), .B2(new_n370), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n403), .B2(KEYINPUT6), .ZN(new_n404));
  NOR4_X1   g203(.A1(new_n396), .A2(KEYINPUT83), .A3(new_n399), .A4(new_n397), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n314), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n260), .B(new_n274), .C1(new_n279), .C2(new_n263), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n359), .B1(new_n408), .B2(new_n317), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n326), .A2(new_n260), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n280), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(G228gat), .B(G233gat), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n359), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n279), .A2(new_n414), .A3(new_n260), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n317), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n279), .B2(new_n260), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n280), .A2(new_n410), .B1(G228gat), .B2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n412), .B2(new_n420), .ZN(new_n425));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(G22gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n420), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n421), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n432), .B2(new_n423), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n315), .B1(new_n389), .B2(new_n369), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT39), .B1(new_n373), .B2(new_n316), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT39), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n382), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n437), .A2(new_n439), .A3(KEYINPUT40), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n383), .A3(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n281), .B(new_n302), .C1(new_n287), .C2(new_n280), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n311), .A3(KEYINPUT30), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n281), .B1(new_n287), .B2(new_n280), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n301), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n434), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT84), .B1(new_n407), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n403), .A2(new_n401), .A3(KEYINPUT6), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT6), .B1(new_n378), .B2(new_n382), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n454), .A2(new_n455), .B1(new_n398), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n310), .A2(new_n313), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n303), .A2(KEYINPUT38), .B1(new_n447), .B2(new_n301), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n429), .B1(new_n424), .B2(new_n425), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n432), .A2(new_n428), .A3(new_n423), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n437), .A2(new_n439), .A3(KEYINPUT40), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT40), .B1(new_n437), .B2(new_n439), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(new_n403), .ZN(new_n466));
  INV_X1    g265(.A(new_n450), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n399), .B1(new_n396), .B2(new_n397), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n378), .A2(new_n382), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n453), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n450), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT81), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT36), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n352), .B1(new_n259), .B2(KEYINPUT67), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n257), .A2(new_n206), .A3(new_n209), .A4(new_n208), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(new_n222), .B1(new_n210), .B2(new_n220), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n235), .A2(new_n231), .A3(new_n236), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n230), .B1(new_n238), .B2(new_n240), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n246), .B(new_n215), .C1(new_n243), .C2(new_n244), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT67), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n229), .A2(new_n489), .A3(new_n248), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n481), .B1(new_n491), .B2(new_n352), .ZN(new_n492));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n229), .A2(new_n489), .A3(new_n248), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n489), .B1(new_n229), .B2(new_n248), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n352), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n481), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n493), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n496), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT33), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  XOR2_X1   g305(.A(G15gat), .B(G43gat), .Z(new_n507));
  XNOR2_X1  g306(.A(G71gat), .B(G99gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n498), .B(new_n505), .C1(new_n506), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n361), .B1(new_n488), .B2(new_n490), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n504), .B1(new_n512), .B2(new_n481), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n497), .B1(new_n492), .B2(new_n493), .ZN(new_n516));
  NOR4_X1   g315(.A1(new_n512), .A2(new_n481), .A3(new_n504), .A4(new_n496), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n515), .B(new_n509), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n513), .A2(KEYINPUT32), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n511), .B2(new_n518), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n480), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n511), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n519), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT36), .A3(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n479), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n526), .A2(new_n462), .A3(new_n461), .A4(new_n521), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT35), .B1(new_n531), .B2(new_n477), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n533));
  INV_X1    g332(.A(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n450), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n457), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT85), .B(KEYINPUT35), .C1(new_n531), .C2(new_n477), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n471), .A2(new_n530), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT12), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  OR2_X1    g347(.A1(G43gat), .A2(G50gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G43gat), .A2(G50gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT87), .B(G50gat), .Z(new_n553));
  OAI211_X1 g352(.A(new_n548), .B(new_n550), .C1(new_n553), .C2(G43gat), .ZN(new_n554));
  OR3_X1    g353(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT88), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n552), .A2(new_n554), .A3(new_n560), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G29gat), .A2(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n556), .A2(KEYINPUT86), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n555), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n556), .A2(KEYINPUT86), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n551), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT16), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G1gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G1gat), .B2(new_n570), .ZN(new_n573));
  INV_X1    g372(.A(G8gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n547), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n559), .A2(new_n561), .B1(new_n551), .B2(new_n567), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n578), .A2(new_n575), .A3(KEYINPUT89), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n577), .A2(new_n579), .B1(new_n569), .B2(new_n576), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT13), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n576), .B1(new_n569), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n578), .A2(KEYINPUT17), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n547), .A3(new_n576), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT89), .B1(new_n578), .B2(new_n575), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT90), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n591), .A2(KEYINPUT18), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n587), .A2(new_n590), .A3(new_n581), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n586), .A2(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n593), .B1(new_n596), .B2(new_n581), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n546), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n575), .B1(new_n578), .B2(KEYINPUT17), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n562), .A2(KEYINPUT17), .A3(new_n568), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n577), .A2(new_n579), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n581), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n592), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(new_n545), .A3(new_n583), .A4(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n540), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G78gat), .ZN(new_n608));
  XOR2_X1   g407(.A(G57gat), .B(G64gat), .Z(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(KEYINPUT9), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(KEYINPUT91), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n617), .B(KEYINPUT92), .Z(new_n618));
  OAI21_X1  g417(.A(new_n611), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(G127gat), .B(G155gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT93), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G183gat), .B(G211gat), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n626), .A2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n575), .B1(new_n620), .B2(new_n619), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OR3_X1    g433(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n634), .B1(new_n629), .B2(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n619), .ZN(new_n640));
  NAND2_X1  g439(.A1(G85gat), .A2(G92gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT7), .ZN(new_n642));
  NAND2_X1  g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(G85gat), .ZN(new_n644));
  INV_X1    g443(.A(G92gat), .ZN(new_n645));
  AOI22_X1  g444(.A1(KEYINPUT8), .A2(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G99gat), .B(G106gat), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n642), .A3(new_n646), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(KEYINPUT98), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n653));
  INV_X1    g452(.A(new_n651), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n642), .B2(new_n646), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n619), .A2(KEYINPUT98), .A3(new_n651), .A4(new_n649), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT10), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT95), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n654), .B2(new_n655), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n649), .A2(KEYINPUT95), .A3(new_n651), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n640), .A2(new_n661), .A3(KEYINPUT10), .A4(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n639), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n657), .A2(new_n658), .ZN(new_n666));
  INV_X1    g465(.A(new_n639), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n665), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT99), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n665), .A2(new_n668), .A3(new_n674), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n665), .B2(new_n668), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT100), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n680), .B(new_n677), .C1(new_n673), .C2(new_n675), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G190gat), .B(G218gat), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT96), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n661), .A2(new_n662), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n578), .B2(KEYINPUT17), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n600), .ZN(new_n688));
  AND2_X1   g487(.A1(G232gat), .A2(G233gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(KEYINPUT41), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n578), .B2(new_n686), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n684), .B(new_n685), .C1(new_n688), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n569), .A2(new_n584), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n586), .A3(new_n686), .ZN(new_n694));
  INV_X1    g493(.A(new_n691), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(KEYINPUT96), .A3(new_n695), .A4(new_n683), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n692), .A2(KEYINPUT94), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT97), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n689), .A2(KEYINPUT41), .ZN(new_n699));
  XNOR2_X1  g498(.A(G134gat), .B(G162gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT97), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n692), .A2(new_n703), .A3(new_n696), .ZN(new_n704));
  INV_X1    g503(.A(new_n701), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n697), .A2(KEYINPUT97), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n638), .A2(new_n682), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n607), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n476), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT101), .B(G1gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1324gat));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n607), .A2(new_n467), .A3(new_n708), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G8gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(KEYINPUT103), .A3(new_n574), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT16), .B(G8gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n607), .A2(new_n720), .A3(new_n467), .A4(new_n708), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n716), .A2(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR4_X1   g522(.A1(new_n714), .A2(new_n720), .A3(KEYINPUT42), .A4(new_n718), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n715), .A2(new_n717), .B1(new_n723), .B2(new_n724), .ZN(G1325gat));
  AND3_X1   g524(.A1(new_n524), .A2(KEYINPUT104), .A3(new_n527), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT104), .B1(new_n524), .B2(new_n527), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G15gat), .B1(new_n709), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n522), .A2(new_n523), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n732), .A2(G15gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n709), .B2(new_n733), .ZN(G1326gat));
  NAND2_X1  g533(.A1(new_n473), .A2(new_n478), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n607), .A2(new_n736), .A3(new_n708), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT43), .B(G22gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1327gat));
  INV_X1    g541(.A(new_n682), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n638), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n606), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n532), .A2(new_n533), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n537), .A2(new_n534), .ZN(new_n747));
  AND3_X1   g546(.A1(new_n746), .A2(new_n539), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n529), .B1(new_n452), .B2(new_n470), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n707), .B(new_n745), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n476), .A2(G29gat), .ZN(new_n751));
  OR3_X1    g550(.A1(new_n750), .A2(KEYINPUT106), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n756));
  INV_X1    g555(.A(new_n707), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n540), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n707), .C1(new_n748), .C2(new_n749), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n745), .ZN(new_n761));
  OAI21_X1  g560(.A(G29gat), .B1(new_n761), .B2(new_n476), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n755), .A2(new_n762), .A3(new_n763), .ZN(G1328gat));
  OAI21_X1  g563(.A(G36gat), .B1(new_n761), .B2(new_n450), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n750), .A2(G36gat), .A3(new_n450), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT46), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1329gat));
  INV_X1    g567(.A(new_n528), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n760), .A2(new_n769), .A3(new_n745), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G43gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n732), .A2(G43gat), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n750), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n471), .A2(new_n530), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n538), .A2(new_n539), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n757), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(KEYINPUT107), .A3(new_n745), .A4(new_n773), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n758), .A2(new_n728), .A3(new_n745), .A4(new_n759), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G43gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n780), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n783), .A2(G43gat), .B1(new_n775), .B2(new_n779), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n788), .A2(KEYINPUT108), .A3(KEYINPUT47), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n781), .B1(new_n787), .B2(new_n789), .ZN(G1330gat));
  NOR4_X1   g589(.A1(new_n744), .A2(new_n553), .A3(new_n735), .A4(new_n757), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n607), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT48), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n758), .A2(new_n463), .A3(new_n745), .A4(new_n759), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n553), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(KEYINPUT109), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n797), .B(new_n793), .C1(new_n794), .C2(new_n553), .ZN(new_n798));
  INV_X1    g597(.A(new_n792), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n760), .A2(new_n736), .A3(new_n745), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n553), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n796), .A2(new_n798), .B1(KEYINPUT48), .B2(new_n801), .ZN(G1331gat));
  NAND2_X1  g601(.A1(new_n776), .A2(new_n777), .ZN(new_n803));
  NOR4_X1   g602(.A1(new_n743), .A2(new_n638), .A3(new_n605), .A4(new_n707), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n476), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g608(.A1(new_n805), .A2(new_n450), .ZN(new_n810));
  NOR2_X1   g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  AND2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n810), .B2(new_n811), .ZN(G1333gat));
  OR3_X1    g613(.A1(new_n805), .A2(KEYINPUT111), .A3(new_n732), .ZN(new_n815));
  INV_X1    g614(.A(G71gat), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT111), .B1(new_n805), .B2(new_n732), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n803), .A2(G71gat), .A3(new_n728), .A4(new_n804), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT110), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1334gat));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n736), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g626(.A1(new_n637), .A2(new_n605), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT112), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n682), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n760), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G85gat), .B1(new_n831), .B2(new_n476), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n778), .A2(KEYINPUT113), .A3(KEYINPUT51), .A4(new_n829), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n803), .A2(new_n707), .A3(new_n829), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(KEYINPUT51), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT113), .B1(new_n834), .B2(KEYINPUT51), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n682), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n807), .A2(new_n644), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n834), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n778), .A2(new_n829), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n450), .A2(G92gat), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n682), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n758), .A2(new_n467), .A3(new_n759), .A4(new_n830), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G92gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n848), .B2(G92gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n845), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n837), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1337gat));
  INV_X1    g654(.A(G99gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n831), .A2(new_n856), .A3(new_n729), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n731), .B(new_n682), .C1(new_n835), .C2(new_n836), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(G1338gat));
  NOR3_X1   g658(.A1(new_n743), .A2(G106gat), .A3(new_n434), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n835), .B2(new_n836), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n862));
  NAND4_X1  g661(.A1(new_n758), .A2(new_n463), .A3(new_n759), .A4(new_n830), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(G106gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT51), .B1(new_n843), .B2(KEYINPUT114), .ZN(new_n866));
  AOI211_X1 g665(.A(new_n841), .B(new_n840), .C1(new_n778), .C2(new_n829), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n758), .A2(new_n736), .A3(new_n759), .A4(new_n830), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n868), .A2(new_n860), .B1(G106gat), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n870), .B2(new_n871), .ZN(G1339gat));
  NOR2_X1   g671(.A1(new_n596), .A2(new_n581), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n580), .A2(new_n582), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n544), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n604), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n679), .B2(new_n681), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n667), .B(new_n663), .C1(new_n666), .C2(KEYINPUT10), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n878), .A2(KEYINPUT54), .A3(new_n665), .ZN(new_n879));
  INV_X1    g678(.A(new_n671), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n639), .C1(new_n659), .C2(new_n664), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n879), .A2(KEYINPUT55), .A3(new_n880), .A4(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n676), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n605), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n707), .B1(new_n877), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n887), .A2(new_n676), .A3(new_n883), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n707), .A2(new_n890), .A3(new_n876), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n638), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n743), .A2(new_n606), .A3(new_n637), .A4(new_n757), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n476), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n894), .A2(new_n450), .A3(new_n534), .ZN(new_n895));
  AOI21_X1  g694(.A(G113gat), .B1(new_n895), .B2(new_n605), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n638), .A2(new_n682), .A3(new_n707), .A4(new_n605), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n877), .A2(new_n888), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n757), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n707), .A2(new_n890), .A3(new_n876), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n901), .B2(new_n638), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n467), .A2(new_n476), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n902), .A2(new_n736), .A3(new_n732), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n606), .A2(new_n344), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(G1340gat));
  AOI21_X1  g706(.A(G120gat), .B1(new_n895), .B2(new_n682), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n743), .A2(new_n345), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n905), .B2(new_n909), .ZN(G1341gat));
  AND2_X1   g709(.A1(new_n895), .A2(new_n637), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(G127gat), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n638), .A2(new_n336), .ZN(new_n915));
  AOI22_X1  g714(.A1(new_n913), .A2(new_n914), .B1(new_n905), .B2(new_n915), .ZN(G1342gat));
  NAND3_X1  g715(.A1(new_n895), .A2(new_n338), .A3(new_n707), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(KEYINPUT56), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n338), .B1(new_n905), .B2(new_n707), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(KEYINPUT56), .B2(new_n917), .ZN(G1343gat));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n769), .A2(new_n904), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n735), .B1(new_n892), .B2(new_n893), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT57), .B(new_n434), .C1(new_n892), .C2(new_n893), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(G141gat), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n606), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n463), .B1(new_n726), .B2(new_n727), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n467), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n894), .A2(new_n933), .A3(new_n605), .A4(new_n934), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n928), .A2(new_n930), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n922), .B1(new_n936), .B2(KEYINPUT58), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT57), .B1(new_n902), .B2(new_n735), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n892), .A2(new_n893), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n925), .A3(new_n463), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n938), .A2(new_n940), .A3(new_n923), .A4(new_n930), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n935), .A2(new_n929), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n943), .A2(KEYINPUT118), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT119), .B1(new_n943), .B2(new_n944), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n947), .B(KEYINPUT58), .C1(new_n941), .C2(new_n942), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n937), .A2(new_n945), .B1(new_n946), .B2(new_n948), .ZN(G1344gat));
  NOR2_X1   g748(.A1(new_n743), .A2(G148gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n894), .A2(new_n933), .A3(new_n934), .A4(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n735), .A2(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n707), .A2(new_n890), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT120), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n876), .B1(new_n954), .B2(KEYINPUT120), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n899), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n638), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n953), .B1(new_n958), .B2(new_n897), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT57), .B1(new_n902), .B2(new_n434), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n959), .A2(new_n682), .A3(new_n923), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n952), .B1(new_n961), .B2(G148gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n952), .A2(G148gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n928), .B2(new_n682), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n951), .B1(new_n962), .B2(new_n964), .ZN(G1345gat));
  INV_X1    g764(.A(new_n928), .ZN(new_n966));
  OAI21_X1  g765(.A(G155gat), .B1(new_n966), .B2(new_n638), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n638), .A2(G155gat), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n894), .A2(new_n933), .A3(new_n934), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n967), .A2(new_n969), .ZN(G1346gat));
  NOR2_X1   g769(.A1(new_n757), .A2(G162gat), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n894), .A2(new_n933), .A3(new_n934), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT121), .B1(new_n966), .B2(new_n757), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G162gat), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n966), .A2(KEYINPUT121), .A3(new_n757), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1347gat));
  NOR2_X1   g775(.A1(new_n902), .A2(new_n736), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n467), .A2(new_n476), .ZN(new_n978));
  XOR2_X1   g777(.A(new_n978), .B(KEYINPUT123), .Z(new_n979));
  NOR2_X1   g778(.A1(new_n979), .A2(new_n732), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n981), .A2(new_n204), .A3(new_n606), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n902), .A2(new_n983), .A3(new_n807), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT122), .B1(new_n939), .B2(new_n476), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n531), .A2(new_n450), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n986), .A2(new_n605), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n982), .B1(new_n988), .B2(new_n204), .ZN(G1348gat));
  OAI21_X1  g788(.A(G176gat), .B1(new_n981), .B2(new_n743), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n987), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n682), .A2(new_n205), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G1349gat));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n637), .A3(new_n980), .ZN(new_n994));
  AOI22_X1  g793(.A1(new_n994), .A2(G183gat), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n995));
  OR2_X1    g794(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n638), .A2(new_n235), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n987), .B(new_n997), .C1(new_n984), .C2(new_n985), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n996), .B1(new_n995), .B2(new_n998), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n999), .A2(new_n1000), .ZN(G1350gat));
  NAND2_X1  g800(.A1(new_n707), .A2(new_n212), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n977), .A2(new_n707), .A3(new_n980), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT61), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1003), .A2(new_n1004), .A3(G190gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n1004), .B1(new_n1003), .B2(G190gat), .ZN(new_n1006));
  OAI22_X1  g805(.A1(new_n991), .A2(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1351gat));
  NOR2_X1   g806(.A1(new_n979), .A2(new_n728), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n959), .A2(new_n960), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(G197gat), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n1009), .A2(new_n1010), .A3(new_n606), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n931), .A2(new_n450), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n986), .A2(new_n605), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1011), .B1(new_n1010), .B2(new_n1013), .ZN(G1352gat));
  XOR2_X1   g813(.A(KEYINPUT125), .B(G204gat), .Z(new_n1015));
  NOR2_X1   g814(.A1(new_n743), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g815(.A(new_n1012), .B(new_n1016), .C1(new_n984), .C2(new_n985), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n1015), .B1(new_n1009), .B2(new_n743), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(G1353gat));
  NAND4_X1  g820(.A1(new_n986), .A2(new_n276), .A3(new_n637), .A4(new_n1012), .ZN(new_n1022));
  NAND4_X1  g821(.A1(new_n959), .A2(new_n637), .A3(new_n960), .A4(new_n1008), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1023), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1023), .B2(G211gat), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(G1354gat));
  NAND2_X1  g825(.A1(new_n707), .A2(new_n270), .ZN(new_n1027));
  AND3_X1   g826(.A1(new_n959), .A2(new_n960), .A3(new_n1008), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT126), .ZN(new_n1029));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1009), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n986), .A2(new_n707), .A3(new_n1012), .ZN(new_n1032));
  AOI22_X1  g831(.A1(new_n1029), .A2(new_n1031), .B1(new_n267), .B2(new_n1032), .ZN(G1355gat));
endmodule


