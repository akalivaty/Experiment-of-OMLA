//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT91), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G15gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G15gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(G15gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(G22gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AND4_X1   g013(.A1(new_n203), .A2(new_n209), .A3(new_n210), .A4(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  AOI21_X1  g015(.A(G8gat), .B1(new_n216), .B2(new_n213), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n203), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(G1gat), .B1(new_n211), .B2(new_n212), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n216), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n223));
  OAI21_X1  g022(.A(G8gat), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT90), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT89), .B1(new_n216), .B2(G1gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n221), .B(new_n204), .C1(new_n206), .C2(new_n208), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n214), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n229), .A3(G8gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n219), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G36gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT14), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G29gat), .B2(G36gat), .ZN(new_n237));
  INV_X1    g036(.A(G29gat), .ZN(new_n238));
  INV_X1    g037(.A(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT14), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n235), .A2(KEYINPUT15), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT15), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n232), .B2(new_n233), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n237), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NOR4_X1   g046(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n242), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT17), .ZN(new_n251));
  INV_X1    g050(.A(new_n246), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n243), .A2(new_n244), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(KEYINPUT15), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n248), .B1(new_n254), .B2(new_n245), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT17), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n231), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n231), .A2(new_n259), .A3(new_n255), .ZN(new_n260));
  INV_X1    g059(.A(new_n218), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n217), .A2(new_n203), .A3(new_n209), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n228), .A2(new_n229), .A3(G8gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n229), .B1(new_n228), .B2(G8gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT92), .B1(new_n266), .B2(new_n250), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n202), .B(new_n258), .C1(new_n260), .C2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT18), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n259), .B1(new_n231), .B2(new_n255), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(KEYINPUT92), .A3(new_n250), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n258), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n231), .A2(new_n255), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n275), .B1(new_n260), .B2(new_n267), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(new_n202), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT87), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G141gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G169gat), .B(G197gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT12), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n280), .A2(KEYINPUT87), .A3(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G190gat), .B(G218gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G134gat), .B(G162gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT41), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(G99gat), .A2(G106gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT98), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G99gat), .ZN(new_n302));
  INV_X1    g101(.A(G106gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305));
  NAND2_X1  g104(.A1(G99gat), .A2(G106gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G92gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT97), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT97), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G92gat), .ZN(new_n312));
  INV_X1    g111(.A(G85gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G85gat), .A2(G92gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT7), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G85gat), .A3(G92gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n306), .A2(KEYINPUT8), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT8), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(G99gat), .B2(G106gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT97), .B(G92gat), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(new_n313), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n301), .A2(new_n307), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n319), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n322), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT99), .A4(new_n319), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n330), .A2(new_n331), .B1(new_n247), .B2(new_n249), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n296), .A2(KEYINPUT41), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT100), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT100), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n332), .B2(new_n334), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n330), .A2(new_n331), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n250), .A2(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n255), .A2(new_n256), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n298), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n297), .B(new_n343), .C1(new_n336), .C2(new_n338), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n295), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n338), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n332), .A2(new_n337), .A3(new_n334), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n297), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n339), .A2(new_n344), .A3(new_n298), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n294), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n355));
  NAND2_X1  g154(.A1(G231gat), .A2(G233gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G183gat), .B(G211gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G64gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G71gat), .ZN(new_n363));
  INV_X1    g162(.A(G78gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G71gat), .A2(G78gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT9), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n366), .B(new_n365), .C1(new_n361), .C2(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT94), .ZN(new_n375));
  XNOR2_X1  g174(.A(G127gat), .B(G155gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n376), .B(KEYINPUT95), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n374), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n372), .A2(new_n373), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT96), .B1(new_n266), .B2(new_n384), .ZN(new_n385));
  OR3_X1    g184(.A1(new_n266), .A2(KEYINPUT96), .A3(new_n384), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n360), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n385), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n378), .A3(new_n382), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n359), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G120gat), .B(G148gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G176gat), .B(G204gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G230gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT10), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n340), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT102), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT102), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n340), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n371), .B(new_n370), .C1(new_n308), .C2(new_n321), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n327), .B1(new_n319), .B2(new_n326), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT101), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n370), .A2(new_n371), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT101), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n328), .A4(new_n322), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT10), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n330), .A2(new_n372), .A3(new_n331), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n400), .B1(new_n407), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n399), .B1(new_n414), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n398), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n405), .B1(new_n340), .B2(new_n402), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT102), .B(new_n401), .C1(new_n330), .C2(new_n331), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n399), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n419), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n397), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n354), .A2(new_n394), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G183gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT27), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G183gat), .ZN(new_n434));
  INV_X1    g233(.A(G190gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT28), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT27), .B(G183gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  NOR2_X1   g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443));
  NAND2_X1  g242(.A1(G169gat), .A2(G176gat), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n441), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n437), .A2(new_n440), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT66), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n445), .A2(new_n446), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n440), .A4(new_n437), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT69), .ZN(new_n453));
  INV_X1    g252(.A(G134gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G127gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT67), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT68), .B1(new_n454), .B2(G127gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n454), .A3(G127gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460));
  INV_X1    g259(.A(G127gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(G134gat), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n456), .A2(new_n457), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464));
  INV_X1    g263(.A(G113gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(G120gat), .ZN(new_n466));
  INV_X1    g265(.A(G120gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(G113gat), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G127gat), .B(G134gat), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(new_n464), .C1(new_n466), .C2(new_n468), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT64), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n441), .B2(KEYINPUT23), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n441), .A2(KEYINPUT23), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n475), .A2(new_n476), .A3(new_n444), .ZN(new_n477));
  NOR2_X1   g276(.A1(G183gat), .A2(G190gat), .ZN(new_n478));
  AND2_X1   g277(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(G190gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G183gat), .A2(G190gat), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT24), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT65), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n485), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT23), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n477), .A2(new_n487), .A3(KEYINPUT25), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n444), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(KEYINPUT23), .B2(new_n441), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n431), .A2(new_n435), .ZN(new_n493));
  NAND3_X1  g292(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n483), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n492), .A2(new_n495), .A3(new_n489), .A4(new_n475), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT25), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n452), .A2(new_n453), .A3(new_n473), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n473), .A3(new_n448), .A4(new_n451), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n448), .A3(new_n451), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n470), .A2(new_n472), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT70), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n508), .A2(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n507), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT33), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G15gat), .B(G43gat), .Z(new_n517));
  XNOR2_X1  g316(.A(G71gat), .B(G99gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT33), .B1(new_n506), .B2(new_n507), .ZN(new_n521));
  INV_X1    g320(.A(new_n519), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n521), .A2(KEYINPUT34), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n511), .B(new_n512), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n513), .A3(new_n519), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT34), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n508), .A2(new_n510), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n508), .A2(new_n510), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n524), .A2(KEYINPUT36), .A3(new_n529), .ZN(new_n533));
  XOR2_X1   g332(.A(G78gat), .B(G106gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT76), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G50gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G155gat), .A2(G162gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT2), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(G141gat), .A2(G148gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(G141gat), .A2(G148gat), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(KEYINPUT72), .A3(KEYINPUT2), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OR3_X1    g346(.A1(KEYINPUT71), .A2(G155gat), .A3(G162gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT71), .B1(G155gat), .B2(G162gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n548), .A2(new_n549), .B1(G155gat), .B2(G162gat), .ZN(new_n550));
  INV_X1    g349(.A(G155gat), .ZN(new_n551));
  INV_X1    g350(.A(G162gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n539), .B1(new_n553), .B2(KEYINPUT2), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n547), .A2(new_n550), .B1(new_n545), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT3), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT29), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G211gat), .A2(G218gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(G211gat), .A2(G218gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G197gat), .A2(G204gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(G197gat), .A2(G204gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G211gat), .B(G218gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G197gat), .B(G204gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n564), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT78), .B1(new_n557), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n572));
  INV_X1    g371(.A(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n550), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n545), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n574), .A2(new_n556), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(KEYINPUT29), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G228gat), .A2(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT3), .B1(new_n570), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT77), .B1(new_n581), .B2(new_n555), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n574), .A2(new_n575), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT77), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT29), .B1(new_n565), .B2(new_n569), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n583), .B(new_n584), .C1(KEYINPUT3), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n579), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n578), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n557), .A2(new_n570), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n581), .A2(new_n555), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n579), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n207), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n578), .A2(KEYINPUT79), .A3(new_n587), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT79), .B1(new_n578), .B2(new_n587), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n207), .B(new_n595), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n538), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(G22gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n599), .A3(new_n537), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT4), .B1(new_n583), .B2(new_n504), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT4), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n555), .A2(new_n609), .A3(new_n470), .A4(new_n472), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n473), .A2(new_n555), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(KEYINPUT73), .A3(KEYINPUT4), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n555), .A2(new_n556), .B1(new_n470), .B2(new_n472), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n583), .A2(KEYINPUT3), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT5), .ZN(new_n618));
  NAND2_X1  g417(.A1(G225gat), .A2(G233gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n606), .B1(new_n614), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  AOI211_X1 g421(.A(KEYINPUT5), .B(new_n622), .C1(new_n615), .C2(new_n616), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(KEYINPUT74), .A3(new_n613), .A4(new_n611), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n504), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n612), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n618), .B1(new_n627), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n610), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n619), .A3(new_n617), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G1gat), .B(G29gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT0), .ZN(new_n634));
  XNOR2_X1  g433(.A(G57gat), .B(G85gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n621), .A2(new_n624), .B1(new_n630), .B2(new_n628), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n636), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n625), .A2(new_n636), .A3(new_n631), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n639), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G8gat), .B(G36gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G64gat), .B(G92gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G226gat), .A2(G233gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(KEYINPUT29), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n448), .A2(new_n451), .ZN(new_n652));
  AND4_X1   g451(.A1(KEYINPUT25), .A2(new_n492), .A3(new_n489), .A4(new_n475), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n653), .A2(new_n487), .B1(new_n496), .B2(new_n497), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n440), .A2(new_n437), .A3(new_n445), .A4(new_n446), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n498), .B2(new_n490), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n650), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n570), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n499), .A2(new_n448), .A3(new_n451), .A4(new_n650), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n573), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n648), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n503), .A2(new_n651), .B1(new_n657), .B2(new_n650), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n573), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n667), .A3(new_n647), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(KEYINPUT30), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n660), .A2(new_n663), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT30), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n671), .A3(new_n647), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n644), .A2(new_n673), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n532), .A2(new_n533), .B1(new_n605), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n676));
  AOI211_X1 g475(.A(KEYINPUT38), .B(new_n647), .C1(new_n670), .C2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT81), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n678), .B1(new_n666), .B2(new_n573), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n659), .A2(KEYINPUT81), .A3(new_n570), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n573), .A3(new_n662), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT82), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT82), .A4(new_n573), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n679), .A2(new_n680), .A3(new_n683), .A4(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT83), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT37), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n685), .B2(KEYINPUT37), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n677), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT37), .B1(new_n660), .B2(new_n663), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n665), .A2(new_n667), .ZN(new_n691));
  INV_X1    g490(.A(new_n676), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n690), .B(new_n648), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  AOI22_X1  g492(.A1(new_n693), .A2(KEYINPUT38), .B1(new_n647), .B2(new_n670), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n632), .A2(new_n637), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n641), .A2(new_n636), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n640), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n689), .A2(new_n694), .A3(new_n639), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n641), .A2(new_n636), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n673), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n611), .A2(new_n613), .A3(new_n617), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n622), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT39), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(new_n636), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(KEYINPUT39), .C1(new_n622), .C2(new_n627), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT80), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .A4(KEYINPUT40), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(new_n705), .A3(new_n636), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT80), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n700), .A2(new_n707), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n605), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT35), .ZN(new_n715));
  INV_X1    g514(.A(new_n530), .ZN(new_n716));
  INV_X1    g515(.A(new_n673), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n697), .B2(new_n639), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n675), .A2(new_n714), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n716), .A2(KEYINPUT85), .A3(new_n713), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n524), .A2(new_n601), .A3(new_n529), .A4(new_n604), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT85), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n674), .A2(new_n715), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI211_X1 g526(.A(new_n291), .B(new_n430), .C1(new_n720), .C2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n644), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT103), .B(G1gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1324gat));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(new_n717), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G8gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G8gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n728), .A2(new_n717), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n733), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n733), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n739), .A2(KEYINPUT105), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT105), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1325gat));
  AND3_X1   g542(.A1(new_n524), .A2(KEYINPUT36), .A3(new_n529), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT36), .B1(new_n524), .B2(new_n529), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n205), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n530), .A2(G15gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n728), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT106), .Z(G1326gat));
  NAND2_X1  g549(.A1(new_n728), .A2(new_n605), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT107), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT43), .B(G22gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1327gat));
  AOI21_X1  g553(.A(new_n354), .B1(new_n720), .B2(new_n727), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n291), .A2(new_n394), .A3(new_n428), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT108), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n234), .B1(new_n761), .B2(new_n644), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n755), .A2(new_n759), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n729), .A3(new_n232), .A4(new_n233), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(new_n765), .ZN(G1328gat));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n239), .A3(new_n717), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT46), .Z(new_n768));
  OAI21_X1  g567(.A(G36gat), .B1(new_n761), .B2(new_n673), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1329gat));
  NAND2_X1  g569(.A1(new_n763), .A2(new_n716), .ZN(new_n771));
  INV_X1    g570(.A(G43gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n746), .A2(G43gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n761), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n777), .B(new_n773), .C1(new_n761), .C2(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1330gat));
  NAND4_X1  g578(.A1(new_n756), .A2(new_n605), .A3(new_n757), .A4(new_n760), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n713), .A2(G50gat), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n780), .A2(G50gat), .B1(new_n763), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g582(.A1(new_n720), .A2(new_n727), .ZN(new_n784));
  AND4_X1   g583(.A1(new_n784), .A2(new_n291), .A3(new_n394), .A4(new_n354), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n785), .A2(new_n428), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n644), .B(KEYINPUT109), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g588(.A1(new_n429), .A2(new_n673), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT49), .B(G64gat), .Z(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(G1333gat));
  NAND3_X1  g593(.A1(new_n786), .A2(G71gat), .A3(new_n746), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n785), .A2(new_n428), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n530), .B(KEYINPUT110), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n363), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1334gat));
  NOR2_X1   g600(.A1(new_n796), .A2(new_n713), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n364), .ZN(G1335gat));
  AND3_X1   g602(.A1(new_n280), .A2(KEYINPUT87), .A3(new_n287), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n287), .B1(new_n280), .B2(KEYINPUT87), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n394), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n428), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n758), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810), .B2(new_n644), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n755), .B2(new_n807), .ZN(new_n812));
  INV_X1    g611(.A(new_n354), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n715), .B1(new_n722), .B2(new_n674), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n698), .A2(new_n712), .A3(new_n713), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n674), .A2(new_n605), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n744), .B2(new_n745), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n726), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n721), .B2(new_n724), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n813), .B(new_n807), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n812), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n729), .A2(new_n313), .A3(new_n428), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n811), .B1(new_n824), .B2(new_n825), .ZN(G1336gat));
  NAND4_X1  g625(.A1(new_n756), .A2(new_n717), .A3(new_n757), .A4(new_n809), .ZN(new_n827));
  INV_X1    g626(.A(new_n325), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n790), .A2(new_n309), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n812), .B2(new_n823), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT112), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n822), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n784), .A2(KEYINPUT51), .A3(new_n813), .A4(new_n807), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n830), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n834), .B(KEYINPUT52), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n833), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n839), .B2(new_n840), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT113), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(new_n829), .A3(new_n832), .A4(new_n841), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(G1337gat));
  INV_X1    g646(.A(new_n746), .ZN(new_n848));
  OAI21_X1  g647(.A(G99gat), .B1(new_n810), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n716), .A2(new_n302), .A3(new_n428), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n824), .B2(new_n850), .ZN(G1338gat));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n756), .A2(new_n605), .A3(new_n757), .A4(new_n809), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G106gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n605), .A2(new_n303), .A3(new_n428), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n824), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI221_X1 g658(.A(new_n854), .B1(new_n855), .B2(new_n852), .C1(new_n824), .C2(new_n857), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1339gat));
  OR2_X1    g660(.A1(new_n806), .A2(new_n430), .ZN(new_n862));
  INV_X1    g661(.A(new_n394), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n397), .B1(new_n418), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n407), .A2(new_n400), .A3(new_n417), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n425), .A2(KEYINPUT54), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n867), .A3(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n427), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n270), .A2(new_n279), .A3(new_n274), .A4(new_n287), .ZN(new_n870));
  INV_X1    g669(.A(new_n278), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n273), .A2(new_n275), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n202), .B1(new_n273), .B2(new_n258), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n286), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT55), .B1(new_n865), .B2(new_n867), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n869), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n863), .B1(new_n877), .B2(new_n354), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n428), .A2(new_n870), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n354), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n869), .A2(new_n876), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n806), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n862), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n787), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n725), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n673), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n465), .B1(new_n886), .B2(new_n291), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n806), .A2(new_n430), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n870), .A2(new_n874), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n865), .A2(new_n867), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT55), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n889), .A2(new_n427), .A3(new_n892), .A4(new_n868), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n394), .B1(new_n893), .B2(new_n813), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n879), .A2(new_n354), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n427), .A3(new_n868), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n291), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n888), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(new_n605), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n729), .A2(new_n673), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n716), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT115), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n806), .A2(G113gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n887), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT116), .ZN(G1340gat));
  NOR3_X1   g705(.A1(new_n903), .A2(new_n467), .A3(new_n429), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n885), .A2(new_n673), .A3(new_n428), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n467), .B2(new_n908), .ZN(G1341gat));
  OAI21_X1  g708(.A(G127gat), .B1(new_n903), .B2(new_n863), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n394), .A2(new_n461), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n886), .B2(new_n911), .ZN(G1342gat));
  NOR2_X1   g711(.A1(new_n354), .A2(new_n717), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n885), .A2(new_n454), .A3(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT56), .Z(new_n915));
  OAI21_X1  g714(.A(G134gat), .B1(new_n903), .B2(new_n354), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1343gat));
  NOR2_X1   g716(.A1(new_n746), .A2(new_n713), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n884), .A2(new_n673), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(G141gat), .A3(new_n291), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT58), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n848), .A2(new_n901), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n883), .A2(KEYINPUT57), .A3(new_n605), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n883), .B2(new_n605), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n927), .A2(new_n291), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n928), .A2(KEYINPUT118), .ZN(new_n929));
  OAI21_X1  g728(.A(G141gat), .B1(new_n928), .B2(KEYINPUT118), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n927), .A2(KEYINPUT117), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n923), .C1(new_n925), .C2(new_n926), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n806), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n920), .B1(new_n936), .B2(G141gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n931), .B1(new_n932), .B2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(G148gat), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n933), .A2(new_n935), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n939), .C1(new_n940), .C2(new_n428), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n898), .B2(new_n713), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n924), .A3(KEYINPUT119), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT119), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n946), .B(new_n943), .C1(new_n898), .C2(new_n713), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n923), .A2(new_n428), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g749(.A1(new_n950), .A2(KEYINPUT120), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n939), .B1(new_n950), .B2(KEYINPUT120), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n942), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n428), .A2(new_n939), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n941), .A2(new_n953), .B1(new_n919), .B2(new_n954), .ZN(G1345gat));
  AND2_X1   g754(.A1(new_n940), .A2(new_n394), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n394), .A2(new_n551), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n956), .A2(new_n551), .B1(new_n919), .B2(new_n957), .ZN(G1346gat));
  NAND4_X1  g757(.A1(new_n884), .A2(new_n552), .A3(new_n913), .A4(new_n918), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n940), .A2(new_n813), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n552), .ZN(G1347gat));
  OR2_X1    g760(.A1(new_n787), .A2(new_n673), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n962), .A2(KEYINPUT121), .A3(new_n797), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT121), .B1(new_n962), .B2(new_n797), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n899), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(G169gat), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(new_n291), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n898), .A2(new_n729), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(new_n725), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n969), .A2(new_n717), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n806), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n967), .B1(new_n971), .B2(new_n966), .ZN(G1348gat));
  OAI21_X1  g771(.A(G176gat), .B1(new_n965), .B2(new_n429), .ZN(new_n973));
  INV_X1    g772(.A(G176gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n969), .A2(new_n974), .A3(new_n790), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1349gat));
  AND2_X1   g775(.A1(new_n394), .A2(new_n438), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n963), .A2(new_n394), .A3(new_n899), .A4(new_n964), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G183gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n981), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT122), .B1(new_n981), .B2(KEYINPUT60), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n981), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n970), .A2(new_n977), .B1(G183gat), .B2(new_n979), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT60), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI22_X1  g787(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n988), .ZN(G1350gat));
  OAI21_X1  g788(.A(G190gat), .B1(new_n965), .B2(new_n354), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT61), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n435), .A3(new_n813), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1351gat));
  AND3_X1   g792(.A1(new_n968), .A2(new_n717), .A3(new_n918), .ZN(new_n994));
  INV_X1    g793(.A(G197gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n994), .A2(new_n995), .A3(new_n806), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n962), .A2(new_n746), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n998), .B1(new_n948), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n945), .A2(KEYINPUT124), .A3(new_n947), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1000), .A2(new_n806), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(KEYINPUT125), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G197gat), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1002), .A2(KEYINPUT125), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(G1352gat));
  NAND2_X1  g805(.A1(new_n948), .A2(new_n999), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n1007), .A2(new_n428), .A3(new_n1001), .A4(new_n997), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G204gat), .ZN(new_n1009));
  INV_X1    g808(.A(G204gat), .ZN(new_n1010));
  NAND4_X1  g809(.A1(new_n968), .A2(new_n1010), .A3(new_n790), .A4(new_n918), .ZN(new_n1011));
  XOR2_X1   g810(.A(new_n1011), .B(KEYINPUT62), .Z(new_n1012));
  NAND2_X1  g811(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT126), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1009), .A2(KEYINPUT126), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(G1353gat));
  INV_X1    g816(.A(G211gat), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n994), .A2(new_n1018), .A3(new_n394), .ZN(new_n1019));
  NAND2_X1  g818(.A1(new_n997), .A2(new_n394), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n948), .A2(new_n1020), .ZN(new_n1021));
  OR2_X1    g820(.A1(new_n1021), .A2(KEYINPUT127), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1018), .B1(new_n1021), .B2(KEYINPUT127), .ZN(new_n1023));
  AND3_X1   g822(.A1(new_n1022), .A2(KEYINPUT63), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g823(.A(KEYINPUT63), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1019), .B1(new_n1024), .B2(new_n1025), .ZN(G1354gat));
  AOI21_X1  g825(.A(G218gat), .B1(new_n994), .B2(new_n813), .ZN(new_n1027));
  AND2_X1   g826(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n813), .A2(G218gat), .ZN(new_n1029));
  AOI21_X1  g828(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(G1355gat));
endmodule


