

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U562 ( .A(n704), .B(KEYINPUT100), .ZN(n708) );
  XNOR2_X1 U563 ( .A(KEYINPUT97), .B(n731), .ZN(n783) );
  AND2_X1 U564 ( .A1(n825), .A2(n839), .ZN(n530) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n531) );
  XNOR2_X1 U566 ( .A(n571), .B(KEYINPUT13), .ZN(n532) );
  NOR2_X1 U567 ( .A1(n826), .A2(n530), .ZN(n533) );
  OR2_X1 U568 ( .A1(n781), .A2(n780), .ZN(n534) );
  NOR2_X1 U569 ( .A1(n1007), .A2(n703), .ZN(n709) );
  NOR2_X1 U570 ( .A1(n998), .A2(n709), .ZN(n710) );
  INV_X1 U571 ( .A(KEYINPUT29), .ZN(n723) );
  XNOR2_X1 U572 ( .A(n724), .B(n723), .ZN(n729) );
  AND2_X1 U573 ( .A1(n732), .A2(n783), .ZN(n757) );
  OR2_X1 U574 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U575 ( .A1(n541), .A2(n643), .ZN(n653) );
  NOR2_X1 U576 ( .A1(G651), .A2(n643), .ZN(n650) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n548) );
  XOR2_X1 U578 ( .A(KEYINPUT76), .B(n577), .Z(n1007) );
  INV_X1 U579 ( .A(G651), .ZN(n541) );
  XNOR2_X1 U580 ( .A(KEYINPUT68), .B(n531), .ZN(n643) );
  NAND2_X1 U581 ( .A1(n653), .A2(G77), .ZN(n535) );
  XOR2_X1 U582 ( .A(KEYINPUT71), .B(n535), .Z(n537) );
  NOR2_X1 U583 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U584 ( .A1(n649), .A2(G90), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U586 ( .A(n538), .B(KEYINPUT9), .ZN(n540) );
  NAND2_X1 U587 ( .A1(G52), .A2(n650), .ZN(n539) );
  NAND2_X1 U588 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U589 ( .A1(G543), .A2(n541), .ZN(n543) );
  XNOR2_X1 U590 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n542) );
  XNOR2_X1 U591 ( .A(n543), .B(n542), .ZN(n657) );
  NAND2_X1 U592 ( .A1(n657), .A2(G64), .ZN(n544) );
  XOR2_X1 U593 ( .A(KEYINPUT70), .B(n544), .Z(n545) );
  NOR2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U595 ( .A(KEYINPUT72), .B(n547), .ZN(G171) );
  INV_X1 U596 ( .A(G171), .ZN(G301) );
  XOR2_X2 U597 ( .A(KEYINPUT17), .B(n548), .Z(n900) );
  NAND2_X1 U598 ( .A1(G137), .A2(n900), .ZN(n549) );
  XNOR2_X1 U599 ( .A(n549), .B(KEYINPUT66), .ZN(n558) );
  INV_X1 U600 ( .A(G2104), .ZN(n553) );
  INV_X1 U601 ( .A(G2105), .ZN(n550) );
  NOR2_X1 U602 ( .A1(n553), .A2(n550), .ZN(n892) );
  NAND2_X1 U603 ( .A1(G113), .A2(n892), .ZN(n552) );
  NOR2_X1 U604 ( .A1(G2104), .A2(n550), .ZN(n893) );
  NAND2_X1 U605 ( .A1(G125), .A2(n893), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n556) );
  NOR2_X2 U607 ( .A1(G2105), .A2(n553), .ZN(n897) );
  NAND2_X1 U608 ( .A1(G101), .A2(n897), .ZN(n554) );
  XNOR2_X1 U609 ( .A(KEYINPUT23), .B(n554), .ZN(n555) );
  NOR2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U612 ( .A(n559), .B(KEYINPUT65), .ZN(n698) );
  BUF_X1 U613 ( .A(n698), .Z(G160) );
  AND2_X1 U614 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U615 ( .A1(G111), .A2(n892), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G135), .A2(n900), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n893), .A2(G123), .ZN(n562) );
  XOR2_X1 U619 ( .A(KEYINPUT18), .B(n562), .Z(n563) );
  NOR2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n897), .A2(G99), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n947) );
  XNOR2_X1 U623 ( .A(G2096), .B(n947), .ZN(n567) );
  OR2_X1 U624 ( .A1(G2100), .A2(n567), .ZN(G156) );
  INV_X1 U625 ( .A(G860), .ZN(n614) );
  NAND2_X1 U626 ( .A1(n649), .A2(G81), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G68), .A2(n653), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G43), .A2(n650), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n532), .A2(n572), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G56), .A2(n657), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT75), .ZN(n574) );
  XNOR2_X1 U634 ( .A(n574), .B(KEYINPUT14), .ZN(n575) );
  NOR2_X1 U635 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U636 ( .A1(n614), .A2(n1007), .ZN(G153) );
  INV_X1 U637 ( .A(G57), .ZN(G237) );
  INV_X1 U638 ( .A(G108), .ZN(G238) );
  NAND2_X1 U639 ( .A1(G89), .A2(n649), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT4), .ZN(n579) );
  XNOR2_X1 U641 ( .A(n579), .B(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G76), .A2(n653), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U644 ( .A(KEYINPUT5), .B(n582), .ZN(n588) );
  XNOR2_X1 U645 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G51), .A2(n650), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G63), .A2(n657), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n586), .B(n585), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U651 ( .A(KEYINPUT7), .B(n589), .ZN(G168) );
  XOR2_X1 U652 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U653 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n591) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G223) );
  INV_X1 U656 ( .A(G567), .ZN(n685) );
  NOR2_X1 U657 ( .A1(G223), .A2(n685), .ZN(n593) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(KEYINPUT11), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n593), .B(n592), .ZN(G234) );
  NAND2_X1 U660 ( .A1(G301), .A2(G868), .ZN(n603) );
  NAND2_X1 U661 ( .A1(G54), .A2(n650), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G92), .A2(n649), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G79), .A2(n653), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U665 ( .A1(G66), .A2(n657), .ZN(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT77), .B(n596), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U669 ( .A(n601), .B(KEYINPUT15), .ZN(n998) );
  OR2_X1 U670 ( .A1(n998), .A2(G868), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G53), .A2(n650), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G65), .A2(n657), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G91), .A2(n649), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G78), .A2(n653), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n995) );
  INV_X1 U679 ( .A(n995), .ZN(G299) );
  INV_X1 U680 ( .A(G868), .ZN(n610) );
  NOR2_X1 U681 ( .A1(G286), .A2(n610), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT80), .ZN(n613) );
  NOR2_X1 U683 ( .A1(G299), .A2(G868), .ZN(n612) );
  NOR2_X1 U684 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n615), .A2(n998), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n616), .B(KEYINPUT16), .ZN(n617) );
  XOR2_X1 U688 ( .A(KEYINPUT81), .B(n617), .Z(G148) );
  NOR2_X1 U689 ( .A1(n1007), .A2(G868), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G868), .A2(n998), .ZN(n618) );
  NOR2_X1 U691 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G559), .A2(n998), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n621), .B(n1007), .ZN(n667) );
  NOR2_X1 U695 ( .A1(G860), .A2(n667), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G55), .A2(n650), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G67), .A2(n657), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U699 ( .A1(G93), .A2(n649), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G80), .A2(n653), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n669) );
  XNOR2_X1 U703 ( .A(n628), .B(n669), .ZN(G145) );
  NAND2_X1 U704 ( .A1(G72), .A2(n653), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G47), .A2(n650), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G85), .A2(n649), .ZN(n631) );
  XNOR2_X1 U708 ( .A(KEYINPUT67), .B(n631), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n657), .A2(G60), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U712 ( .A1(G86), .A2(n649), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G48), .A2(n650), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n653), .A2(G73), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n638), .Z(n639) );
  NOR2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n657), .A2(G61), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G49), .A2(n650), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G87), .A2(n643), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U723 ( .A1(n657), .A2(n646), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G651), .A2(G74), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G88), .A2(n649), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G50), .A2(n650), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U729 ( .A1(n653), .A2(G75), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT82), .B(n654), .Z(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n657), .A2(G62), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U735 ( .A(n995), .B(G290), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n660), .B(G305), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n662) );
  XNOR2_X1 U738 ( .A(G288), .B(KEYINPUT84), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U740 ( .A(n664), .B(n663), .Z(n666) );
  XNOR2_X1 U741 ( .A(G166), .B(n669), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n666), .B(n665), .ZN(n919) );
  XNOR2_X1 U743 ( .A(n667), .B(n919), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n668), .A2(G868), .ZN(n671) );
  OR2_X1 U745 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XNOR2_X1 U748 ( .A(n672), .B(KEYINPUT85), .ZN(n673) );
  XNOR2_X1 U749 ( .A(KEYINPUT20), .B(n673), .ZN(n674) );
  NAND2_X1 U750 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(KEYINPUT22), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT86), .ZN(n679) );
  NOR2_X1 U757 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G96), .A2(n680), .ZN(n850) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n850), .ZN(n681) );
  XNOR2_X1 U760 ( .A(n681), .B(KEYINPUT87), .ZN(n687) );
  NAND2_X1 U761 ( .A1(G120), .A2(G69), .ZN(n682) );
  NOR2_X1 U762 ( .A1(G237), .A2(n682), .ZN(n683) );
  XOR2_X1 U763 ( .A(KEYINPUT88), .B(n683), .Z(n684) );
  NOR2_X1 U764 ( .A1(G238), .A2(n684), .ZN(n852) );
  NOR2_X1 U765 ( .A1(n685), .A2(n852), .ZN(n686) );
  NOR2_X1 U766 ( .A1(n687), .A2(n686), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n688) );
  XOR2_X1 U769 ( .A(KEYINPUT89), .B(n688), .Z(n689) );
  NOR2_X1 U770 ( .A1(n690), .A2(n689), .ZN(n849) );
  NAND2_X1 U771 ( .A1(n849), .A2(G36), .ZN(G176) );
  NAND2_X1 U772 ( .A1(G114), .A2(n892), .ZN(n692) );
  NAND2_X1 U773 ( .A1(G102), .A2(n897), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U775 ( .A1(G138), .A2(n900), .ZN(n693) );
  XNOR2_X1 U776 ( .A(n693), .B(KEYINPUT90), .ZN(n695) );
  NAND2_X1 U777 ( .A1(n893), .A2(G126), .ZN(n694) );
  NAND2_X1 U778 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U779 ( .A1(n697), .A2(n696), .ZN(G164) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n791) );
  NAND2_X1 U781 ( .A1(n698), .A2(G40), .ZN(n699) );
  XNOR2_X1 U782 ( .A(n699), .B(KEYINPUT91), .ZN(n790) );
  NAND2_X1 U783 ( .A1(n791), .A2(n790), .ZN(n730) );
  INV_X1 U784 ( .A(G1996), .ZN(n827) );
  NOR2_X1 U785 ( .A1(n730), .A2(n827), .ZN(n700) );
  XNOR2_X1 U786 ( .A(n700), .B(KEYINPUT26), .ZN(n702) );
  AND2_X1 U787 ( .A1(n730), .A2(G1341), .ZN(n701) );
  OR2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n709), .A2(n998), .ZN(n704) );
  INV_X1 U790 ( .A(n730), .ZN(n725) );
  INV_X1 U791 ( .A(n725), .ZN(n740) );
  NOR2_X1 U792 ( .A1(G2067), .A2(n740), .ZN(n706) );
  NOR2_X1 U793 ( .A1(n725), .A2(G1348), .ZN(n705) );
  NOR2_X1 U794 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n712) );
  XNOR2_X1 U796 ( .A(n710), .B(KEYINPUT101), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U798 ( .A1(G2072), .A2(n725), .ZN(n713) );
  XNOR2_X1 U799 ( .A(n713), .B(KEYINPUT98), .ZN(n714) );
  XNOR2_X1 U800 ( .A(n714), .B(KEYINPUT27), .ZN(n716) );
  XNOR2_X1 U801 ( .A(G1956), .B(KEYINPUT99), .ZN(n1018) );
  NOR2_X1 U802 ( .A1(n1018), .A2(n725), .ZN(n715) );
  NOR2_X1 U803 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U804 ( .A1(n995), .A2(n719), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U806 ( .A1(n995), .A2(n719), .ZN(n720) );
  XOR2_X1 U807 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n724) );
  INV_X1 U809 ( .A(G1961), .ZN(n1033) );
  NAND2_X1 U810 ( .A1(n740), .A2(n1033), .ZN(n727) );
  XNOR2_X1 U811 ( .A(KEYINPUT25), .B(G2078), .ZN(n971) );
  NAND2_X1 U812 ( .A1(n725), .A2(n971), .ZN(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n736) );
  NAND2_X1 U814 ( .A1(n736), .A2(G171), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n755) );
  INV_X1 U816 ( .A(G1966), .ZN(n732) );
  NAND2_X1 U817 ( .A1(G8), .A2(n730), .ZN(n731) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n740), .ZN(n756) );
  NOR2_X1 U819 ( .A1(n757), .A2(n756), .ZN(n733) );
  NAND2_X1 U820 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U822 ( .A1(n735), .A2(G168), .ZN(n738) );
  NOR2_X1 U823 ( .A1(G171), .A2(n736), .ZN(n737) );
  NOR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n739), .Z(n754) );
  INV_X1 U826 ( .A(G8), .ZN(n746) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n740), .ZN(n742) );
  INV_X1 U828 ( .A(n783), .ZN(n767) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n767), .ZN(n741) );
  NOR2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT102), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n744), .A2(G303), .ZN(n745) );
  OR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n748) );
  AND2_X1 U834 ( .A1(n754), .A2(n748), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n755), .A2(n747), .ZN(n752) );
  INV_X1 U836 ( .A(n748), .ZN(n750) );
  AND2_X1 U837 ( .A1(G286), .A2(G8), .ZN(n749) );
  OR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n753), .B(KEYINPUT32), .ZN(n762) );
  AND2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n760) );
  AND2_X1 U842 ( .A1(G8), .A2(n756), .ZN(n758) );
  OR2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U844 ( .A1(n762), .A2(n761), .ZN(n775) );
  NOR2_X1 U845 ( .A1(G288), .A2(G1976), .ZN(n763) );
  XOR2_X1 U846 ( .A(n763), .B(KEYINPUT103), .Z(n782) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n764) );
  NOR2_X1 U848 ( .A1(n782), .A2(n764), .ZN(n1002) );
  NAND2_X1 U849 ( .A1(n775), .A2(n1002), .ZN(n765) );
  XNOR2_X1 U850 ( .A(n765), .B(KEYINPUT104), .ZN(n769) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U852 ( .A(n994), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U855 ( .A(n770), .B(KEYINPUT64), .ZN(n781) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  AND2_X1 U858 ( .A1(n772), .A2(n783), .ZN(n787) );
  OR2_X1 U859 ( .A1(KEYINPUT33), .A2(n787), .ZN(n779) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(KEYINPUT105), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n746), .A2(n774), .ZN(n777) );
  INV_X1 U863 ( .A(n775), .ZN(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U865 ( .A1(n783), .A2(n778), .ZN(n789) );
  OR2_X1 U866 ( .A1(n779), .A2(n789), .ZN(n780) );
  XNOR2_X1 U867 ( .A(G1981), .B(G305), .ZN(n991) );
  AND2_X1 U868 ( .A1(n782), .A2(KEYINPUT33), .ZN(n784) );
  AND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n991), .A2(n785), .ZN(n786) );
  OR2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n813) );
  INV_X1 U873 ( .A(n790), .ZN(n792) );
  NOR2_X1 U874 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U875 ( .A(n793), .B(KEYINPUT92), .ZN(n839) );
  INV_X1 U876 ( .A(n839), .ZN(n811) );
  NAND2_X1 U877 ( .A1(G105), .A2(n897), .ZN(n794) );
  XNOR2_X1 U878 ( .A(n794), .B(KEYINPUT38), .ZN(n801) );
  NAND2_X1 U879 ( .A1(G117), .A2(n892), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G141), .A2(n900), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G129), .A2(n893), .ZN(n797) );
  XNOR2_X1 U883 ( .A(KEYINPUT95), .B(n797), .ZN(n798) );
  NOR2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U886 ( .A(KEYINPUT96), .B(n802), .Z(n888) );
  NOR2_X1 U887 ( .A1(n827), .A2(n888), .ZN(n810) );
  NAND2_X1 U888 ( .A1(G95), .A2(n897), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G131), .A2(n900), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G107), .A2(n892), .ZN(n806) );
  NAND2_X1 U892 ( .A1(G119), .A2(n893), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n910) );
  INV_X1 U895 ( .A(G1991), .ZN(n964) );
  NOR2_X1 U896 ( .A1(n910), .A2(n964), .ZN(n809) );
  NOR2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n946) );
  NOR2_X1 U898 ( .A1(n811), .A2(n946), .ZN(n831) );
  INV_X1 U899 ( .A(n831), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n813), .A2(n812), .ZN(n826) );
  XOR2_X1 U901 ( .A(G1986), .B(G290), .Z(n996) );
  XNOR2_X1 U902 ( .A(G2067), .B(KEYINPUT37), .ZN(n837) );
  NAND2_X1 U903 ( .A1(n892), .A2(G116), .ZN(n814) );
  XNOR2_X1 U904 ( .A(n814), .B(KEYINPUT94), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G128), .A2(n893), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U907 ( .A(n817), .B(KEYINPUT35), .ZN(n823) );
  XNOR2_X1 U908 ( .A(KEYINPUT34), .B(KEYINPUT93), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G104), .A2(n897), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G140), .A2(n900), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U914 ( .A(KEYINPUT36), .B(n824), .Z(n890) );
  NOR2_X1 U915 ( .A1(n837), .A2(n890), .ZN(n835) );
  INV_X1 U916 ( .A(n835), .ZN(n952) );
  NAND2_X1 U917 ( .A1(n996), .A2(n952), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n534), .A2(n533), .ZN(n842) );
  AND2_X1 U919 ( .A1(n827), .A2(n888), .ZN(n943) );
  AND2_X1 U920 ( .A1(n964), .A2(n910), .ZN(n950) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n828) );
  XNOR2_X1 U922 ( .A(KEYINPUT106), .B(n828), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n950), .A2(n829), .ZN(n830) );
  NOR2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U925 ( .A1(n943), .A2(n832), .ZN(n833) );
  XOR2_X1 U926 ( .A(KEYINPUT39), .B(n833), .Z(n834) );
  NOR2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U928 ( .A(n836), .B(KEYINPUT107), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n837), .A2(n890), .ZN(n954) );
  NAND2_X1 U930 ( .A1(n838), .A2(n954), .ZN(n840) );
  NAND2_X1 U931 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U933 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U934 ( .A(G223), .ZN(n844) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n844), .ZN(G217) );
  INV_X1 U936 ( .A(G661), .ZN(n846) );
  NAND2_X1 U937 ( .A1(G2), .A2(G15), .ZN(n845) );
  NOR2_X1 U938 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(n847), .Z(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U943 ( .A(G132), .ZN(G219) );
  INV_X1 U944 ( .A(G120), .ZN(G236) );
  INV_X1 U945 ( .A(G82), .ZN(G220) );
  INV_X1 U946 ( .A(G69), .ZN(G235) );
  INV_X1 U947 ( .A(n850), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(G261) );
  INV_X1 U949 ( .A(G261), .ZN(G325) );
  XOR2_X1 U950 ( .A(KEYINPUT42), .B(G2090), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(G2100), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(G2096), .B(KEYINPUT43), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2678), .B(KEYINPUT109), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(G227) );
  XNOR2_X1 U960 ( .A(G1981), .B(G2474), .ZN(n871) );
  XOR2_X1 U961 ( .A(G1956), .B(G1961), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1986), .B(G1966), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U964 ( .A(G1976), .B(G1971), .Z(n865) );
  XNOR2_X1 U965 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U968 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U971 ( .A1(n897), .A2(G100), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n872), .Z(n874) );
  NAND2_X1 U973 ( .A1(n892), .A2(G112), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(KEYINPUT112), .B(n875), .ZN(n880) );
  NAND2_X1 U976 ( .A1(n893), .A2(G124), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT44), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G136), .A2(n900), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U980 ( .A1(n880), .A2(n879), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G118), .A2(n892), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G130), .A2(n893), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G106), .A2(n897), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G142), .A2(n900), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U987 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n914) );
  XOR2_X1 U990 ( .A(G160), .B(n890), .Z(n891) );
  XNOR2_X1 U991 ( .A(n891), .B(G162), .ZN(n906) );
  NAND2_X1 U992 ( .A1(G115), .A2(n892), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G127), .A2(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(KEYINPUT47), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G103), .A2(n897), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n900), .A2(G139), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT114), .B(n901), .Z(n902) );
  NOR2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n938) );
  XOR2_X1 U1001 ( .A(G164), .B(n938), .Z(n904) );
  XNOR2_X1 U1002 ( .A(n947), .B(n904), .ZN(n905) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n912) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n908) );
  XNOR2_X1 U1005 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n914), .B(n913), .Z(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G395) );
  XOR2_X1 U1011 ( .A(G286), .B(n1007), .Z(n917) );
  XNOR2_X1 U1012 ( .A(G301), .B(n998), .ZN(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n919), .B(n918), .Z(n920) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n920), .ZN(G397) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n922), .B(n921), .ZN(n933) );
  XOR2_X1 U1019 ( .A(G2451), .B(G2430), .Z(n924) );
  XNOR2_X1 U1020 ( .A(G2438), .B(G2443), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n924), .B(n923), .ZN(n930) );
  XOR2_X1 U1022 ( .A(G2435), .B(G2454), .Z(n926) );
  XNOR2_X1 U1023 ( .A(G1348), .B(G1341), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n926), .B(n925), .ZN(n928) );
  XOR2_X1 U1025 ( .A(G2446), .B(G2427), .Z(n927) );
  XNOR2_X1 U1026 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(n930), .B(n929), .Z(n931) );
  NAND2_X1 U1028 ( .A1(G14), .A2(n931), .ZN(n936) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n936), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G96), .ZN(G221) );
  INV_X1 U1035 ( .A(n936), .ZN(G401) );
  XNOR2_X1 U1036 ( .A(G164), .B(G2078), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT119), .ZN(n940) );
  XOR2_X1 U1038 ( .A(G2072), .B(n938), .Z(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT50), .B(n941), .Z(n960) );
  XOR2_X1 U1041 ( .A(G2090), .B(G162), .Z(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1043 ( .A(KEYINPUT51), .B(n944), .Z(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n957) );
  XNOR2_X1 U1045 ( .A(G160), .B(G2084), .ZN(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT117), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1052 ( .A(KEYINPUT118), .B(n958), .Z(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n961), .ZN(n962) );
  INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n986) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n986), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(G29), .ZN(n1046) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G35), .ZN(n981) );
  XNOR2_X1 U1059 ( .A(n964), .B(G25), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n965), .A2(G28), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n966), .B(KEYINPUT120), .ZN(n978) );
  XNOR2_X1 U1062 ( .A(KEYINPUT121), .B(G2072), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(n967), .B(G33), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G1996), .B(G32), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(n968), .B(KEYINPUT123), .ZN(n970) );
  XOR2_X1 U1066 ( .A(G2067), .B(G26), .Z(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n974) );
  XOR2_X1 U1068 ( .A(G27), .B(n971), .Z(n972) );
  XNOR2_X1 U1069 ( .A(KEYINPUT122), .B(n972), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT53), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G2084), .B(KEYINPUT54), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G34), .B(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n988) );
  INV_X1 U1079 ( .A(G29), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n989), .ZN(n1044) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1013) );
  XOR2_X1 U1083 ( .A(G168), .B(G1966), .Z(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n992), .Z(n1011) );
  XNOR2_X1 U1086 ( .A(G301), .B(n1033), .ZN(n1006) );
  NAND2_X1 U1087 ( .A1(G1971), .A2(G303), .ZN(n993) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(n995), .B(G1956), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1091 ( .A(G1348), .B(n998), .Z(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G1341), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1042) );
  INV_X1 U1100 ( .A(G16), .ZN(n1040) );
  XNOR2_X1 U1101 ( .A(KEYINPUT59), .B(G1348), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(n1014), .B(G4), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(G1341), .B(G19), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(G1981), .B(G6), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1106 ( .A(KEYINPUT124), .B(n1017), .Z(n1020) );
  XOR2_X1 U1107 ( .A(n1018), .B(G20), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(KEYINPUT60), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1024), .B(KEYINPUT125), .ZN(n1032) );
  XOR2_X1 U1112 ( .A(G1971), .B(KEYINPUT126), .Z(n1025) );
  XNOR2_X1 U1113 ( .A(G22), .B(n1025), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(G1986), .B(G24), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(G23), .B(G1976), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1118 ( .A(KEYINPUT58), .B(n1030), .Z(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1037) );
  XOR2_X1 U1120 ( .A(G1966), .B(G21), .Z(n1035) );
  XNOR2_X1 U1121 ( .A(n1033), .B(G5), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(KEYINPUT61), .B(n1038), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1127 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1128 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1047), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

