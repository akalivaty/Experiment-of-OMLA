//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G1gat), .B2(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n214), .C1(G1gat), .C2(new_n208), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT91), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n218), .B2(KEYINPUT14), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G43gat), .ZN(new_n224));
  INV_X1    g023(.A(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G43gat), .A2(G50gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT15), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n231), .A3(new_n227), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n226), .A2(KEYINPUT89), .A3(new_n231), .A4(new_n227), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n234), .A2(new_n223), .A3(new_n229), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n230), .A2(new_n236), .A3(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n236), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n236), .A3(KEYINPUT90), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n217), .A2(new_n237), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(new_n216), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT92), .Z(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT18), .A4(new_n250), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n250), .B(KEYINPUT13), .Z(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n246), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n207), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n251), .A2(new_n252), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(new_n206), .A3(new_n254), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT34), .ZN(new_n265));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT65), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(KEYINPUT23), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n274), .A2(G169gat), .A3(G176gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  OAI211_X1 g077(.A(KEYINPUT65), .B(new_n277), .C1(new_n278), .C2(new_n271), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n280), .B(new_n283), .C1(new_n285), .C2(KEYINPUT24), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT67), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT68), .B(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n282), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n280), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n273), .A2(new_n298), .A3(new_n275), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n291), .A2(new_n292), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n285), .B1(KEYINPUT26), .B2(new_n271), .ZN(new_n302));
  INV_X1    g101(.A(new_n272), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n306));
  AOI21_X1  g105(.A(G190gat), .B1(new_n306), .B2(KEYINPUT69), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n281), .A2(KEYINPUT68), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(KEYINPUT27), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n311), .A3(KEYINPUT70), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT28), .A3(new_n282), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n305), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT71), .B(G134gat), .Z(new_n323));
  INV_X1    g122(.A(G127gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G134gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n325), .A2(new_n328), .B1(KEYINPUT1), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT74), .B1(new_n332), .B2(G113gat), .ZN(new_n333));
  AND2_X1   g132(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n333), .B1(new_n336), .B2(G113gat), .ZN(new_n337));
  INV_X1    g136(.A(G113gat), .ZN(new_n338));
  NOR4_X1   g137(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT74), .A4(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n331), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n335), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g141(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n341), .A2(new_n342), .A3(G113gat), .A4(new_n343), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n344), .B(KEYINPUT75), .C1(new_n345), .C2(new_n333), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n324), .A2(new_n327), .ZN(new_n347));
  NAND2_X1  g146(.A1(G127gat), .A2(G134gat), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT1), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n340), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n322), .A2(new_n330), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n330), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n301), .A2(new_n352), .A3(new_n321), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n269), .B1(new_n354), .B2(new_n266), .ZN(new_n355));
  INV_X1    g154(.A(new_n266), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n356), .B(new_n268), .C1(new_n351), .C2(new_n353), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n356), .A3(new_n353), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n360), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n368), .A2(KEYINPUT33), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(KEYINPUT32), .A3(new_n370), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n358), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n357), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n266), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n268), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n367), .A2(new_n371), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT36), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n367), .A2(new_n371), .ZN(new_n379));
  INV_X1    g178(.A(new_n358), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n358), .A2(new_n367), .A3(new_n371), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT36), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n378), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G22gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT22), .ZN(new_n388));
  INV_X1    g187(.A(G211gat), .ZN(new_n389));
  INV_X1    g188(.A(G218gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT78), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G211gat), .B(G218gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n396), .A2(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n387), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  XNOR2_X1  g202(.A(G141gat), .B(G148gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(G155gat), .B2(G162gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G155gat), .B(G162gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n412));
  OR2_X1    g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(new_n403), .A3(new_n408), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n415), .A2(new_n403), .A3(new_n408), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n408), .B1(new_n415), .B2(new_n403), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n387), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(KEYINPUT83), .A3(new_n387), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XOR2_X1   g225(.A(G211gat), .B(G218gat), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT79), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(new_n392), .A3(new_n394), .A4(new_n395), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n397), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n396), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n386), .B(new_n419), .C1(new_n426), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n399), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n435), .B2(new_n387), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n424), .A2(new_n425), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n399), .ZN(new_n438));
  INV_X1    g237(.A(new_n433), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n385), .B(new_n434), .C1(new_n440), .C2(new_n386), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n426), .A2(new_n433), .ZN(new_n444));
  OAI211_X1 g243(.A(G228gat), .B(G233gat), .C1(new_n444), .C2(new_n436), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n385), .B1(new_n445), .B2(new_n434), .ZN(new_n446));
  OAI21_X1  g245(.A(G78gat), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n434), .B1(new_n440), .B2(new_n386), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(G78gat), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n442), .A3(new_n450), .A4(new_n441), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT31), .B(G50gat), .Z(new_n452));
  XNOR2_X1  g251(.A(new_n452), .B(G106gat), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n447), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n447), .B2(new_n451), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n352), .A2(KEYINPUT82), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n350), .A2(new_n459), .A3(new_n330), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n418), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n350), .A2(new_n417), .A3(new_n330), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G225gat), .A2(G233gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n457), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n420), .A2(new_n421), .A3(new_n387), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n424), .B2(new_n425), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n458), .A3(new_n460), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n462), .A2(KEYINPUT4), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n350), .A2(new_n471), .A3(new_n417), .A4(new_n330), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n473), .A3(new_n464), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n464), .B1(new_n461), .B2(new_n462), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT84), .B(new_n474), .C1(new_n477), .C2(new_n457), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT87), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT0), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n461), .A2(new_n464), .A3(new_n462), .ZN(new_n489));
  INV_X1    g288(.A(new_n460), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n459), .B1(new_n350), .B2(new_n330), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n492), .A2(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT39), .B(new_n489), .C1(new_n493), .C2(new_n464), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n464), .B1(new_n469), .B2(new_n473), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT39), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n488), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT40), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT40), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n483), .A2(new_n488), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n287), .A2(KEYINPUT66), .A3(new_n288), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT66), .B1(new_n287), .B2(new_n288), .ZN(new_n510));
  INV_X1    g309(.A(new_n300), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT80), .B1(new_n512), .B2(new_n320), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT80), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n301), .A2(new_n514), .A3(new_n321), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n513), .A2(new_n515), .A3(G226gat), .A4(G233gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(G226gat), .A2(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n399), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n322), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n516), .A2(new_n520), .A3(new_n439), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n301), .A2(new_n514), .A3(new_n321), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n514), .B1(new_n301), .B2(new_n321), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n322), .A2(new_n517), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n439), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n508), .B1(new_n521), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(new_n520), .A3(new_n439), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n515), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n530), .B2(new_n519), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n529), .B(new_n507), .C1(new_n531), .C2(new_n439), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(KEYINPUT30), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n527), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(new_n529), .A3(new_n535), .A4(new_n507), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n456), .B1(new_n504), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n476), .A2(new_n478), .A3(new_n488), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n476), .A2(new_n481), .A3(new_n478), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n481), .B1(new_n476), .B2(new_n478), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n488), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT6), .B1(new_n479), .B2(new_n487), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n508), .A2(KEYINPUT37), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT38), .B1(new_n528), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n439), .A3(new_n526), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n439), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n516), .A2(new_n520), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n433), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT37), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n529), .B1(new_n531), .B2(new_n439), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n508), .B1(new_n558), .B2(KEYINPUT37), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT37), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n534), .B2(new_n529), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT38), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n532), .A3(new_n557), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n384), .B1(new_n538), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n545), .A2(new_n539), .ZN(new_n565));
  INV_X1    g364(.A(new_n541), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n565), .A2(new_n566), .B1(new_n533), .B2(new_n536), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n454), .A2(new_n455), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n381), .A2(new_n382), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n456), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT35), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n546), .A2(new_n456), .A3(new_n570), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n537), .A2(KEYINPUT35), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n264), .B1(new_n569), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G57gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G64gat), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(G57gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n580), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR3_X1   g390(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n580), .A2(new_n582), .ZN(new_n593));
  OAI221_X1 g392(.A(new_n584), .B1(new_n591), .B2(new_n592), .C1(new_n593), .C2(new_n583), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n216), .B1(new_n595), .B2(KEYINPUT21), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT97), .Z(new_n597));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT96), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(KEYINPUT95), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n611), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n606), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n612), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n602), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n613), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(new_n617), .A3(new_n601), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n245), .ZN(new_n630));
  NAND2_X1  g429(.A1(G85gat), .A2(G92gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT7), .ZN(new_n632));
  XNOR2_X1  g431(.A(G99gat), .B(G106gat), .ZN(new_n633));
  NOR2_X1   g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(KEYINPUT8), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n632), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n633), .B1(new_n632), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n630), .A2(new_n639), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n637), .A2(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n243), .A2(new_n237), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n640), .B2(new_n644), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n629), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n628), .A3(new_n645), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n624), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n633), .A2(KEYINPUT98), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n589), .A2(new_n594), .A3(new_n639), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n587), .A2(new_n588), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT94), .B1(new_n585), .B2(new_n586), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n594), .B(new_n654), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n643), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n594), .A4(new_n639), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n655), .A2(new_n659), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n668), .A3(new_n672), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n653), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n578), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n541), .B1(new_n545), .B2(new_n539), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT99), .B(G1gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1324gat));
  NAND3_X1  g482(.A1(new_n578), .A2(new_n537), .A3(new_n677), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT100), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(G8gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(G1325gat));
  OR2_X1    g490(.A1(new_n378), .A2(new_n383), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n678), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n570), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n678), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n568), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NOR3_X1   g497(.A1(new_n624), .A2(new_n652), .A3(new_n676), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n680), .A2(G29gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n578), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT101), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  AOI22_X1  g503(.A1(KEYINPUT35), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n487), .B1(new_n480), .B2(new_n482), .ZN(new_n706));
  INV_X1    g505(.A(new_n545), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n566), .B(new_n532), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n528), .A2(new_n547), .B1(KEYINPUT37), .B2(new_n558), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT38), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n549), .A2(new_n550), .B1(new_n553), .B2(new_n433), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n560), .B1(new_n711), .B2(new_n552), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n710), .B(new_n508), .C1(new_n558), .C2(KEYINPUT37), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n709), .A2(new_n710), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n502), .A2(new_n503), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n716), .A2(new_n536), .A3(new_n533), .A4(new_n544), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n568), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n692), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT103), .B1(new_n567), .B2(new_n568), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n721), .B(new_n456), .C1(new_n537), .C2(new_n679), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT104), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n564), .A2(new_n725), .A3(new_n722), .A4(new_n720), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n705), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n648), .A2(new_n650), .A3(KEYINPUT105), .ZN(new_n728));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n648), .B2(new_n650), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n704), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n569), .A2(new_n577), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n263), .B(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n624), .A2(new_n676), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n680), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n703), .A2(new_n740), .ZN(G1328gat));
  INV_X1    g540(.A(new_n537), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n578), .A2(new_n699), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n537), .A2(new_n221), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n744), .A2(KEYINPUT106), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n743), .A2(new_n750), .ZN(G1329gat));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n384), .A3(new_n734), .A4(new_n738), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n570), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n578), .A2(new_n224), .A3(new_n756), .A4(new_n699), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n753), .B(new_n757), .C1(new_n754), .C2(KEYINPUT47), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1330gat));
  NOR2_X1   g561(.A1(new_n568), .A2(new_n225), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n735), .A2(new_n738), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n225), .B1(new_n746), .B2(new_n568), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT48), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1331gat));
  NAND2_X1  g569(.A1(new_n724), .A2(new_n726), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n577), .ZN(new_n772));
  INV_X1    g571(.A(new_n676), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n263), .B(KEYINPUT102), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n653), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n680), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(new_n579), .ZN(G1332gat));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n742), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  AND2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n779), .B2(new_n780), .ZN(G1333gat));
  OAI21_X1  g582(.A(G71gat), .B1(new_n776), .B2(new_n692), .ZN(new_n784));
  INV_X1    g583(.A(G71gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n756), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n776), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1334gat));
  NOR2_X1   g588(.A1(new_n776), .A2(new_n568), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(new_n450), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n624), .A2(new_n774), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n676), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n735), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795), .B2(new_n680), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n651), .A4(new_n792), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n792), .A2(new_n651), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n727), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OR3_X1    g601(.A1(new_n680), .A2(G85gat), .A3(new_n773), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NAND4_X1  g603(.A1(new_n732), .A2(new_n537), .A3(new_n734), .A4(new_n794), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G92gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n742), .A2(G92gat), .A3(new_n773), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n795), .B2(new_n692), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n570), .A2(G99gat), .A3(new_n773), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n802), .B2(new_n815), .ZN(G1338gat));
  NAND4_X1  g615(.A1(new_n732), .A2(new_n456), .A3(new_n734), .A4(new_n794), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n568), .A2(G106gat), .A3(new_n773), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n820), .B(KEYINPUT108), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n817), .A2(G106gat), .B1(new_n801), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n819), .B2(new_n824), .ZN(G1339gat));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n624), .A2(new_n652), .A3(new_n773), .A4(new_n737), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n661), .A2(new_n667), .A3(new_n662), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n663), .A2(new_n830), .A3(new_n664), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n831), .A2(KEYINPUT109), .A3(new_n673), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT109), .B1(new_n831), .B2(new_n673), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n675), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT55), .B(new_n829), .C1(new_n832), .C2(new_n833), .ZN(new_n838));
  INV_X1    g637(.A(new_n255), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n248), .A2(new_n256), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT110), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n250), .B1(new_n244), .B2(new_n248), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n205), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n262), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n837), .A2(new_n730), .A3(new_n838), .A4(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n676), .A3(new_n262), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n837), .A2(new_n838), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n737), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n731), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n827), .B1(new_n850), .B2(new_n624), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n680), .A2(new_n456), .A3(new_n570), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n826), .B1(new_n853), .B2(new_n537), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n851), .A2(KEYINPUT111), .A3(new_n742), .A4(new_n852), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n338), .A3(new_n264), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n742), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n774), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n857), .B1(new_n862), .B2(new_n338), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n856), .B2(new_n773), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n676), .A2(new_n336), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n860), .B2(new_n865), .ZN(G1341gat));
  NAND2_X1  g665(.A1(new_n620), .A2(new_n623), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n326), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n326), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n860), .B2(new_n869), .ZN(G1342gat));
  OR2_X1    g669(.A1(new_n652), .A2(new_n323), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n860), .A2(new_n871), .B1(new_n872), .B2(KEYINPUT56), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(KEYINPUT114), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n872), .B(KEYINPUT56), .C1(new_n860), .C2(new_n871), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n854), .A2(new_n651), .A3(new_n855), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(KEYINPUT113), .A3(G134gat), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT113), .B1(new_n877), .B2(G134gat), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n875), .B(new_n876), .C1(new_n878), .C2(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n384), .A2(new_n680), .A3(new_n537), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n568), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n867), .A2(new_n774), .A3(new_n651), .A4(new_n676), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n836), .A2(new_n263), .A3(new_n675), .A4(new_n838), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n651), .B1(new_n888), .B2(new_n847), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n845), .B1(new_n889), .B2(KEYINPUT115), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n891));
  AOI211_X1 g690(.A(new_n891), .B(new_n651), .C1(new_n888), .C2(new_n847), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n867), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT116), .B(new_n867), .C1(new_n890), .C2(new_n892), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n851), .B2(new_n456), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n774), .B(new_n883), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n264), .A2(G141gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n851), .A2(new_n456), .A3(new_n883), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n882), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT58), .B1(new_n902), .B2(KEYINPUT117), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n774), .A2(new_n838), .A3(new_n837), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n730), .B1(new_n905), .B2(new_n847), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n867), .B1(new_n906), .B2(new_n846), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n568), .B1(new_n907), .B2(new_n827), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n883), .A4(new_n901), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n263), .B(new_n883), .C1(new_n897), .C2(new_n898), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(G141gat), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n881), .B1(new_n903), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(G141gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n910), .A3(new_n904), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n908), .A2(new_n883), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n899), .A2(G141gat), .B1(new_n917), .B2(new_n901), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n916), .B(KEYINPUT118), .C1(new_n882), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n914), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(G148gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n921), .A3(new_n676), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  AND4_X1   g722(.A1(new_n651), .A2(new_n837), .A3(new_n838), .A4(new_n844), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(new_n889), .ZN(new_n925));
  AOI22_X1  g724(.A1(new_n677), .A2(new_n264), .B1(new_n867), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n884), .B1(new_n926), .B2(new_n568), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n851), .A2(new_n885), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT119), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n851), .A2(new_n930), .A3(new_n885), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n676), .A3(new_n883), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n923), .B1(new_n933), .B2(G148gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n935), .A2(new_n773), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(KEYINPUT59), .A3(new_n921), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n922), .B1(new_n934), .B2(new_n937), .ZN(G1345gat));
  INV_X1    g737(.A(G155gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n624), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(KEYINPUT120), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(KEYINPUT120), .B2(new_n940), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n935), .A2(new_n939), .A3(new_n867), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  OAI21_X1  g743(.A(G162gat), .B1(new_n935), .B2(new_n731), .ZN(new_n945));
  INV_X1    g744(.A(G162gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n917), .A2(new_n946), .A3(new_n651), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT121), .ZN(G1347gat));
  NAND2_X1  g748(.A1(new_n851), .A2(new_n680), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n742), .A2(new_n570), .A3(new_n456), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n737), .A2(G169gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(KEYINPUT123), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n680), .A2(new_n537), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT124), .Z(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(new_n571), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n851), .A3(new_n263), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(G169gat), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n956), .B1(new_n955), .B2(new_n962), .ZN(G1348gat));
  NAND2_X1  g762(.A1(new_n960), .A2(new_n851), .ZN(new_n964));
  INV_X1    g763(.A(G176gat), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n964), .A2(new_n965), .A3(new_n773), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n952), .A2(new_n676), .A3(new_n953), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(new_n965), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n965), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n966), .B1(new_n970), .B2(new_n971), .ZN(G1349gat));
  NOR2_X1   g771(.A1(new_n964), .A2(new_n867), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(new_n295), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n953), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n624), .A2(new_n318), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT60), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT60), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n974), .B(new_n979), .C1(new_n975), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1350gat));
  OAI21_X1  g780(.A(G190gat), .B1(new_n964), .B2(new_n652), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n730), .A2(new_n282), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n975), .B2(new_n984), .ZN(G1351gat));
  NOR3_X1   g784(.A1(new_n384), .A2(new_n742), .A3(new_n568), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n952), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  XOR2_X1   g787(.A(KEYINPUT126), .B(G197gat), .Z(new_n989));
  NAND3_X1  g788(.A1(new_n988), .A2(new_n774), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n959), .A2(new_n692), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n991), .B(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n932), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n993), .A2(new_n264), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n994), .B2(new_n989), .ZN(G1352gat));
  NOR2_X1   g794(.A1(new_n773), .A2(G204gat), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  OR3_X1    g796(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n932), .A2(new_n676), .A3(new_n992), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(G204gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(KEYINPUT62), .B1(new_n987), .B2(new_n997), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n988), .A2(new_n389), .A3(new_n624), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n932), .A2(new_n624), .A3(new_n992), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(G218gat), .B1(new_n993), .B2(new_n652), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n730), .A2(new_n390), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n987), .B2(new_n1009), .ZN(G1355gat));
endmodule


