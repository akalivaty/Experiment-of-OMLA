//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n202));
  XNOR2_X1  g001(.A(G155gat), .B(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n203), .A2(new_n206), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n212), .A3(new_n210), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n202), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n211), .A2(new_n217), .A3(new_n219), .ZN(new_n221));
  OR2_X1    g020(.A1(G127gat), .A2(G134gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n223), .A2(KEYINPUT69), .B1(G127gat), .B2(G134gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G113gat), .B(G120gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n222), .B(new_n224), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g025(.A(G120gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G113gat), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G120gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT1), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(KEYINPUT69), .ZN(new_n232));
  NAND2_X1  g031(.A1(G127gat), .A2(G134gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n222), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n217), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n226), .A2(new_n235), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n218), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT4), .B1(new_n236), .B2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n236), .B(new_n238), .ZN(new_n248));
  INV_X1    g047(.A(new_n241), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n252));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT0), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n247), .B2(new_n250), .ZN(new_n261));
  AOI211_X1 g060(.A(new_n202), .B(new_n219), .C1(new_n211), .C2(new_n217), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n221), .A2(new_n236), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n264), .A2(new_n220), .B1(new_n245), .B2(new_n244), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT5), .B1(new_n265), .B2(new_n241), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n256), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n252), .A2(KEYINPUT6), .A3(new_n257), .A4(new_n259), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n261), .A2(new_n266), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT6), .A4(new_n257), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n269), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT35), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277));
  AND3_X1   g076(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(G169gat), .B2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n277), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n285), .A2(G169gat), .A3(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n287), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n287), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n282), .A2(new_n283), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n277), .B1(new_n295), .B2(new_n285), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n299), .B1(new_n298), .B2(new_n300), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n289), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT27), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G183gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n314), .A3(new_n309), .ZN(new_n315));
  AND2_X1   g114(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(new_n282), .A3(new_n283), .A4(KEYINPUT68), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n287), .A2(new_n321), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n295), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n327), .A3(new_n298), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n236), .ZN(new_n330));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT64), .Z(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n306), .A2(new_n328), .A3(new_n242), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT34), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n306), .A2(new_n328), .A3(new_n242), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n242), .B1(new_n306), .B2(new_n328), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT33), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G15gat), .B(G43gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n340), .B(KEYINPUT32), .C1(new_n342), .C2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n337), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n335), .A2(KEYINPUT34), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n335), .A2(KEYINPUT34), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n347), .A2(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G204gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G197gat), .ZN(new_n356));
  INV_X1    g155(.A(G197gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G204gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT22), .ZN(new_n359));
  AND2_X1   g158(.A1(G211gat), .A2(G218gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G211gat), .A2(G218gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT71), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(KEYINPUT71), .A3(new_n362), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n366), .A2(new_n356), .A3(new_n370), .A4(new_n358), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n364), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n329), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n374), .B1(new_n306), .B2(new_n328), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n329), .A2(new_n375), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n306), .B2(new_n328), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n380), .B(new_n372), .C1(new_n375), .C2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(KEYINPUT72), .ZN(new_n384));
  XOR2_X1   g183(.A(G64gat), .B(G92gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT73), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n379), .A2(KEYINPUT73), .A3(new_n382), .A4(new_n386), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n379), .B2(new_n382), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n379), .A2(new_n382), .A3(new_n386), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n393), .B1(new_n394), .B2(KEYINPUT30), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401));
  INV_X1    g200(.A(G50gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(KEYINPUT77), .B(KEYINPUT31), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT80), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n221), .A2(new_n409), .A3(new_n376), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n221), .B2(new_n376), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n373), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n365), .A2(new_n371), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n376), .B1(new_n414), .B2(new_n363), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n219), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n416), .B2(new_n238), .ZN(new_n417));
  AOI211_X1 g216(.A(KEYINPUT79), .B(new_n218), .C1(new_n415), .C2(new_n219), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n408), .B(new_n412), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n359), .A2(KEYINPUT78), .A3(new_n362), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n371), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT78), .B1(new_n359), .B2(new_n362), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n376), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n219), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n238), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n221), .A2(new_n376), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n373), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n408), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n419), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n419), .B2(new_n429), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n406), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT82), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n436), .B(new_n406), .C1(new_n432), .C2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n408), .ZN(new_n439));
  INV_X1    g238(.A(new_n418), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n238), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n443), .B2(new_n428), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n419), .A2(new_n429), .A3(G22gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n405), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n435), .A2(new_n437), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n276), .A2(new_n354), .A3(new_n400), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n437), .A2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n430), .B1(new_n443), .B2(new_n428), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n419), .A2(new_n429), .A3(new_n431), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n436), .B1(new_n452), .B2(new_n406), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n354), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n396), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n269), .A2(new_n271), .A3(new_n274), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT35), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n350), .B2(new_n353), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n347), .A2(new_n349), .ZN(new_n463));
  INV_X1    g262(.A(new_n337), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n337), .A2(new_n347), .A3(new_n349), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n449), .A2(new_n453), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n379), .A2(new_n472), .A3(new_n382), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT85), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n379), .A2(new_n475), .A3(new_n382), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n379), .A2(new_n382), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n386), .B1(new_n478), .B2(KEYINPUT37), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT38), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n477), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n389), .A2(new_n390), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(new_n269), .A3(new_n271), .A4(new_n274), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n447), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n248), .A2(new_n249), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(KEYINPUT39), .C1(new_n265), .C2(new_n241), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n240), .A2(new_n246), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n249), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n256), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT84), .A2(KEYINPUT40), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n260), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n397), .A2(new_n498), .A3(new_n399), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n471), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n459), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G134gat), .B(G162gat), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n502), .B(KEYINPUT97), .Z(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n505));
  NAND2_X1  g304(.A1(G85gat), .A2(G92gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT7), .ZN(new_n507));
  XOR2_X1   g306(.A(G99gat), .B(G106gat), .Z(new_n508));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509));
  INV_X1    g308(.A(G85gat), .ZN(new_n510));
  INV_X1    g309(.A(G92gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(KEYINPUT8), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n508), .B1(new_n507), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n505), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n515), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT98), .A3(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT15), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  INV_X1    g325(.A(G36gat), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT87), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(G29gat), .A3(G36gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT14), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT88), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n534), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n524), .A4(new_n522), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(KEYINPUT15), .A3(new_n523), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n540), .A2(KEYINPUT89), .A3(KEYINPUT17), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT17), .B1(new_n540), .B2(KEYINPUT89), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n519), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n516), .A3(new_n518), .ZN(new_n544));
  INV_X1    g343(.A(G232gat), .ZN(new_n545));
  INV_X1    g344(.A(G233gat), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n544), .A2(KEYINPUT99), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT99), .B1(new_n544), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT100), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n543), .B(new_n554), .C1(new_n550), .C2(new_n551), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n547), .A2(KEYINPUT41), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT96), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n560), .B1(new_n556), .B2(new_n557), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n504), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n563), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n503), .A3(new_n561), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT20), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G57gat), .B(G64gat), .Z(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  AND2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n576), .A2(new_n575), .A3(KEYINPUT9), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n578), .A2(new_n579), .B1(KEYINPUT91), .B2(new_n576), .ZN(new_n580));
  XNOR2_X1  g379(.A(G71gat), .B(G78gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT93), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n581), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n573), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n583), .A2(new_n589), .A3(new_n586), .A4(new_n572), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n591));
  AND3_X1   g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n571), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(new_n590), .ZN(new_n595));
  INV_X1    g394(.A(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n570), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT16), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(G1gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(G15gat), .B(G22gat), .ZN(new_n602));
  MUX2_X1   g401(.A(G1gat), .B(new_n601), .S(new_n602), .Z(new_n603));
  INV_X1    g402(.A(G8gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT95), .Z(new_n607));
  AND3_X1   g406(.A1(new_n594), .A2(new_n599), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n594), .B2(new_n599), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n568), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n599), .ZN(new_n611));
  INV_X1    g410(.A(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n599), .A3(new_n607), .ZN(new_n614));
  INV_X1    g413(.A(new_n568), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n567), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n501), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n583), .A2(new_n586), .A3(new_n517), .A4(new_n513), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n507), .A2(new_n512), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT101), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n508), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n582), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(KEYINPUT103), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT102), .B1(new_n624), .B2(new_n626), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n628), .B(new_n625), .C1(new_n619), .C2(new_n623), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n636), .A3(new_n623), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n516), .A4(new_n518), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n626), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(new_n635), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n630), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n625), .B(KEYINPUT104), .Z(new_n646));
  AOI21_X1  g445(.A(new_n646), .B1(new_n637), .B2(new_n638), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n603), .B(G8gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n540), .ZN(new_n651));
  NAND2_X1  g450(.A1(G229gat), .A2(G233gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT13), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n541), .B2(new_n542), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n605), .A2(new_n540), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n656), .A2(KEYINPUT18), .A3(new_n652), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G113gat), .B(G141gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G169gat), .B(G197gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT12), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n655), .A2(new_n658), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n656), .A2(new_n652), .A3(new_n657), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(KEYINPUT90), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT90), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n666), .B2(new_n667), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n665), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n668), .A2(new_n655), .A3(new_n658), .ZN(new_n673));
  INV_X1    g472(.A(new_n664), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n649), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n618), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n275), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g481(.A(G8gat), .B1(new_n679), .B2(new_n400), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n679), .A2(new_n400), .A3(new_n685), .ZN(new_n686));
  MUX2_X1   g485(.A(new_n684), .B(KEYINPUT42), .S(new_n686), .Z(G1325gat));
  INV_X1    g486(.A(G15gat), .ZN(new_n688));
  INV_X1    g487(.A(new_n354), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n679), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n692));
  INV_X1    g491(.A(new_n469), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n679), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n470), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n567), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n459), .B2(new_n500), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n610), .A2(new_n616), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n701), .A2(new_n678), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n526), .A3(new_n275), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT45), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n706), .A2(new_n501), .A3(KEYINPUT44), .A4(new_n567), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT44), .B1(new_n701), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n678), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n275), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G29gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT108), .ZN(G1328gat));
  INV_X1    g514(.A(new_n400), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n703), .A2(new_n527), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT109), .Z(new_n719));
  NOR2_X1   g518(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT110), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n707), .A2(new_n708), .A3(new_n400), .A4(new_n710), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n719), .B(new_n721), .C1(new_n527), .C2(new_n722), .ZN(G1329gat));
  NAND3_X1  g522(.A1(new_n709), .A2(new_n469), .A3(new_n711), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT47), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n703), .A2(new_n728), .A3(new_n354), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n727), .B(new_n730), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n501), .A2(new_n706), .A3(new_n567), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n701), .A2(new_n706), .A3(KEYINPUT44), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n734), .A2(new_n470), .A3(new_n735), .A4(new_n711), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n703), .A2(new_n402), .A3(new_n470), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n739), .A2(KEYINPUT48), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n736), .A2(KEYINPUT112), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n736), .A2(KEYINPUT112), .ZN(new_n743));
  OAI21_X1  g542(.A(G50gat), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n738), .A2(KEYINPUT48), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n741), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n709), .A2(new_n748), .A3(new_n470), .A4(new_n711), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n736), .A2(KEYINPUT112), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n402), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(KEYINPUT113), .A3(new_n745), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n740), .B1(new_n747), .B2(new_n752), .ZN(G1331gat));
  INV_X1    g552(.A(new_n649), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n676), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n618), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n275), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n716), .ZN(new_n760));
  NOR2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n761), .B2(new_n760), .ZN(G1333gat));
  NAND3_X1  g563(.A1(new_n618), .A2(new_n354), .A3(new_n755), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT114), .ZN(new_n766));
  INV_X1    g565(.A(G71gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G71gat), .B1(new_n756), .B2(new_n693), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n470), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g575(.A1(new_n701), .A2(new_n677), .A3(new_n702), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n649), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n275), .A2(new_n510), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n610), .A2(new_n616), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n784), .A2(new_n676), .A3(new_n754), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n709), .A2(new_n275), .A3(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n782), .A2(new_n783), .B1(new_n510), .B2(new_n786), .ZN(G1336gat));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n400), .A2(G92gat), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n649), .B(new_n789), .C1(new_n779), .C2(new_n780), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n709), .A2(new_n716), .A3(new_n785), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n788), .B(new_n790), .C1(new_n791), .C2(new_n511), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g592(.A1(new_n709), .A2(new_n469), .A3(new_n785), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G99gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n689), .A2(G99gat), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n796), .A2(new_n797), .B1(new_n782), .B2(new_n798), .ZN(G1338gat));
  NOR3_X1   g598(.A1(new_n754), .A2(G106gat), .A3(new_n447), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT119), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n734), .A2(new_n785), .A3(new_n470), .A4(new_n735), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT118), .B1(new_n803), .B2(G106gat), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n803), .A2(new_n808), .ZN(new_n810));
  OAI21_X1  g609(.A(G106gat), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n812), .A3(new_n802), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n807), .A2(new_n813), .ZN(G1339gat));
  AND3_X1   g613(.A1(new_n631), .A2(new_n635), .A3(new_n643), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n637), .A2(new_n638), .A3(new_n646), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n639), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n647), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n642), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT55), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n639), .A2(new_n817), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n637), .A2(new_n638), .A3(new_n646), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  INV_X1    g624(.A(new_n642), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n647), .B2(new_n817), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n815), .B1(new_n821), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n676), .A2(new_n564), .A3(new_n566), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n651), .A2(new_n654), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n663), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n672), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n566), .B2(new_n564), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n829), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n700), .A2(new_n672), .A3(new_n649), .A4(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n702), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n649), .A2(new_n676), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n617), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n716), .A2(new_n456), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n454), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n676), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n649), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n784), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(G127gat), .ZN(G1342gat));
  INV_X1    g652(.A(new_n846), .ZN(new_n854));
  INV_X1    g653(.A(new_n454), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n700), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n857), .B(new_n858), .Z(G1343gat));
  NOR2_X1   g658(.A1(new_n447), .A2(new_n469), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(G141gat), .B1(new_n861), .B2(new_n676), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n784), .B1(new_n838), .B2(new_n839), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n784), .A2(new_n700), .A3(new_n842), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n470), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n716), .A2(new_n456), .A3(new_n469), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n869), .B(new_n870), .C1(KEYINPUT57), .C2(new_n866), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n676), .A2(G141gat), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n863), .B(KEYINPUT58), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n871), .A2(new_n872), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n862), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n205), .A3(new_n649), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n205), .A2(KEYINPUT59), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n871), .B2(new_n754), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT57), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n470), .B(new_n867), .C1(new_n864), .C2(new_n865), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n882), .A2(new_n649), .A3(new_n870), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT124), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI211_X1 g686(.A(KEYINPUT124), .B(new_n881), .C1(new_n884), .C2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(G1345gat));
  NOR3_X1   g688(.A1(new_n871), .A2(new_n207), .A3(new_n702), .ZN(new_n890));
  INV_X1    g689(.A(new_n861), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(new_n702), .ZN(new_n892));
  AOI21_X1  g691(.A(G155gat), .B1(new_n892), .B2(KEYINPUT125), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n891), .B2(new_n702), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n893), .B2(new_n895), .ZN(G1346gat));
  OAI21_X1  g695(.A(G162gat), .B1(new_n871), .B2(new_n700), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n861), .A2(new_n208), .A3(new_n567), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n400), .A2(new_n275), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n844), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(new_n855), .ZN(new_n902));
  AOI21_X1  g701(.A(G169gat), .B1(new_n902), .B2(new_n676), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n900), .B(KEYINPUT126), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n844), .A2(new_n855), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n677), .A2(new_n282), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n902), .A2(new_n283), .A3(new_n649), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n905), .A2(new_n649), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n283), .B2(new_n909), .ZN(G1349gat));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT60), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n784), .A2(new_n307), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n901), .A2(new_n855), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n311), .B1(new_n905), .B2(new_n784), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n912), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n905), .A2(new_n784), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G183gat), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n920), .A2(new_n911), .A3(KEYINPUT60), .A4(new_n915), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n918), .A2(new_n921), .ZN(G1350gat));
  AOI21_X1  g721(.A(new_n309), .B1(new_n905), .B2(new_n567), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n902), .A2(new_n309), .A3(new_n567), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n904), .A2(new_n693), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n883), .A3(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n357), .A3(new_n677), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n901), .A2(new_n860), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n676), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(new_n357), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n754), .A2(G204gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n901), .A2(new_n860), .A3(new_n935), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  NAND3_X1  g736(.A1(new_n882), .A2(new_n649), .A3(new_n883), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n938), .B2(new_n928), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1353gat));
  NAND3_X1  g739(.A1(new_n932), .A2(new_n368), .A3(new_n784), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n882), .A2(new_n784), .A3(new_n883), .A4(new_n929), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n369), .A3(new_n567), .ZN(new_n946));
  OAI21_X1  g745(.A(G218gat), .B1(new_n930), .B2(new_n700), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1355gat));
endmodule


