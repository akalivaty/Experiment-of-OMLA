//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT85), .A2(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT85), .A2(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT18), .A2(G131), .ZN(new_n196));
  NOR2_X1   g010(.A1(G237), .A2(G953), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n204), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(new_n206), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT87), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n195), .A2(new_n198), .ZN(new_n216));
  INV_X1    g030(.A(new_n196), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT86), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n219));
  AOI211_X1 g033(.A(new_n219), .B(new_n196), .C1(new_n195), .C2(new_n198), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n201), .B(new_n215), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n195), .A2(new_n198), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT89), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT89), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n225), .A3(G131), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n223), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G146), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n211), .B(KEYINPUT19), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n189), .B1(new_n221), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n215), .B1(new_n218), .B2(new_n220), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n199), .B(KEYINPUT88), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(new_n224), .B2(new_n226), .ZN(new_n241));
  INV_X1    g055(.A(new_n231), .ZN(new_n242));
  AOI21_X1  g056(.A(G146), .B1(new_n229), .B2(new_n230), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT90), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(new_n231), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n224), .A2(new_n240), .A3(new_n226), .A4(new_n227), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n239), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n236), .B1(new_n251), .B2(new_n189), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT20), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n225), .B1(new_n216), .B2(G131), .ZN(new_n256));
  AOI211_X1 g070(.A(KEYINPUT89), .B(new_n223), .C1(new_n195), .C2(new_n198), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT17), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(new_n258), .A3(new_n244), .A4(new_n247), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n189), .A3(new_n221), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n216), .A2(G131), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n256), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  OAI22_X1  g076(.A1(new_n262), .A2(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n263));
  INV_X1    g077(.A(new_n189), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT20), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n253), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  XNOR2_X1  g084(.A(G128), .B(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT13), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G128), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n272), .B(G134), .C1(KEYINPUT13), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n276));
  OR2_X1    g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n275), .B2(new_n276), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT92), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G122), .ZN(new_n283));
  INV_X1    g097(.A(G122), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT92), .A3(G116), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g102(.A1(KEYINPUT66), .A2(G116), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(G122), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT93), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G107), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n286), .B2(new_n290), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n290), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT93), .ZN(new_n298));
  AOI21_X1  g112(.A(G107), .B1(new_n298), .B2(new_n292), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n277), .B(new_n280), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT9), .B(G234), .ZN(new_n301));
  INV_X1    g115(.A(G217), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n301), .A2(new_n302), .A3(G953), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n290), .A2(KEYINPUT14), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n286), .B1(new_n290), .B2(KEYINPUT14), .ZN(new_n306));
  OAI21_X1  g120(.A(G107), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n271), .A2(new_n278), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n304), .B(new_n307), .C1(new_n279), .C2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n300), .A2(new_n303), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n303), .B1(new_n300), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n270), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT15), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G478), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT91), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n260), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n189), .B1(new_n259), .B2(new_n221), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n259), .A2(new_n221), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT91), .A3(new_n264), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n270), .ZN(new_n323));
  OAI21_X1  g137(.A(G475), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT95), .B(G952), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(G234), .A2(G237), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT21), .B(G898), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(G902), .A3(G953), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AND4_X1   g146(.A1(new_n269), .A2(new_n316), .A3(new_n324), .A4(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G214), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n288), .A2(G119), .A3(new_n289), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT67), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n288), .A2(new_n338), .A3(G119), .A4(new_n289), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n282), .A2(G119), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT2), .B(G113), .Z(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n337), .A2(new_n343), .A3(new_n339), .A4(new_n341), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(KEYINPUT68), .A3(new_n344), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n294), .A3(G104), .ZN(new_n352));
  INV_X1    g166(.A(G101), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n188), .A2(G107), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n350), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n353), .A2(KEYINPUT78), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n348), .A2(new_n349), .A3(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n337), .A2(KEYINPUT5), .A3(new_n339), .A4(new_n341), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n341), .A2(KEYINPUT5), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(G113), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n188), .B2(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n294), .A2(KEYINPUT79), .A3(G104), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n354), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G101), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(new_n355), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n347), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G122), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(new_n375), .A3(new_n373), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G143), .B(G146), .ZN(new_n380));
  AND2_X1   g194(.A1(KEYINPUT0), .A2(G128), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n273), .A2(G146), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT64), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(new_n207), .B2(G143), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n273), .A2(KEYINPUT64), .A3(G146), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT0), .A2(G128), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n382), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n207), .A2(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n273), .A2(G146), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT1), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .A4(G128), .ZN(new_n396));
  INV_X1    g210(.A(G128), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n393), .B2(KEYINPUT1), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n205), .B(new_n396), .C1(new_n387), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n400), .A3(G125), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n374), .A2(new_n406), .A3(new_n376), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n379), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n375), .B(KEYINPUT83), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT8), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n372), .A2(new_n347), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n364), .A2(KEYINPUT84), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n365), .A2(G113), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n364), .B2(KEYINPUT84), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n372), .B1(new_n366), .B2(new_n347), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT7), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n404), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n392), .A2(new_n399), .A3(new_n401), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n391), .A2(new_n399), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n418), .B2(new_n404), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n423), .A3(new_n378), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(new_n270), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n408), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G210), .B1(G237), .B2(G902), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n408), .A2(new_n425), .A3(new_n427), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n335), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  INV_X1    g248(.A(G227), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(G953), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n434), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT11), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n278), .B2(G137), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n278), .A2(G137), .ZN(new_n441));
  INV_X1    g255(.A(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(KEYINPUT11), .A3(G134), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G131), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n440), .A2(new_n443), .A3(new_n223), .A4(new_n441), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n371), .A2(new_n355), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n395), .A2(new_n393), .A3(new_n394), .A4(G128), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G128), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n393), .A2(new_n394), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT80), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n448), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n396), .B1(new_n387), .B2(new_n398), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n355), .B2(new_n371), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n447), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n454), .B1(new_n398), .B2(new_n380), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n396), .A3(new_n456), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n372), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n273), .A2(KEYINPUT64), .A3(G146), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT64), .B1(new_n273), .B2(G146), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n393), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n449), .B1(new_n468), .B2(new_n451), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n448), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT12), .A3(new_n447), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT10), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n447), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n381), .A2(new_n388), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n468), .A2(new_n477), .B1(new_n380), .B2(new_n381), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n355), .A2(KEYINPUT4), .B1(new_n357), .B2(new_n358), .ZN(new_n479));
  INV_X1    g293(.A(new_n361), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n372), .A2(KEYINPUT10), .A3(new_n458), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n475), .A2(new_n476), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n438), .B1(new_n473), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT12), .B1(new_n471), .B2(new_n447), .ZN(new_n485));
  AOI211_X1 g299(.A(new_n461), .B(new_n476), .C1(new_n465), .C2(new_n470), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n438), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n437), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT10), .B1(new_n372), .B2(new_n464), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n469), .A2(new_n448), .A3(new_n474), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n390), .B1(new_n360), .B2(new_n361), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n437), .B1(new_n493), .B2(new_n476), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n481), .B(new_n482), .C1(new_n457), .C2(KEYINPUT10), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n447), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(G469), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n270), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n483), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n437), .ZN(new_n502));
  INV_X1    g316(.A(new_n437), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n483), .C1(new_n485), .C2(new_n486), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n505), .B2(new_n499), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n433), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n333), .A2(new_n431), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n302), .B1(G234), .B2(new_n270), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT24), .B(G110), .Z(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  INV_X1    g326(.A(G119), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(G128), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n397), .A2(G119), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n397), .A2(G119), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT74), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n511), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n397), .A2(KEYINPUT23), .A3(G119), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n521), .C1(new_n514), .C2(KEYINPUT23), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G110), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n231), .B(new_n213), .C1(new_n520), .C2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n516), .A2(new_n519), .A3(new_n511), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(G110), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(new_n242), .C2(new_n243), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT22), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(G137), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n524), .B(new_n534), .C1(new_n529), .C2(new_n530), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n270), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT25), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT25), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(KEYINPUT76), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n510), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n509), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n537), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT77), .Z(new_n546));
  NOR2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n348), .A2(new_n349), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n478), .A2(new_n447), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT65), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n278), .B2(G137), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n442), .A2(KEYINPUT65), .A3(G134), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n441), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G131), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n458), .A2(new_n446), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT30), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT69), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n549), .A2(new_n555), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n548), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n197), .A2(G210), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT27), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT26), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G101), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT26), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n566), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n353), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n556), .B1(new_n349), .B2(new_n348), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n563), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n573), .A2(KEYINPUT28), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n554), .A2(new_n446), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n576), .A2(new_n458), .B1(new_n478), .B2(new_n447), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n347), .A2(new_n346), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n340), .B1(new_n336), .B2(KEYINPUT67), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n343), .B1(new_n579), .B2(new_n339), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n349), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n556), .A2(new_n348), .A3(new_n349), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT28), .B1(new_n585), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n575), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n574), .B1(new_n588), .B2(new_n572), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n270), .B1(new_n589), .B2(KEYINPUT29), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(KEYINPUT72), .A3(new_n585), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT72), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n548), .A2(new_n592), .A3(new_n577), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(KEYINPUT28), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n568), .A2(new_n571), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT29), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n575), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT73), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n594), .A2(KEYINPUT73), .A3(new_n575), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n590), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(G472), .A2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT71), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n581), .A2(new_n582), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT69), .B(new_n559), .C1(new_n549), .C2(new_n555), .ZN(new_n608));
  AND4_X1   g422(.A1(new_n549), .A2(new_n555), .A3(new_n560), .A4(new_n561), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n572), .A3(new_n583), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT31), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n558), .A2(new_n562), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n573), .B1(new_n613), .B2(new_n607), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT31), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(new_n615), .A3(new_n572), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n607), .A2(KEYINPUT70), .A3(new_n556), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(KEYINPUT28), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n572), .B1(new_n620), .B2(new_n575), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n606), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n588), .A2(new_n595), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT71), .A3(new_n612), .A4(new_n616), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n605), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n603), .B1(new_n625), .B2(KEYINPUT32), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT32), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n627), .B(new_n605), .C1(new_n622), .C2(new_n624), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n508), .B(new_n547), .C1(new_n626), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  AOI21_X1  g444(.A(new_n615), .B1(new_n614), .B2(new_n572), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n563), .A2(new_n595), .A3(KEYINPUT31), .A4(new_n573), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT71), .B1(new_n633), .B2(new_n623), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n617), .A2(new_n621), .A3(new_n606), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n270), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n604), .B1(new_n634), .B2(new_n635), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n547), .ZN(new_n640));
  INV_X1    g454(.A(new_n507), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n267), .B1(new_n266), .B2(new_n253), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT20), .B(new_n254), .C1(new_n260), .C2(new_n265), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G475), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n321), .A2(new_n264), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n317), .A3(new_n260), .ZN(new_n648));
  AOI21_X1  g462(.A(G902), .B1(new_n319), .B2(KEYINPUT91), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(new_n311), .B2(new_n312), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n300), .A2(new_n309), .ZN(new_n654));
  INV_X1    g468(.A(new_n303), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n656), .A2(KEYINPUT33), .A3(new_n310), .ZN(new_n657));
  INV_X1    g471(.A(G478), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n313), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n431), .A3(new_n332), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n642), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  NAND3_X1  g483(.A1(new_n255), .A2(KEYINPUT96), .A3(new_n268), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT96), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(new_n643), .B2(new_n644), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n316), .A2(new_n650), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n332), .A2(new_n431), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n642), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  AND3_X1   g492(.A1(new_n538), .A2(KEYINPUT76), .A3(new_n541), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n541), .B1(new_n538), .B2(KEYINPUT76), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n509), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n531), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n531), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n544), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT97), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n531), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(KEYINPUT97), .A3(new_n544), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n681), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n333), .A2(new_n431), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n638), .A3(new_n507), .A4(new_n637), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  NAND2_X1  g510(.A1(new_n638), .A2(new_n627), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n625), .A2(KEYINPUT32), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n603), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n431), .A2(new_n507), .A3(new_n692), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n328), .B1(G900), .B2(new_n331), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n674), .A2(new_n673), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n699), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  INV_X1    g518(.A(new_n430), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n427), .B1(new_n408), .B2(new_n425), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n705), .A2(KEYINPUT98), .A3(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT98), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n429), .B2(new_n430), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT38), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT38), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n707), .B2(new_n709), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n701), .B(KEYINPUT39), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n507), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT40), .Z(new_n717));
  INV_X1    g531(.A(new_n614), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n572), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n270), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n572), .B1(new_n591), .B2(new_n593), .ZN(new_n721));
  OAI21_X1  g535(.A(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n697), .A2(new_n698), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n269), .A2(new_n324), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n313), .A2(new_n314), .A3(G478), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n270), .B(new_n315), .C1(new_n311), .C2(new_n312), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n728), .A2(new_n692), .A3(new_n335), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n714), .A2(new_n717), .A3(new_n723), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n273), .ZN(G45));
  OAI211_X1 g545(.A(new_n662), .B(new_n701), .C1(new_n645), .C2(new_n650), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n699), .A2(new_n700), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  AOI21_X1  g549(.A(new_n595), .B1(new_n620), .B2(new_n575), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n596), .B1(new_n736), .B2(new_n574), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n270), .A3(new_n600), .A4(new_n601), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n638), .A2(new_n627), .B1(G472), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n640), .B1(new_n739), .B2(new_n698), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n437), .A2(new_n501), .B1(new_n494), .B2(new_n473), .ZN(new_n741));
  OAI21_X1  g555(.A(G469), .B1(new_n741), .B2(G902), .ZN(new_n742));
  INV_X1    g556(.A(new_n504), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n503), .B1(new_n496), .B2(new_n483), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n499), .B(new_n270), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n432), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT99), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT99), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n742), .A2(new_n748), .A3(new_n432), .A4(new_n745), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n747), .A2(KEYINPUT100), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT100), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n740), .A2(new_n666), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n699), .A3(new_n547), .A4(new_n675), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT101), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n740), .A2(KEYINPUT101), .A3(new_n675), .A4(new_n752), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  AND3_X1   g575(.A1(new_n431), .A2(new_n747), .A3(new_n749), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n651), .A2(new_n332), .A3(new_n316), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n687), .A2(new_n690), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n543), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n762), .B(new_n766), .C1(new_n626), .C2(new_n628), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(KEYINPUT102), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n572), .B1(new_n594), .B2(new_n575), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n631), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n616), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n770), .A2(new_n631), .A3(new_n769), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n604), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(G472), .ZN(new_n775));
  AOI21_X1  g589(.A(G902), .B1(new_n622), .B2(new_n624), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n774), .B(new_n547), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n724), .A2(new_n431), .A3(new_n332), .A4(new_n727), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n752), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  INV_X1    g595(.A(new_n773), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n616), .A3(new_n771), .ZN(new_n783));
  AOI22_X1  g597(.A1(new_n636), .A2(G472), .B1(new_n783), .B2(new_n604), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n732), .A2(KEYINPUT103), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT103), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n724), .A2(new_n786), .A3(new_n662), .A4(new_n701), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n784), .A2(new_n788), .A3(new_n762), .A4(new_n692), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n626), .B1(new_n791), .B2(new_n698), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n628), .A2(KEYINPUT105), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n640), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n498), .A2(KEYINPUT104), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT104), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n489), .A2(new_n796), .A3(G469), .A4(new_n497), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n506), .A3(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n705), .A2(new_n335), .A3(new_n706), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n432), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(KEYINPUT42), .A3(new_n788), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT42), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n699), .A2(new_n800), .A3(new_n547), .A4(new_n788), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n794), .A2(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(new_n223), .ZN(G33));
  AND4_X1   g619(.A1(new_n699), .A2(new_n800), .A3(new_n547), .A4(new_n702), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n278), .ZN(G36));
  OAI21_X1  g621(.A(KEYINPUT43), .B1(new_n724), .B2(new_n663), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n724), .A2(new_n663), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT43), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n639), .A2(new_n692), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT44), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT107), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n799), .B(KEYINPUT108), .Z(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n812), .B2(KEYINPUT44), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n485), .A2(new_n486), .ZN(new_n819));
  INV_X1    g633(.A(new_n483), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT81), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n503), .B1(new_n821), .B2(new_n487), .ZN(new_n822));
  INV_X1    g636(.A(new_n497), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n497), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(G469), .ZN(new_n826));
  INV_X1    g640(.A(new_n500), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT46), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT106), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(KEYINPUT46), .A3(new_n827), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n745), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(KEYINPUT106), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n432), .B(new_n715), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  OAI21_X1  g650(.A(new_n432), .B1(new_n831), .B2(new_n832), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT47), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n432), .C1(new_n831), .C2(new_n832), .ZN(new_n840));
  INV_X1    g654(.A(new_n799), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n699), .A2(new_n547), .A3(new_n732), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(G140), .ZN(G42));
  OR2_X1    g658(.A1(G952), .A2(G953), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n799), .A2(new_n749), .A3(new_n747), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n723), .A2(new_n640), .A3(new_n846), .A4(new_n328), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n664), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n326), .ZN(new_n849));
  INV_X1    g663(.A(new_n328), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n811), .A2(new_n850), .A3(new_n808), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n777), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n762), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT117), .Z(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n846), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n794), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n849), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n852), .A2(new_n815), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n838), .A2(new_n840), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n742), .A2(new_n433), .A3(new_n745), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n747), .A2(new_n335), .A3(new_n749), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n711), .B2(new_n713), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n866), .B1(new_n868), .B2(new_n852), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT50), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n724), .A2(new_n662), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n784), .A2(new_n692), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n847), .A2(new_n872), .B1(new_n874), .B2(new_n855), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n870), .A2(new_n871), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n860), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n871), .A3(new_n875), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n864), .A2(new_n878), .A3(KEYINPUT51), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n859), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT118), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n859), .B(new_n882), .C1(new_n877), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n794), .A2(new_n801), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n803), .A2(new_n802), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n841), .A2(new_n765), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n784), .A2(new_n788), .A3(new_n432), .A4(new_n798), .ZN(new_n892));
  INV_X1    g706(.A(new_n701), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n727), .A2(new_n650), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n507), .A2(new_n673), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n626), .B2(new_n628), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n891), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(new_n806), .A3(KEYINPUT112), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT112), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n895), .B1(new_n739), .B2(new_n698), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n798), .A2(new_n785), .A3(new_n787), .A4(new_n432), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n890), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n740), .A2(new_n702), .A3(new_n800), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n889), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n780), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n629), .A2(new_n694), .A3(new_n767), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n665), .A2(KEYINPUT110), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n724), .A2(KEYINPUT111), .A3(new_n316), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT111), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n651), .B2(new_n727), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n332), .B(new_n431), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT110), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n664), .A2(new_n431), .A3(new_n917), .A4(new_n332), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n912), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n642), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n760), .A2(new_n911), .A3(new_n753), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n908), .A2(new_n921), .ZN(new_n922));
  OAI221_X1 g736(.A(new_n700), .B1(new_n702), .B2(new_n733), .C1(new_n626), .C2(new_n628), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n543), .A2(new_n764), .A3(new_n893), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n798), .A2(new_n924), .A3(new_n432), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n431), .A2(new_n724), .A3(new_n727), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n723), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n927), .A3(new_n789), .ZN(new_n928));
  XOR2_X1   g742(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT115), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n923), .A2(new_n927), .A3(KEYINPUT52), .A4(new_n789), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(KEYINPUT113), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(KEYINPUT113), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n931), .B(new_n933), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n886), .B1(new_n922), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n760), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n629), .A2(new_n767), .A3(new_n694), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(new_n753), .A3(new_n780), .A4(new_n920), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT112), .B1(new_n898), .B2(new_n806), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n905), .A2(new_n906), .A3(new_n900), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n804), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT52), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n928), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n934), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n886), .A2(new_n942), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n885), .B1(new_n938), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n942), .A2(new_n945), .A3(new_n948), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT53), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n922), .A2(new_n937), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n952), .B(KEYINPUT54), .C1(new_n953), .C2(KEYINPUT53), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n845), .B1(new_n884), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n640), .A2(new_n335), .A3(new_n433), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n742), .A2(new_n745), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT49), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n809), .A3(new_n959), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n714), .A2(new_n960), .A3(new_n723), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT109), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n956), .A2(new_n962), .ZN(G75));
  NAND2_X1  g777(.A1(new_n931), .A2(new_n933), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT113), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n934), .B(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n943), .A2(new_n944), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n431), .A2(new_n747), .A3(new_n749), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n969), .A2(new_n763), .A3(new_n765), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n776), .A2(new_n775), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n971), .A2(new_n625), .A3(new_n641), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n970), .A2(new_n699), .B1(new_n972), .B2(new_n693), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n753), .A3(new_n780), .A4(new_n629), .ZN(new_n974));
  INV_X1    g788(.A(new_n920), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n968), .A2(new_n976), .A3(new_n760), .A4(new_n889), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT53), .B1(new_n967), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n922), .A2(new_n886), .A3(new_n948), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n978), .A2(new_n979), .A3(G210), .A4(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n405), .B(KEYINPUT55), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT120), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n379), .A2(new_n407), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT119), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n982), .B(new_n984), .Z(new_n985));
  XOR2_X1   g799(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n986));
  AND3_X1   g800(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT56), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n191), .A2(G952), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(G51));
  XNOR2_X1  g805(.A(new_n500), .B(KEYINPUT57), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n938), .A2(new_n949), .A3(new_n885), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT54), .B1(new_n978), .B2(new_n979), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n741), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n978), .A2(new_n979), .ZN(new_n998));
  OR3_X1    g812(.A1(new_n998), .A2(new_n270), .A3(new_n826), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(G54));
  INV_X1    g814(.A(new_n990), .ZN(new_n1001));
  NAND2_X1  g815(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT122), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n978), .A2(new_n979), .A3(G902), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1001), .B1(new_n1004), .B2(new_n252), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n252), .B2(new_n1004), .ZN(G60));
  NOR2_X1   g820(.A1(new_n993), .A2(new_n994), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n653), .A2(new_n657), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G478), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT59), .Z(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1001), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n955), .B2(new_n1011), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(new_n1014), .ZN(G63));
  NAND2_X1  g829(.A1(G217), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT60), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n978), .A2(new_n979), .A3(new_n689), .A4(new_n1018), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n938), .A2(new_n949), .A3(new_n1017), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n536), .A2(new_n537), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1001), .B(new_n1019), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g837(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1021), .B1(new_n998), .B2(new_n1017), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1027), .A2(new_n1001), .A3(new_n1024), .A4(new_n1019), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1026), .A2(new_n1028), .ZN(G66));
  OAI21_X1  g843(.A(G953), .B1(new_n329), .B2(new_n403), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT124), .Z(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n942), .B2(G953), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT125), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n984), .B1(G898), .B2(new_n191), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1033), .B(new_n1034), .Z(G69));
  AND2_X1   g849(.A1(new_n794), .A2(new_n926), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n834), .B1(new_n817), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n923), .A2(new_n789), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n804), .A2(new_n806), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1037), .A2(new_n843), .A3(new_n1039), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n1040), .A2(G953), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n613), .B(KEYINPUT126), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(new_n232), .Z(new_n1043));
  NAND3_X1  g857(.A1(new_n435), .A2(KEYINPUT127), .A3(G900), .ZN(new_n1044));
  OAI21_X1  g858(.A(G953), .B1(KEYINPUT127), .B2(G900), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1043), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1048));
  NOR3_X1   g862(.A1(new_n913), .A2(new_n915), .A3(new_n664), .ZN(new_n1049));
  NOR3_X1   g863(.A1(new_n1049), .A2(new_n716), .A3(new_n841), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n740), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n835), .A2(new_n191), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g866(.A1(new_n730), .A2(new_n1038), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1054), .A2(new_n843), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1048), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g871(.A1(new_n1041), .A2(new_n1047), .B1(new_n1043), .B2(new_n1057), .ZN(G72));
  NAND2_X1  g872(.A1(G472), .A2(G902), .ZN(new_n1059));
  XOR2_X1   g873(.A(new_n1059), .B(KEYINPUT63), .Z(new_n1060));
  OAI21_X1  g874(.A(new_n1060), .B1(new_n1040), .B2(new_n921), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n574), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n835), .A2(new_n942), .A3(new_n1051), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1060), .B1(new_n1063), .B2(new_n1056), .ZN(new_n1064));
  INV_X1    g878(.A(new_n719), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n990), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(new_n574), .ZN(new_n1067));
  AND3_X1   g881(.A1(new_n719), .A2(new_n1067), .A3(new_n1060), .ZN(new_n1068));
  OAI211_X1 g882(.A(new_n952), .B(new_n1068), .C1(new_n953), .C2(KEYINPUT53), .ZN(new_n1069));
  AND3_X1   g883(.A1(new_n1062), .A2(new_n1066), .A3(new_n1069), .ZN(G57));
endmodule


