

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755;

  AND2_X1 U369 ( .A1(n425), .A2(n456), .ZN(n721) );
  AND2_X1 U370 ( .A1(n707), .A2(n596), .ZN(n598) );
  AND2_X1 U371 ( .A1(n376), .A2(n573), .ZN(n596) );
  XNOR2_X1 U372 ( .A(n512), .B(n511), .ZN(n547) );
  XNOR2_X1 U373 ( .A(G131), .B(G143), .ZN(n475) );
  NOR2_X1 U374 ( .A1(G953), .A2(G237), .ZN(n504) );
  XNOR2_X2 U375 ( .A(n494), .B(n493), .ZN(n509) );
  XNOR2_X2 U376 ( .A(n574), .B(KEYINPUT78), .ZN(n605) );
  AND2_X1 U377 ( .A1(n368), .A2(n370), .ZN(n367) );
  XNOR2_X1 U378 ( .A(n598), .B(n597), .ZN(n753) );
  BUF_X2 U379 ( .A(n547), .Z(n696) );
  INV_X2 U380 ( .A(G125), .ZN(n384) );
  NOR2_X2 U381 ( .A1(n686), .A2(n685), .ZN(n422) );
  XNOR2_X2 U382 ( .A(n470), .B(KEYINPUT4), .ZN(n494) );
  NOR2_X1 U383 ( .A1(n413), .A2(n584), .ZN(n668) );
  XNOR2_X1 U384 ( .A(n442), .B(G953), .ZN(n745) );
  AND2_X1 U385 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U386 ( .A(n668), .B(n412), .ZN(n411) );
  XNOR2_X1 U387 ( .A(n583), .B(KEYINPUT112), .ZN(n413) );
  AND2_X1 U388 ( .A1(n403), .A2(n669), .ZN(n398) );
  AND2_X1 U389 ( .A1(n581), .A2(n580), .ZN(n599) );
  AND2_X1 U390 ( .A1(n573), .A2(n405), .ZN(n530) );
  INV_X1 U391 ( .A(n549), .ZN(n346) );
  INV_X1 U392 ( .A(n564), .ZN(n572) );
  XNOR2_X1 U393 ( .A(n444), .B(n443), .ZN(n508) );
  XNOR2_X1 U394 ( .A(KEYINPUT69), .B(G101), .ZN(n507) );
  XOR2_X1 U395 ( .A(G137), .B(G146), .Z(n506) );
  BUF_X1 U396 ( .A(n590), .Z(n347) );
  BUF_X1 U397 ( .A(n656), .Z(n348) );
  NOR2_X2 U398 ( .A1(n438), .A2(n431), .ZN(n727) );
  XNOR2_X1 U399 ( .A(n547), .B(KEYINPUT108), .ZN(n577) );
  BUF_X1 U400 ( .A(n582), .Z(n618) );
  XNOR2_X1 U401 ( .A(n569), .B(KEYINPUT81), .ZN(n576) );
  OR2_X1 U402 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U403 ( .A(G119), .B(KEYINPUT3), .ZN(n443) );
  XOR2_X1 U404 ( .A(G113), .B(G116), .Z(n444) );
  XNOR2_X1 U405 ( .A(n495), .B(G137), .ZN(n515) );
  INV_X1 U406 ( .A(G140), .ZN(n495) );
  XNOR2_X1 U407 ( .A(G134), .B(G131), .ZN(n493) );
  XNOR2_X1 U408 ( .A(n391), .B(KEYINPUT105), .ZN(n685) );
  XNOR2_X1 U409 ( .A(n526), .B(n525), .ZN(n564) );
  NOR2_X1 U410 ( .A1(n383), .A2(n415), .ZN(n382) );
  INV_X1 U411 ( .A(KEYINPUT107), .ZN(n409) );
  XNOR2_X1 U412 ( .A(n441), .B(n352), .ZN(n387) );
  XNOR2_X1 U413 ( .A(n474), .B(KEYINPUT18), .ZN(n441) );
  XNOR2_X1 U414 ( .A(n454), .B(n453), .ZN(n582) );
  XNOR2_X1 U415 ( .A(n452), .B(n451), .ZN(n453) );
  INV_X1 U416 ( .A(KEYINPUT80), .ZN(n451) );
  INV_X1 U417 ( .A(n576), .ZN(n423) );
  NAND2_X1 U418 ( .A1(n572), .A2(n571), .ZN(n586) );
  NOR2_X1 U419 ( .A1(n576), .A2(n570), .ZN(n571) );
  OR2_X1 U420 ( .A1(n652), .A2(G902), .ZN(n503) );
  XNOR2_X1 U421 ( .A(n509), .B(n373), .ZN(n637) );
  XNOR2_X1 U422 ( .A(n372), .B(n508), .ZN(n373) );
  XNOR2_X1 U423 ( .A(n375), .B(n374), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n506), .B(n505), .ZN(n374) );
  XNOR2_X1 U425 ( .A(n407), .B(n406), .ZN(n731) );
  XNOR2_X1 U426 ( .A(G104), .B(G107), .ZN(n406) );
  XNOR2_X1 U427 ( .A(n408), .B(G110), .ZN(n407) );
  INV_X1 U428 ( .A(KEYINPUT92), .ZN(n408) );
  XNOR2_X1 U429 ( .A(n445), .B(G122), .ZN(n446) );
  XOR2_X1 U430 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n445) );
  INV_X1 U431 ( .A(G128), .ZN(n447) );
  XNOR2_X1 U432 ( .A(n731), .B(n507), .ZN(n498) );
  OR2_X1 U433 ( .A1(n599), .A2(n404), .ZN(n403) );
  NOR2_X1 U434 ( .A1(n401), .A2(n350), .ZN(n400) );
  AND2_X1 U435 ( .A1(n599), .A2(n402), .ZN(n401) );
  XNOR2_X1 U436 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n491) );
  INV_X1 U437 ( .A(KEYINPUT64), .ZN(n442) );
  XNOR2_X1 U438 ( .A(n520), .B(n416), .ZN(n729) );
  XNOR2_X1 U439 ( .A(n518), .B(n417), .ZN(n416) );
  XNOR2_X1 U440 ( .A(n419), .B(n418), .ZN(n417) );
  INV_X1 U441 ( .A(KEYINPUT86), .ZN(n412) );
  NAND2_X1 U442 ( .A1(n353), .A2(n575), .ZN(n380) );
  NAND2_X1 U443 ( .A1(n575), .A2(n360), .ZN(n381) );
  NOR2_X1 U444 ( .A1(n565), .A2(n745), .ZN(n395) );
  INV_X1 U445 ( .A(G237), .ZN(n450) );
  INV_X1 U446 ( .A(G902), .ZN(n510) );
  XNOR2_X1 U447 ( .A(n507), .B(KEYINPUT5), .ZN(n375) );
  XOR2_X1 U448 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n480) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  XNOR2_X1 U450 ( .A(n396), .B(n356), .ZN(n458) );
  XNOR2_X1 U451 ( .A(KEYINPUT75), .B(KEYINPUT14), .ZN(n396) );
  INV_X1 U452 ( .A(n601), .ZN(n404) );
  XNOR2_X1 U453 ( .A(n515), .B(n516), .ZN(n418) );
  XNOR2_X1 U454 ( .A(n517), .B(n514), .ZN(n419) );
  XNOR2_X1 U455 ( .A(G116), .B(G122), .ZN(n463) );
  XOR2_X1 U456 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n464) );
  XNOR2_X1 U457 ( .A(G134), .B(G107), .ZN(n462) );
  XNOR2_X1 U458 ( .A(n509), .B(n515), .ZN(n744) );
  XNOR2_X1 U459 ( .A(n386), .B(n498), .ZN(n449) );
  XNOR2_X1 U460 ( .A(n387), .B(n440), .ZN(n386) );
  XNOR2_X1 U461 ( .A(n536), .B(KEYINPUT33), .ZN(n716) );
  NAND2_X1 U462 ( .A1(n582), .A2(n683), .ZN(n590) );
  AND2_X1 U463 ( .A1(n530), .A2(n423), .ZN(n581) );
  XNOR2_X1 U464 ( .A(n377), .B(KEYINPUT28), .ZN(n376) );
  NOR2_X1 U465 ( .A1(n577), .A2(n586), .ZN(n377) );
  XNOR2_X1 U466 ( .A(n590), .B(KEYINPUT19), .ZN(n385) );
  INV_X1 U467 ( .A(n699), .ZN(n405) );
  NAND2_X1 U468 ( .A1(n700), .A2(n346), .ZN(n430) );
  XNOR2_X1 U469 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U470 ( .A(n644), .B(n643), .ZN(n645) );
  AND2_X1 U471 ( .A1(n726), .A2(G210), .ZN(n437) );
  AND2_X1 U472 ( .A1(n433), .A2(n647), .ZN(n432) );
  NAND2_X1 U473 ( .A1(n435), .A2(n434), .ZN(n433) );
  INV_X1 U474 ( .A(G210), .ZN(n434) );
  INV_X1 U475 ( .A(n681), .ZN(n427) );
  XNOR2_X1 U476 ( .A(n388), .B(KEYINPUT82), .ZN(n362) );
  XNOR2_X1 U477 ( .A(n728), .B(n729), .ZN(n394) );
  AND2_X1 U478 ( .A1(n622), .A2(KEYINPUT2), .ZN(n349) );
  AND2_X1 U479 ( .A1(n399), .A2(n601), .ZN(n350) );
  XOR2_X1 U480 ( .A(G113), .B(G122), .Z(n351) );
  NAND2_X1 U481 ( .A1(n429), .A2(n700), .ZN(n546) );
  XNOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT17), .ZN(n352) );
  AND2_X1 U483 ( .A1(n605), .A2(n415), .ZN(n353) );
  AND2_X1 U484 ( .A1(n692), .A2(KEYINPUT107), .ZN(n354) );
  AND2_X1 U485 ( .A1(n575), .A2(n382), .ZN(n355) );
  AND2_X1 U486 ( .A1(G234), .A2(G237), .ZN(n356) );
  AND2_X1 U487 ( .A1(n534), .A2(n409), .ZN(n357) );
  AND2_X1 U488 ( .A1(n378), .A2(n381), .ZN(n358) );
  XNOR2_X1 U489 ( .A(n449), .B(n448), .ZN(n723) );
  XOR2_X1 U490 ( .A(n461), .B(KEYINPUT68), .Z(n359) );
  AND2_X1 U491 ( .A1(n383), .A2(n415), .ZN(n360) );
  OR2_X1 U492 ( .A1(n745), .A2(G952), .ZN(n647) );
  INV_X1 U493 ( .A(KEYINPUT47), .ZN(n383) );
  NAND2_X1 U494 ( .A1(n361), .A2(n720), .ZN(n426) );
  NAND2_X1 U495 ( .A1(n362), .A2(n427), .ZN(n361) );
  XNOR2_X1 U496 ( .A(n563), .B(n562), .ZN(n363) );
  XNOR2_X1 U497 ( .A(n563), .B(n562), .ZN(n738) );
  XNOR2_X2 U498 ( .A(n628), .B(KEYINPUT65), .ZN(n364) );
  NAND2_X2 U499 ( .A1(n627), .A2(n365), .ZN(n628) );
  XNOR2_X2 U500 ( .A(n573), .B(KEYINPUT1), .ZN(n592) );
  NAND2_X1 U501 ( .A1(n385), .A2(n439), .ZN(n428) );
  XNOR2_X1 U502 ( .A(n426), .B(KEYINPUT125), .ZN(n425) );
  NAND2_X1 U503 ( .A1(n410), .A2(n623), .ZN(n365) );
  NAND2_X1 U504 ( .A1(n410), .A2(n623), .ZN(n388) );
  NAND2_X1 U505 ( .A1(n367), .A2(n366), .ZN(n389) );
  NAND2_X1 U506 ( .A1(n656), .A2(n357), .ZN(n366) );
  NAND2_X1 U507 ( .A1(n369), .A2(n692), .ZN(n656) );
  NAND2_X1 U508 ( .A1(n369), .A2(n354), .ZN(n368) );
  XNOR2_X1 U509 ( .A(n513), .B(KEYINPUT88), .ZN(n369) );
  NAND2_X1 U510 ( .A1(n371), .A2(KEYINPUT107), .ZN(n370) );
  INV_X1 U511 ( .A(n534), .ZN(n371) );
  XNOR2_X2 U512 ( .A(n424), .B(n447), .ZN(n470) );
  NAND2_X1 U513 ( .A1(n379), .A2(n355), .ZN(n378) );
  INV_X1 U514 ( .A(n605), .ZN(n379) );
  NAND2_X1 U515 ( .A1(n358), .A2(n380), .ZN(n414) );
  XNOR2_X2 U516 ( .A(n384), .B(G146), .ZN(n474) );
  AND2_X1 U517 ( .A1(n385), .A2(n596), .ZN(n574) );
  NAND2_X1 U518 ( .A1(n389), .A2(n544), .ZN(n545) );
  NOR2_X2 U519 ( .A1(n681), .A2(n625), .ZN(n627) );
  XNOR2_X1 U520 ( .A(n390), .B(n484), .ZN(n485) );
  NOR2_X1 U521 ( .A1(n644), .A2(G902), .ZN(n390) );
  NOR2_X1 U522 ( .A1(n540), .A2(n539), .ZN(n391) );
  XNOR2_X1 U523 ( .A(n478), .B(n392), .ZN(n482) );
  XNOR2_X1 U524 ( .A(n477), .B(n351), .ZN(n392) );
  NAND2_X1 U525 ( .A1(n752), .A2(KEYINPUT44), .ZN(n544) );
  XNOR2_X2 U526 ( .A(n543), .B(KEYINPUT35), .ZN(n752) );
  AND2_X1 U527 ( .A1(n535), .A2(n592), .ZN(n536) );
  XNOR2_X1 U528 ( .A(n393), .B(KEYINPUT99), .ZN(n531) );
  NAND2_X1 U529 ( .A1(n529), .A2(n530), .ZN(n393) );
  NAND2_X1 U530 ( .A1(n658), .A2(n673), .ZN(n533) );
  NAND2_X1 U531 ( .A1(n397), .A2(n622), .ZN(n420) );
  NOR2_X1 U532 ( .A1(n394), .A2(n730), .ZN(G66) );
  XNOR2_X1 U533 ( .A(n395), .B(KEYINPUT109), .ZN(n566) );
  NAND2_X1 U534 ( .A1(n397), .A2(n349), .ZN(n624) );
  XNOR2_X2 U535 ( .A(n613), .B(n612), .ZN(n397) );
  NAND2_X1 U536 ( .A1(n400), .A2(n403), .ZN(n621) );
  NAND2_X1 U537 ( .A1(n400), .A2(n398), .ZN(n603) );
  INV_X1 U538 ( .A(n682), .ZN(n399) );
  AND2_X1 U539 ( .A1(n682), .A2(n404), .ZN(n402) );
  XNOR2_X2 U540 ( .A(n503), .B(n502), .ZN(n573) );
  INV_X1 U541 ( .A(n626), .ZN(n410) );
  NAND2_X1 U542 ( .A1(n414), .A2(n411), .ZN(n585) );
  INV_X1 U543 ( .A(KEYINPUT85), .ZN(n415) );
  NOR2_X1 U544 ( .A1(n738), .A2(n420), .ZN(n626) );
  XNOR2_X1 U545 ( .A(n420), .B(n747), .ZN(n746) );
  XNOR2_X1 U546 ( .A(n422), .B(n421), .ZN(n707) );
  INV_X1 U547 ( .A(KEYINPUT41), .ZN(n421) );
  NAND2_X1 U548 ( .A1(n682), .A2(n683), .ZN(n686) );
  XNOR2_X2 U549 ( .A(n618), .B(n595), .ZN(n682) );
  XNOR2_X2 U550 ( .A(KEYINPUT79), .B(G143), .ZN(n424) );
  XNOR2_X2 U551 ( .A(n428), .B(n359), .ZN(n537) );
  INV_X1 U552 ( .A(n552), .ZN(n429) );
  NOR2_X1 U553 ( .A1(n552), .A2(n430), .ZN(n513) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n552) );
  NAND2_X1 U555 ( .A1(n364), .A2(n437), .ZN(n436) );
  XNOR2_X2 U556 ( .A(n628), .B(KEYINPUT65), .ZN(n722) );
  NAND2_X1 U557 ( .A1(n436), .A2(n432), .ZN(n431) );
  INV_X1 U558 ( .A(n726), .ZN(n435) );
  NOR2_X1 U559 ( .A1(n364), .A2(n726), .ZN(n438) );
  OR2_X1 U560 ( .A1(n567), .A2(n460), .ZN(n439) );
  AND2_X1 U561 ( .A1(G224), .A2(n745), .ZN(n440) );
  NOR2_X1 U562 ( .A1(n753), .A2(n634), .ZN(n604) );
  INV_X1 U563 ( .A(n693), .ZN(n570) );
  XNOR2_X1 U564 ( .A(n557), .B(KEYINPUT90), .ZN(n555) );
  XNOR2_X1 U565 ( .A(n556), .B(n555), .ZN(n559) );
  INV_X1 U566 ( .A(KEYINPUT45), .ZN(n562) );
  XNOR2_X1 U567 ( .A(n508), .B(n446), .ZN(n732) );
  XNOR2_X1 U568 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X1 U569 ( .A1(n632), .A2(n730), .ZN(G63) );
  XNOR2_X1 U570 ( .A(n732), .B(n494), .ZN(n448) );
  NAND2_X1 U571 ( .A1(n723), .A2(n625), .ZN(n454) );
  NAND2_X1 U572 ( .A1(n510), .A2(n450), .ZN(n455) );
  NAND2_X1 U573 ( .A1(G210), .A2(n455), .ZN(n452) );
  NAND2_X1 U574 ( .A1(n455), .A2(G214), .ZN(n683) );
  NAND2_X1 U575 ( .A1(G952), .A2(n458), .ZN(n714) );
  NOR2_X1 U576 ( .A1(G953), .A2(n714), .ZN(n567) );
  INV_X1 U577 ( .A(G953), .ZN(n456) );
  NOR2_X1 U578 ( .A1(G898), .A2(n456), .ZN(n457) );
  XOR2_X1 U579 ( .A(KEYINPUT94), .B(n457), .Z(n734) );
  NAND2_X1 U580 ( .A1(G902), .A2(n458), .ZN(n565) );
  NOR2_X1 U581 ( .A1(n734), .A2(n565), .ZN(n459) );
  XOR2_X1 U582 ( .A(KEYINPUT95), .B(n459), .Z(n460) );
  INV_X1 U583 ( .A(KEYINPUT0), .ZN(n461) );
  XNOR2_X1 U584 ( .A(n462), .B(KEYINPUT7), .ZN(n466) );
  XNOR2_X1 U585 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U586 ( .A(n466), .B(n465), .Z(n469) );
  NAND2_X1 U587 ( .A1(n745), .A2(G234), .ZN(n467) );
  XOR2_X1 U588 ( .A(KEYINPUT8), .B(n467), .Z(n519) );
  NAND2_X1 U589 ( .A1(G217), .A2(n519), .ZN(n468) );
  XNOR2_X1 U590 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U591 ( .A(n470), .B(n471), .ZN(n629) );
  NAND2_X1 U592 ( .A1(n629), .A2(n510), .ZN(n473) );
  XNOR2_X1 U593 ( .A(KEYINPUT104), .B(G478), .ZN(n472) );
  XNOR2_X1 U594 ( .A(n473), .B(n472), .ZN(n539) );
  XNOR2_X1 U595 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n484) );
  XOR2_X1 U596 ( .A(n474), .B(KEYINPUT10), .Z(n518) );
  XOR2_X1 U597 ( .A(G140), .B(G104), .Z(n476) );
  XNOR2_X1 U598 ( .A(n476), .B(n475), .ZN(n478) );
  XOR2_X1 U599 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n477) );
  NAND2_X1 U600 ( .A1(G214), .A2(n504), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U602 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U603 ( .A(n518), .B(n483), .ZN(n644) );
  XNOR2_X1 U604 ( .A(n485), .B(G475), .ZN(n540) );
  INV_X1 U605 ( .A(n685), .ZN(n489) );
  NAND2_X1 U606 ( .A1(G234), .A2(n625), .ZN(n486) );
  XNOR2_X1 U607 ( .A(KEYINPUT20), .B(n486), .ZN(n521) );
  NAND2_X1 U608 ( .A1(n521), .A2(G221), .ZN(n488) );
  XOR2_X1 U609 ( .A(KEYINPUT98), .B(KEYINPUT21), .Z(n487) );
  XNOR2_X1 U610 ( .A(n488), .B(n487), .ZN(n693) );
  NAND2_X1 U611 ( .A1(n489), .A2(n693), .ZN(n490) );
  NOR2_X1 U612 ( .A1(n537), .A2(n490), .ZN(n492) );
  NAND2_X1 U613 ( .A1(n745), .A2(G227), .ZN(n496) );
  XNOR2_X1 U614 ( .A(n496), .B(G146), .ZN(n497) );
  XNOR2_X1 U615 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U616 ( .A(n744), .B(n499), .ZN(n652) );
  XNOR2_X1 U617 ( .A(KEYINPUT71), .B(G469), .ZN(n501) );
  INV_X1 U618 ( .A(KEYINPUT70), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U620 ( .A(n592), .ZN(n700) );
  NAND2_X1 U621 ( .A1(n504), .A2(G210), .ZN(n505) );
  NAND2_X1 U622 ( .A1(n637), .A2(n510), .ZN(n512) );
  INV_X1 U623 ( .A(G472), .ZN(n511) );
  XNOR2_X1 U624 ( .A(n696), .B(KEYINPUT6), .ZN(n549) );
  XNOR2_X1 U625 ( .A(G128), .B(G110), .ZN(n514) );
  XOR2_X1 U626 ( .A(KEYINPUT96), .B(KEYINPUT24), .Z(n517) );
  XNOR2_X1 U627 ( .A(G119), .B(KEYINPUT23), .ZN(n516) );
  NAND2_X1 U628 ( .A1(G221), .A2(n519), .ZN(n520) );
  NOR2_X1 U629 ( .A1(n729), .A2(G902), .ZN(n526) );
  XOR2_X1 U630 ( .A(KEYINPUT76), .B(KEYINPUT97), .Z(n523) );
  NAND2_X1 U631 ( .A1(n521), .A2(G217), .ZN(n522) );
  XNOR2_X1 U632 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U633 ( .A(KEYINPUT25), .B(n524), .ZN(n525) );
  XNOR2_X1 U634 ( .A(n564), .B(KEYINPUT106), .ZN(n692) );
  NAND2_X1 U635 ( .A1(n564), .A2(n693), .ZN(n699) );
  NOR2_X1 U636 ( .A1(n696), .A2(n699), .ZN(n527) );
  NAND2_X1 U637 ( .A1(n592), .A2(n527), .ZN(n704) );
  NOR2_X1 U638 ( .A1(n537), .A2(n704), .ZN(n528) );
  XNOR2_X1 U639 ( .A(n528), .B(KEYINPUT31), .ZN(n673) );
  INV_X1 U640 ( .A(n537), .ZN(n529) );
  NAND2_X1 U641 ( .A1(n531), .A2(n696), .ZN(n658) );
  INV_X1 U642 ( .A(n539), .ZN(n532) );
  AND2_X1 U643 ( .A1(n532), .A2(n540), .ZN(n669) );
  INV_X1 U644 ( .A(n669), .ZN(n671) );
  OR2_X1 U645 ( .A1(n540), .A2(n532), .ZN(n674) );
  NAND2_X1 U646 ( .A1(n671), .A2(n674), .ZN(n606) );
  NAND2_X1 U647 ( .A1(n533), .A2(n606), .ZN(n534) );
  NOR2_X1 U648 ( .A1(n346), .A2(n699), .ZN(n535) );
  NOR2_X1 U649 ( .A1(n537), .A2(n716), .ZN(n538) );
  XNOR2_X1 U650 ( .A(n538), .B(KEYINPUT34), .ZN(n542) );
  NAND2_X1 U651 ( .A1(n540), .A2(n539), .ZN(n584) );
  XNOR2_X1 U652 ( .A(n584), .B(KEYINPUT77), .ZN(n541) );
  NAND2_X1 U653 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U654 ( .A(n545), .B(KEYINPUT89), .ZN(n561) );
  NAND2_X1 U655 ( .A1(n577), .A2(n572), .ZN(n548) );
  NOR2_X1 U656 ( .A1(n546), .A2(n548), .ZN(n635) );
  NOR2_X1 U657 ( .A1(n692), .A2(n549), .ZN(n550) );
  NAND2_X1 U658 ( .A1(n550), .A2(n592), .ZN(n551) );
  OR2_X1 U659 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U660 ( .A(KEYINPUT32), .ZN(n553) );
  XNOR2_X1 U661 ( .A(n554), .B(n553), .ZN(n755) );
  NOR2_X1 U662 ( .A1(n635), .A2(n755), .ZN(n556) );
  INV_X1 U663 ( .A(KEYINPUT44), .ZN(n557) );
  NAND2_X1 U664 ( .A1(n557), .A2(n752), .ZN(n558) );
  NAND2_X1 U665 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U666 ( .A1(n561), .A2(n560), .ZN(n563) );
  NOR2_X1 U667 ( .A1(G900), .A2(n566), .ZN(n568) );
  INV_X1 U668 ( .A(n606), .ZN(n687) );
  NAND2_X1 U669 ( .A1(n687), .A2(KEYINPUT47), .ZN(n575) );
  INV_X1 U670 ( .A(n683), .ZN(n614) );
  OR2_X1 U671 ( .A1(n577), .A2(n614), .ZN(n579) );
  INV_X1 U672 ( .A(KEYINPUT30), .ZN(n578) );
  XNOR2_X1 U673 ( .A(n579), .B(n578), .ZN(n580) );
  NAND2_X1 U674 ( .A1(n599), .A2(n618), .ZN(n583) );
  XNOR2_X1 U675 ( .A(n585), .B(KEYINPUT84), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n346), .A2(n586), .ZN(n587) );
  XOR2_X1 U677 ( .A(KEYINPUT110), .B(n587), .Z(n588) );
  NOR2_X1 U678 ( .A1(n671), .A2(n588), .ZN(n589) );
  XNOR2_X1 U679 ( .A(KEYINPUT111), .B(n589), .ZN(n615) );
  NOR2_X1 U680 ( .A1(n347), .A2(n615), .ZN(n591) );
  XNOR2_X1 U681 ( .A(n591), .B(KEYINPUT36), .ZN(n593) );
  AND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n676) );
  NOR2_X1 U683 ( .A1(n594), .A2(n676), .ZN(n611) );
  INV_X1 U684 ( .A(KEYINPUT38), .ZN(n595) );
  XNOR2_X1 U685 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n597) );
  INV_X1 U686 ( .A(KEYINPUT72), .ZN(n600) );
  XNOR2_X1 U687 ( .A(n600), .B(KEYINPUT39), .ZN(n601) );
  XNOR2_X1 U688 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n602) );
  XNOR2_X1 U689 ( .A(n603), .B(n602), .ZN(n634) );
  XNOR2_X1 U690 ( .A(n604), .B(KEYINPUT46), .ZN(n609) );
  AND2_X1 U691 ( .A1(n606), .A2(n383), .ZN(n607) );
  NAND2_X1 U692 ( .A1(n605), .A2(n607), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n613) );
  XNOR2_X1 U694 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n616), .A2(n700), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n617), .B(KEYINPUT43), .ZN(n620) );
  INV_X1 U698 ( .A(n618), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n679) );
  OR2_X1 U700 ( .A1(n621), .A2(n674), .ZN(n633) );
  AND2_X1 U701 ( .A1(n679), .A2(n633), .ZN(n622) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n623) );
  NOR2_X2 U703 ( .A1(n363), .A2(n624), .ZN(n681) );
  NAND2_X1 U704 ( .A1(n364), .A2(G478), .ZN(n631) );
  INV_X1 U705 ( .A(n629), .ZN(n630) );
  INV_X1 U706 ( .A(n647), .ZN(n730) );
  XNOR2_X1 U707 ( .A(n633), .B(G134), .ZN(G36) );
  XOR2_X1 U708 ( .A(G131), .B(n634), .Z(G33) );
  XOR2_X1 U709 ( .A(G110), .B(n635), .Z(G12) );
  NAND2_X1 U710 ( .A1(n722), .A2(G472), .ZN(n639) );
  XOR2_X1 U711 ( .A(KEYINPUT115), .B(KEYINPUT62), .Z(n636) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n640), .A2(n647), .ZN(n642) );
  XOR2_X1 U714 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n722), .A2(G475), .ZN(n646) );
  XNOR2_X1 U717 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(G60) );
  NAND2_X1 U722 ( .A1(n364), .A2(G469), .ZN(n654) );
  XOR2_X1 U723 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U726 ( .A1(n655), .A2(n730), .ZN(G54) );
  XNOR2_X1 U727 ( .A(n348), .B(G101), .ZN(G3) );
  NOR2_X1 U728 ( .A1(n658), .A2(n671), .ZN(n657) );
  XOR2_X1 U729 ( .A(G104), .B(n657), .Z(G6) );
  NOR2_X1 U730 ( .A1(n658), .A2(n674), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n660) );
  XNOR2_X1 U732 ( .A(G107), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT116), .B(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G9) );
  XOR2_X1 U736 ( .A(KEYINPUT118), .B(KEYINPUT29), .Z(n666) );
  INV_X1 U737 ( .A(n674), .ZN(n664) );
  NAND2_X1 U738 ( .A1(n664), .A2(n605), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U740 ( .A(G128), .B(n667), .ZN(G30) );
  XOR2_X1 U741 ( .A(G143), .B(n668), .Z(G45) );
  NAND2_X1 U742 ( .A1(n605), .A2(n669), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n670), .B(G146), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n671), .A2(n673), .ZN(n672) );
  XOR2_X1 U745 ( .A(G113), .B(n672), .Z(G15) );
  NOR2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U747 ( .A(G116), .B(n675), .Z(G18) );
  XOR2_X1 U748 ( .A(KEYINPUT119), .B(KEYINPUT37), .Z(n678) );
  XNOR2_X1 U749 ( .A(G125), .B(n676), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n678), .B(n677), .ZN(G27) );
  XNOR2_X1 U751 ( .A(G140), .B(KEYINPUT120), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(G42) );
  NOR2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n688), .B(KEYINPUT122), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n691), .A2(n716), .ZN(n710) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n695) );
  XNOR2_X1 U760 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n695), .B(n694), .ZN(n698) );
  INV_X1 U762 ( .A(n696), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n703) );
  NAND2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U765 ( .A(n701), .B(KEYINPUT50), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U768 ( .A(KEYINPUT51), .B(n706), .ZN(n708) );
  INV_X1 U769 ( .A(n707), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n708), .A2(n717), .ZN(n709) );
  NOR2_X1 U771 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U772 ( .A(n711), .B(KEYINPUT52), .Z(n712) );
  XNOR2_X1 U773 ( .A(KEYINPUT123), .B(n712), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U775 ( .A(n715), .B(KEYINPUT124), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U777 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U778 ( .A(KEYINPUT53), .B(n721), .ZN(G75) );
  XNOR2_X1 U779 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n725) );
  XNOR2_X1 U780 ( .A(n723), .B(KEYINPUT83), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U782 ( .A(KEYINPUT56), .B(n727), .ZN(G51) );
  NAND2_X1 U783 ( .A1(n364), .A2(G217), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n731), .B(G101), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n742) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  AND2_X1 U789 ( .A1(n737), .A2(G898), .ZN(n740) );
  NOR2_X1 U790 ( .A1(G953), .A2(n363), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U793 ( .A(KEYINPUT126), .B(n743), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n744), .B(n518), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U796 ( .A(n747), .B(G227), .ZN(n748) );
  NAND2_X1 U797 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U800 ( .A(G122), .B(n752), .Z(G24) );
  XNOR2_X1 U801 ( .A(G137), .B(n753), .ZN(n754) );
  XNOR2_X1 U802 ( .A(n754), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U803 ( .A(G119), .B(n755), .Z(G21) );
endmodule

