//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(new_n468), .ZN(G160));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n459), .A2(G112), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n472), .A2(new_n473), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G138), .A4(new_n459), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n459), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n492), .A2(new_n496), .B1(new_n476), .B2(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT71), .B(G88), .Z(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n500), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n506), .A2(new_n505), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n518), .ZN(new_n524));
  OAI21_X1  g099(.A(G651), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n509), .A2(new_n510), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n504), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n537));
  AND3_X1   g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G89), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n503), .A2(G51), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n536), .A2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n530), .A2(new_n532), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n540), .A2(G90), .B1(new_n503), .B2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AOI22_X1  g128(.A1(new_n540), .A2(G81), .B1(new_n503), .B2(G43), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n547), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n555), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n503), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n521), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(new_n540), .B2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n566), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G166), .ZN(G303));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n547), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G87), .B2(new_n540), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n503), .A2(G49), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G288));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n509), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n514), .B2(new_n515), .ZN(new_n584));
  INV_X1    g159(.A(G73), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n500), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n503), .A2(G48), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n501), .A2(new_n502), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n589), .A2(new_n516), .A3(KEYINPUT77), .A4(G86), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n582), .A2(new_n587), .A3(new_n588), .A4(new_n590), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT78), .ZN(G305));
  AND2_X1   g167(.A1(new_n530), .A2(new_n532), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n512), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n503), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n509), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n509), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n521), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n503), .B2(G54), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(KEYINPUT79), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G299), .B2(new_n609), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n614), .B1(new_n613), .B2(new_n616), .ZN(G297));
  AOI21_X1  g192(.A(new_n614), .B1(new_n613), .B2(new_n616), .ZN(G280));
  INV_X1    g193(.A(new_n608), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR2_X1   g196(.A1(new_n608), .A2(G559), .ZN(new_n622));
  OR3_X1    g197(.A1(new_n622), .A2(KEYINPUT80), .A3(new_n609), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT80), .B1(new_n622), .B2(new_n609), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n623), .B(new_n624), .C1(G868), .C2(new_n559), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g201(.A1(new_n471), .A2(G2105), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n485), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n474), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n476), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n459), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT81), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  INV_X1    g218(.A(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(KEYINPUT86), .ZN(new_n655));
  INV_X1    g230(.A(new_n652), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT84), .ZN(new_n660));
  XOR2_X1   g235(.A(G2443), .B(G2446), .Z(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n653), .A2(new_n657), .A3(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(new_n666), .ZN(new_n672));
  AOI211_X1 g247(.A(KEYINPUT87), .B(new_n667), .C1(new_n664), .C2(new_n665), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(KEYINPUT17), .ZN(new_n682));
  INV_X1    g257(.A(new_n676), .ZN(new_n683));
  INV_X1    g258(.A(new_n677), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n679), .A3(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n678), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n681), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1961), .B(G1966), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n694), .B1(new_n699), .B2(KEYINPUT89), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(KEYINPUT89), .B2(new_n699), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n694), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n696), .A2(new_n698), .ZN(new_n704));
  MUX2_X1   g279(.A(new_n703), .B(new_n694), .S(new_n704), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT90), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT91), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n702), .A2(new_n708), .A3(new_n705), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n713), .B1(new_n710), .B2(new_n714), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n692), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n719), .A2(new_n691), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(G229));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n619), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G4), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1348), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(G164), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G27), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n724), .A2(new_n725), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n729), .A2(new_n730), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n726), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n727), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n474), .A2(G139), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n485), .A2(G127), .ZN(new_n740));
  NAND2_X1  g315(.A1(G115), .A2(G2104), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n459), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(new_n727), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G2072), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n727), .A2(G32), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n627), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n476), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(new_n727), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  INV_X1    g331(.A(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G160), .B2(new_n727), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G11), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT30), .B(G28), .Z(new_n764));
  NOR2_X1   g339(.A1(new_n636), .A2(new_n727), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n763), .B1(G29), .B2(new_n764), .C1(new_n765), .C2(KEYINPUT96), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(KEYINPUT96), .B2(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n745), .A2(new_n755), .A3(new_n762), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n722), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n722), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G1961), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n722), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n771), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n734), .A2(new_n768), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n727), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n727), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT29), .B(G2090), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n727), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n474), .A2(G140), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT92), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  INV_X1    g362(.A(G116), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G2105), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n476), .A2(G128), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT93), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n476), .A2(new_n792), .A3(G128), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n789), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n784), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2067), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n722), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n559), .B2(new_n722), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1341), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n782), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n722), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n722), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n778), .B(new_n802), .C1(G1966), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(G1966), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n722), .A2(G24), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n599), .B2(new_n722), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G1986), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(G1986), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n727), .A2(G25), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n474), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n476), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(G95), .A2(G2105), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n820), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n823), .B2(new_n727), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT35), .B(G1991), .Z(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n815), .A2(new_n816), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n722), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(G288), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n722), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT33), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1976), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n722), .A2(G22), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G166), .B2(new_n722), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1971), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT32), .B(G1981), .ZN(new_n838));
  MUX2_X1   g413(.A(G6), .B(G305), .S(G16), .Z(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n838), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n834), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n829), .B1(new_n842), .B2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n834), .A2(new_n840), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n811), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n811), .A3(new_n845), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n810), .B1(new_n847), .B2(new_n848), .ZN(G311));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n809), .B1(new_n850), .B2(new_n846), .ZN(G150));
  NAND3_X1  g426(.A1(new_n530), .A2(new_n532), .A3(G67), .ZN(new_n852));
  NAND2_X1  g427(.A1(G80), .A2(G543), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G651), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n503), .A2(G55), .ZN(new_n856));
  INV_X1    g431(.A(G93), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n509), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n619), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n855), .A2(new_n865), .A3(new_n859), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n512), .B1(new_n852), .B2(new_n853), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT97), .B1(new_n867), .B2(new_n858), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n866), .A2(new_n559), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n559), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n864), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n862), .B1(new_n874), .B2(new_n876), .ZN(G145));
  XOR2_X1   g452(.A(new_n498), .B(KEYINPUT98), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n795), .A2(new_n751), .ZN(new_n880));
  INV_X1    g455(.A(new_n743), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n752), .A2(new_n786), .A3(new_n794), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n743), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n878), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n474), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n476), .A2(G130), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n459), .A2(G118), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n629), .B(new_n895), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n823), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT99), .B1(new_n890), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n896), .B(new_n822), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n886), .A2(new_n889), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n886), .B2(new_n889), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n636), .B(G160), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n481), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n903), .A2(KEYINPUT100), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n907), .B1(new_n903), .B2(KEYINPUT100), .ZN(new_n911));
  AND4_X1   g486(.A1(KEYINPUT101), .A2(new_n902), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n884), .A2(new_n885), .A3(new_n879), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n878), .B1(new_n888), .B2(new_n883), .ZN(new_n914));
  OAI211_X1 g489(.A(KEYINPUT100), .B(new_n897), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n907), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(new_n909), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT101), .B1(new_n918), .B2(new_n902), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n908), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g496(.A1(new_n558), .A2(G651), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n554), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n865), .B1(new_n855), .B2(new_n859), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n867), .A2(KEYINPUT97), .A3(new_n858), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n866), .A2(new_n559), .A3(new_n868), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(new_n622), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n622), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n608), .A2(G299), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n603), .A2(new_n566), .A3(new_n570), .A4(new_n607), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT102), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n931), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n929), .A3(new_n930), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n937), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n599), .B(G166), .ZN(new_n949));
  XNOR2_X1  g524(.A(G305), .B(G288), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n599), .B(G303), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n831), .B(G305), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT42), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n948), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n937), .A2(KEYINPUT103), .A3(new_n939), .A4(new_n945), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n948), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n860), .A2(new_n609), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(G295));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n961), .ZN(G331));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  AND4_X1   g539(.A1(new_n536), .A2(new_n550), .A3(new_n543), .A4(new_n551), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n536), .A2(new_n543), .B1(new_n550), .B2(new_n551), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n928), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT104), .ZN(new_n969));
  NAND2_X1  g544(.A1(G286), .A2(G301), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n536), .A2(new_n550), .A3(new_n543), .A4(new_n551), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n934), .B1(new_n871), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n928), .A2(new_n967), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n927), .A3(new_n926), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n944), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n979), .A3(new_n955), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n968), .A2(new_n977), .A3(new_n935), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(new_n977), .A3(new_n975), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n944), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n964), .B(new_n980), .C1(new_n983), .C2(new_n955), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT105), .B1(new_n984), .B2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n944), .ZN(new_n986));
  INV_X1    g561(.A(new_n981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n955), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n980), .A2(new_n964), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n980), .A2(new_n964), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n955), .B1(new_n976), .B2(new_n979), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT43), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n985), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n995), .A2(new_n996), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n984), .A2(new_n993), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT44), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n498), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT106), .B(G40), .Z(new_n1010));
  NAND3_X1  g585(.A1(G160), .A2(KEYINPUT107), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G125), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n472), .B2(new_n473), .ZN(new_n1013));
  INV_X1    g588(.A(new_n463), .ZN(new_n1014));
  OAI21_X1  g589(.A(G2105), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n466), .B1(new_n474), .B2(G137), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n1010), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1009), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(G1996), .A3(new_n751), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT108), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n795), .B(new_n797), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G1996), .B2(new_n751), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n823), .A2(new_n825), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n822), .A2(new_n826), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1020), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n599), .B(G1986), .Z(new_n1030));
  AOI21_X1  g605(.A(new_n1029), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n488), .B2(new_n497), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT107), .B1(G160), .B2(new_n1010), .ZN(new_n1033));
  AND4_X1   g608(.A1(KEYINPUT107), .A2(new_n1015), .A3(new_n1016), .A4(new_n1010), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n574), .A2(G651), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n540), .A2(G87), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n578), .A3(G1976), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(G8), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1035), .A2(G8), .A3(new_n1038), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT112), .B(G1976), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n575), .B2(new_n578), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1040), .A2(KEYINPUT113), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n1047));
  NOR4_X1   g622(.A1(new_n1039), .A2(new_n1047), .A3(KEYINPUT52), .A4(new_n1044), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n582), .A2(new_n590), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n521), .A2(new_n583), .B1(new_n585), .B2(new_n500), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1052), .A2(G651), .B1(new_n503), .B2(G48), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1050), .A2(KEYINPUT114), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n591), .B2(G1981), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n588), .B1(new_n581), .B2(new_n509), .ZN(new_n1058));
  INV_X1    g633(.A(new_n587), .ZN(new_n1059));
  OAI21_X1  g634(.A(G1981), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1019), .A2(new_n1011), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1032), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT116), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n1062), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n1073), .A3(new_n1067), .A4(new_n1064), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1032), .A2(KEYINPUT45), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1009), .A2(new_n1066), .A3(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT109), .B(G1971), .Z(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1080));
  AOI22_X1  g655(.A1(new_n1011), .A2(new_n1019), .B1(new_n1032), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(G2090), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n520), .A2(new_n528), .A3(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT111), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1084), .A2(new_n1088), .A3(G8), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1049), .A2(new_n1075), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1080), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1007), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n1066), .C1(KEYINPUT50), .C2(new_n1007), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1079), .B1(G2090), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1065), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1079), .B(KEYINPUT117), .C1(G2090), .C2(new_n1097), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1087), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1009), .A2(new_n1076), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n730), .A3(new_n1066), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g681(.A(G1961), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1083), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G301), .B(KEYINPUT54), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1016), .A2(KEYINPUT53), .A3(G40), .A4(new_n730), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n462), .A2(KEYINPUT125), .A3(new_n463), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT125), .B1(new_n462), .B2(new_n463), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n459), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1104), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1104), .A2(KEYINPUT126), .A3(new_n1115), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1110), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1109), .A2(new_n1110), .B1(new_n1120), .B2(new_n1108), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1032), .A2(new_n1080), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1082), .A2(new_n1066), .A3(new_n761), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1966), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1077), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1081), .A2(KEYINPUT118), .A3(new_n761), .A4(new_n1082), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1126), .A2(new_n1128), .A3(G168), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1122), .B1(new_n1130), .B2(G8), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1129), .A3(new_n1128), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1122), .B1(new_n1132), .B2(G286), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(G8), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1103), .B(new_n1121), .C1(new_n1131), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n1138));
  INV_X1    g713(.A(G1996), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1009), .A2(new_n1066), .A3(new_n1139), .A4(new_n1076), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1035), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT122), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1138), .B1(new_n1147), .B2(new_n559), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1140), .A2(new_n1142), .A3(KEYINPUT122), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT122), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1138), .B(new_n559), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G299), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1956), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1033), .A2(new_n1034), .B1(new_n1032), .B2(new_n1080), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1007), .A2(KEYINPUT50), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1009), .A2(new_n1066), .A3(new_n1076), .A4(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1157), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1154), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1161), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT121), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1168), .A2(new_n1169), .A3(new_n1157), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1164), .A2(KEYINPUT61), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1137), .B1(new_n1153), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n559), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1151), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1171), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1169), .A2(new_n1157), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1168), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1176), .A2(new_n1179), .A3(KEYINPUT124), .A4(new_n1167), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1083), .A2(new_n725), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1066), .A2(new_n797), .A3(new_n1032), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1181), .B(new_n1182), .C1(KEYINPUT60), .C2(new_n619), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n619), .A2(KEYINPUT60), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1173), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n608), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1170), .B1(new_n1164), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1136), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT62), .B1(new_n1135), .B2(new_n1131), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1134), .A2(KEYINPUT51), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1191), .B(new_n1192), .C1(new_n1134), .C2(new_n1133), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1109), .A2(G171), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1103), .A2(new_n1190), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(G288), .A2(G1976), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1196), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1057), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1067), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1093), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n1075), .A3(new_n1049), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(G286), .A2(new_n1065), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1132), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT119), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1204), .B(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n1103), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1049), .A2(new_n1075), .A3(new_n1093), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1087), .B1(new_n1084), .B2(G8), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1208), .A2(new_n1206), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g787(.A(new_n1195), .B(new_n1202), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1031), .B1(new_n1189), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1020), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1023), .B2(new_n752), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT46), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1020), .A2(new_n1139), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT47), .Z(new_n1221));
  NAND2_X1  g796(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n786), .A2(new_n794), .A3(new_n797), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1215), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g799(.A1(new_n1215), .A2(G1986), .A3(G290), .ZN(new_n1225));
  XOR2_X1   g800(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1226));
  XNOR2_X1  g801(.A(new_n1225), .B(new_n1226), .ZN(new_n1227));
  NOR2_X1   g802(.A1(new_n1029), .A2(new_n1227), .ZN(new_n1228));
  NOR3_X1   g803(.A1(new_n1221), .A2(new_n1224), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1214), .A2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g805(.A(G319), .ZN(new_n1232));
  NOR2_X1   g806(.A1(G227), .A2(new_n1232), .ZN(new_n1233));
  AND4_X1   g807(.A1(new_n674), .A2(new_n720), .A3(new_n718), .A4(new_n1233), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n998), .A2(new_n1234), .A3(new_n920), .ZN(G225));
  INV_X1    g809(.A(G225), .ZN(G308));
endmodule


