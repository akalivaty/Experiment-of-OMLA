

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778;

  XNOR2_X1 U373 ( .A(G140), .B(G122), .ZN(n569) );
  XNOR2_X1 U374 ( .A(n523), .B(n460), .ZN(n758) );
  XNOR2_X1 U375 ( .A(n398), .B(n553), .ZN(n516) );
  XNOR2_X1 U376 ( .A(n461), .B(G146), .ZN(n523) );
  XNOR2_X1 U377 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X2 U378 ( .A(G953), .ZN(n769) );
  XNOR2_X2 U379 ( .A(n759), .B(n521), .ZN(n735) );
  XNOR2_X2 U380 ( .A(n400), .B(n611), .ZN(n775) );
  XNOR2_X1 U381 ( .A(n505), .B(n523), .ZN(n421) );
  NOR2_X2 U382 ( .A1(n775), .A2(n778), .ZN(n619) );
  NAND2_X2 U383 ( .A1(n427), .A2(n424), .ZN(n587) );
  XNOR2_X1 U384 ( .A(n516), .B(n421), .ZN(n420) );
  XOR2_X1 U385 ( .A(G137), .B(G140), .Z(n527) );
  NOR2_X1 U386 ( .A1(n768), .A2(KEYINPUT83), .ZN(n370) );
  NAND2_X1 U387 ( .A1(n375), .A2(n374), .ZN(n777) );
  AND2_X1 U388 ( .A1(n376), .A2(n430), .ZN(n375) );
  AND2_X1 U389 ( .A1(n579), .A2(n582), .ZN(n366) );
  XNOR2_X1 U390 ( .A(n382), .B(n381), .ZN(n717) );
  AND2_X1 U391 ( .A1(n429), .A2(n428), .ZN(n427) );
  OR2_X1 U392 ( .A1(n613), .A2(n355), .ZN(n635) );
  NOR2_X2 U393 ( .A1(n598), .A2(n687), .ZN(n693) );
  XNOR2_X1 U394 ( .A(n537), .B(n536), .ZN(n598) );
  XNOR2_X1 U395 ( .A(n422), .B(n420), .ZN(n726) );
  XNOR2_X1 U396 ( .A(n464), .B(n463), .ZN(n576) );
  AND2_X1 U397 ( .A1(n481), .A2(n480), .ZN(n479) );
  OR2_X1 U398 ( .A1(n740), .A2(G902), .ZN(n464) );
  INV_X1 U399 ( .A(n504), .ZN(n505) );
  XNOR2_X1 U400 ( .A(n744), .B(KEYINPUT75), .ZN(n520) );
  XNOR2_X1 U401 ( .A(n554), .B(KEYINPUT16), .ZN(n423) );
  XNOR2_X1 U402 ( .A(n495), .B(n494), .ZN(n744) );
  XNOR2_X1 U403 ( .A(n399), .B(G143), .ZN(n553) );
  XNOR2_X1 U404 ( .A(n496), .B(G104), .ZN(n495) );
  XNOR2_X1 U405 ( .A(n612), .B(KEYINPUT1), .ZN(n692) );
  AND2_X1 U406 ( .A1(n435), .A2(n434), .ZN(n415) );
  NAND2_X1 U407 ( .A1(n403), .A2(G217), .ZN(n653) );
  BUF_X1 U408 ( .A(n592), .Z(n634) );
  XNOR2_X2 U409 ( .A(KEYINPUT90), .B(G101), .ZN(n496) );
  XNOR2_X2 U410 ( .A(KEYINPUT66), .B(KEYINPUT70), .ZN(n397) );
  OR2_X1 U411 ( .A1(G902), .A2(G237), .ZN(n507) );
  INV_X1 U412 ( .A(n576), .ZN(n589) );
  NAND2_X1 U413 ( .A1(n402), .A2(n659), .ZN(n389) );
  NAND2_X1 U414 ( .A1(n777), .A2(n668), .ZN(n591) );
  INV_X1 U415 ( .A(G128), .ZN(n399) );
  INV_X1 U416 ( .A(G125), .ZN(n461) );
  XNOR2_X1 U417 ( .A(n416), .B(n361), .ZN(n414) );
  XNOR2_X1 U418 ( .A(n506), .B(n354), .ZN(n592) );
  NAND2_X2 U419 ( .A1(n479), .A2(n475), .ZN(n612) );
  NAND2_X1 U420 ( .A1(n478), .A2(n476), .ZN(n475) );
  AND2_X1 U421 ( .A1(n522), .A2(n477), .ZN(n476) );
  AND2_X1 U422 ( .A1(n615), .A2(n578), .ZN(n493) );
  XNOR2_X1 U423 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n528) );
  XNOR2_X1 U424 ( .A(n462), .B(n459), .ZN(n574) );
  INV_X1 U425 ( .A(n527), .ZN(n482) );
  AND2_X1 U426 ( .A1(n389), .A2(n448), .ZN(n447) );
  NOR2_X1 U427 ( .A1(n449), .A2(n742), .ZN(n448) );
  XOR2_X1 U428 ( .A(KEYINPUT5), .B(KEYINPUT78), .Z(n546) );
  XOR2_X1 U429 ( .A(n411), .B(G116), .Z(n542) );
  XNOR2_X1 U430 ( .A(G146), .B(G137), .ZN(n541) );
  XOR2_X1 U431 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n564) );
  NOR2_X1 U432 ( .A1(G953), .A2(G237), .ZN(n566) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT91), .ZN(n473) );
  XNOR2_X1 U434 ( .A(KEYINPUT82), .B(KEYINPUT17), .ZN(n471) );
  INV_X1 U435 ( .A(KEYINPUT88), .ZN(n373) );
  INV_X1 U436 ( .A(n701), .ZN(n380) );
  OR2_X1 U437 ( .A1(n658), .A2(G902), .ZN(n490) );
  NAND2_X1 U438 ( .A1(n659), .A2(n458), .ZN(n457) );
  INV_X1 U439 ( .A(n684), .ZN(n441) );
  INV_X1 U440 ( .A(KEYINPUT10), .ZN(n460) );
  XNOR2_X1 U441 ( .A(G128), .B(G110), .ZN(n524) );
  XNOR2_X1 U442 ( .A(n520), .B(n743), .ZN(n422) );
  INV_X1 U443 ( .A(n685), .ZN(n413) );
  NOR2_X1 U444 ( .A1(n585), .A2(n599), .ZN(n474) );
  INV_X1 U445 ( .A(KEYINPUT101), .ZN(n419) );
  XNOR2_X1 U446 ( .A(n401), .B(KEYINPUT39), .ZN(n643) );
  NAND2_X1 U447 ( .A1(n630), .A2(n702), .ZN(n401) );
  NAND2_X1 U448 ( .A1(n673), .A2(n701), .ZN(n364) );
  OR2_X1 U449 ( .A1(n439), .A2(n431), .ZN(n430) );
  NAND2_X1 U450 ( .A1(n426), .A2(n425), .ZN(n424) );
  XNOR2_X1 U451 ( .A(n575), .B(G475), .ZN(n463) );
  NAND2_X1 U452 ( .A1(n454), .A2(n453), .ZN(n452) );
  XOR2_X1 U453 ( .A(KEYINPUT99), .B(G134), .Z(n559) );
  INV_X1 U454 ( .A(KEYINPUT115), .ZN(n499) );
  NAND2_X2 U455 ( .A1(n415), .A2(n432), .ZN(n403) );
  NAND2_X1 U456 ( .A1(n651), .A2(KEYINPUT67), .ZN(n434) );
  XOR2_X1 U457 ( .A(G146), .B(G107), .Z(n518) );
  XOR2_X1 U458 ( .A(KEYINPUT89), .B(n654), .Z(n742) );
  NOR2_X1 U459 ( .A1(n443), .A2(n629), .ZN(n442) );
  XNOR2_X1 U460 ( .A(n369), .B(n368), .ZN(n640) );
  INV_X1 U461 ( .A(KEYINPUT77), .ZN(n368) );
  NAND2_X1 U462 ( .A1(n442), .A2(n444), .ZN(n369) );
  NAND2_X1 U463 ( .A1(n624), .A2(KEYINPUT84), .ZN(n444) );
  NAND2_X1 U464 ( .A1(n591), .A2(KEYINPUT68), .ZN(n378) );
  NOR2_X1 U465 ( .A1(n591), .A2(KEYINPUT68), .ZN(n409) );
  INV_X1 U466 ( .A(G469), .ZN(n477) );
  NAND2_X1 U467 ( .A1(G902), .A2(G469), .ZN(n480) );
  XNOR2_X1 U468 ( .A(n491), .B(n544), .ZN(n658) );
  XNOR2_X1 U469 ( .A(n549), .B(n543), .ZN(n491) );
  XNOR2_X1 U470 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U471 ( .A(G104), .B(G143), .Z(n570) );
  INV_X1 U472 ( .A(n758), .ZN(n459) );
  XNOR2_X1 U473 ( .A(n565), .B(n567), .ZN(n462) );
  XNOR2_X1 U474 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n563) );
  XNOR2_X1 U475 ( .A(n472), .B(n470), .ZN(n504) );
  XNOR2_X1 U476 ( .A(n471), .B(KEYINPUT81), .ZN(n470) );
  XNOR2_X1 U477 ( .A(n503), .B(n473), .ZN(n472) );
  INV_X1 U478 ( .A(KEYINPUT4), .ZN(n396) );
  INV_X1 U479 ( .A(KEYINPUT44), .ZN(n408) );
  NAND2_X1 U480 ( .A1(G237), .A2(G234), .ZN(n509) );
  NAND2_X1 U481 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U482 ( .A1(n513), .A2(n358), .ZN(n425) );
  NAND2_X1 U483 ( .A1(n692), .A2(n693), .ZN(n585) );
  NOR2_X1 U484 ( .A1(n603), .A2(n602), .ZN(n605) );
  INV_X1 U485 ( .A(G472), .ZN(n458) );
  XNOR2_X1 U486 ( .A(KEYINPUT79), .B(G110), .ZN(n494) );
  INV_X1 U487 ( .A(KEYINPUT41), .ZN(n381) );
  NOR2_X1 U488 ( .A1(n704), .A2(n380), .ZN(n379) );
  AND2_X1 U489 ( .A1(n393), .A2(n357), .ZN(n392) );
  INV_X1 U490 ( .A(KEYINPUT19), .ZN(n508) );
  NAND2_X1 U491 ( .A1(n592), .A2(n701), .ZN(n465) );
  NOR2_X1 U492 ( .A1(n613), .A2(n691), .ZN(n367) );
  NAND2_X1 U493 ( .A1(n612), .A2(n693), .ZN(n603) );
  XOR2_X1 U494 ( .A(n532), .B(n533), .Z(n652) );
  XNOR2_X1 U495 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U496 ( .A1(n418), .A2(n412), .ZN(n600) );
  XNOR2_X1 U497 ( .A(n635), .B(n419), .ZN(n418) );
  NOR2_X1 U498 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U499 ( .A(n484), .B(n483), .ZN(n774) );
  INV_X1 U500 ( .A(KEYINPUT35), .ZN(n483) );
  NAND2_X1 U501 ( .A1(n392), .A2(n390), .ZN(n484) );
  NAND2_X1 U502 ( .A1(n391), .A2(n350), .ZN(n390) );
  NAND2_X1 U503 ( .A1(n407), .A2(n404), .ZN(n374) );
  NOR2_X2 U504 ( .A1(n622), .A2(n621), .ZN(n674) );
  BUF_X1 U505 ( .A(n620), .Z(n621) );
  NOR2_X1 U506 ( .A1(n583), .A2(n406), .ZN(n405) );
  INV_X1 U507 ( .A(n691), .ZN(n406) );
  BUF_X1 U508 ( .A(G101), .Z(n411) );
  XNOR2_X1 U509 ( .A(n366), .B(n365), .ZN(n580) );
  INV_X1 U510 ( .A(KEYINPUT87), .ZN(n365) );
  NOR2_X1 U511 ( .A1(n456), .A2(n452), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n741), .B(n499), .ZN(n498) );
  INV_X1 U513 ( .A(KEYINPUT60), .ZN(n466) );
  NAND2_X1 U514 ( .A1(n468), .A2(n454), .ZN(n467) );
  XNOR2_X1 U515 ( .A(n737), .B(n736), .ZN(n738) );
  AND2_X1 U516 ( .A1(n587), .A2(n486), .ZN(n350) );
  XOR2_X1 U517 ( .A(n606), .B(KEYINPUT6), .Z(n586) );
  OR2_X1 U518 ( .A1(n582), .A2(n688), .ZN(n351) );
  AND2_X1 U519 ( .A1(n437), .A2(n487), .ZN(n352) );
  XOR2_X1 U520 ( .A(KEYINPUT3), .B(KEYINPUT74), .Z(n353) );
  AND2_X1 U521 ( .A1(G210), .A2(n507), .ZN(n354) );
  XNOR2_X1 U522 ( .A(n474), .B(KEYINPUT33), .ZN(n718) );
  NOR2_X1 U523 ( .A1(n590), .A2(n576), .ZN(n673) );
  OR2_X1 U524 ( .A1(n599), .A2(n364), .ZN(n355) );
  AND2_X1 U525 ( .A1(n389), .A2(n457), .ZN(n356) );
  AND2_X1 U526 ( .A1(n394), .A2(n485), .ZN(n357) );
  XOR2_X1 U527 ( .A(n514), .B(KEYINPUT0), .Z(n358) );
  INV_X1 U528 ( .A(G902), .ZN(n522) );
  INV_X1 U529 ( .A(n651), .ZN(n437) );
  XNOR2_X1 U530 ( .A(G902), .B(KEYINPUT15), .ZN(n651) );
  INV_X1 U531 ( .A(n742), .ZN(n454) );
  XOR2_X1 U532 ( .A(n740), .B(n739), .Z(n359) );
  XOR2_X1 U533 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n360) );
  XNOR2_X1 U534 ( .A(KEYINPUT48), .B(KEYINPUT73), .ZN(n361) );
  NOR2_X1 U535 ( .A1(n659), .A2(n458), .ZN(n362) );
  INV_X1 U536 ( .A(KEYINPUT67), .ZN(n487) );
  XNOR2_X1 U537 ( .A(KEYINPUT63), .B(KEYINPUT106), .ZN(n363) );
  NAND2_X1 U538 ( .A1(n774), .A2(n378), .ZN(n377) );
  XNOR2_X1 U539 ( .A(n591), .B(n373), .ZN(n372) );
  NAND2_X1 U540 ( .A1(n581), .A2(n660), .ZN(n410) );
  XNOR2_X1 U541 ( .A(n367), .B(KEYINPUT28), .ZN(n488) );
  NAND2_X1 U542 ( .A1(n370), .A2(n648), .ZN(n489) );
  XNOR2_X1 U543 ( .A(n469), .B(n359), .ZN(n468) );
  NAND2_X1 U544 ( .A1(n371), .A2(KEYINPUT68), .ZN(n385) );
  NAND2_X1 U545 ( .A1(n372), .A2(n774), .ZN(n371) );
  INV_X1 U546 ( .A(n584), .ZN(n407) );
  NAND2_X1 U547 ( .A1(n584), .A2(KEYINPUT32), .ZN(n376) );
  NAND2_X1 U548 ( .A1(n377), .A2(KEYINPUT44), .ZN(n383) );
  NAND2_X1 U549 ( .A1(n379), .A2(n702), .ZN(n382) );
  NOR2_X1 U550 ( .A1(n717), .A2(n622), .ZN(n616) );
  AND2_X1 U551 ( .A1(n384), .A2(n383), .ZN(n387) );
  NOR2_X1 U552 ( .A1(n409), .A2(n410), .ZN(n384) );
  NAND2_X1 U553 ( .A1(n385), .A2(n408), .ZN(n388) );
  XNOR2_X2 U554 ( .A(n386), .B(n360), .ZN(n648) );
  NAND2_X1 U555 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U556 ( .A1(n718), .A2(n588), .ZN(n393) );
  INV_X1 U557 ( .A(n718), .ZN(n391) );
  NAND2_X1 U558 ( .A1(n395), .A2(n588), .ZN(n394) );
  INV_X1 U559 ( .A(n587), .ZN(n395) );
  NAND2_X1 U560 ( .A1(n643), .A2(n673), .ZN(n400) );
  NAND2_X1 U561 ( .A1(n403), .A2(G475), .ZN(n469) );
  INV_X1 U562 ( .A(n403), .ZN(n402) );
  NAND2_X1 U563 ( .A1(n403), .A2(G469), .ZN(n737) );
  NAND2_X1 U564 ( .A1(n403), .A2(G478), .ZN(n500) );
  AND2_X1 U565 ( .A1(n403), .A2(n362), .ZN(n456) );
  AND2_X1 U566 ( .A1(n439), .A2(n431), .ZN(n404) );
  NAND2_X1 U567 ( .A1(n407), .A2(n405), .ZN(n668) );
  NAND2_X1 U568 ( .A1(n587), .A2(n493), .ZN(n492) );
  NAND2_X1 U569 ( .A1(n414), .A2(n440), .ZN(n768) );
  INV_X1 U570 ( .A(n631), .ZN(n485) );
  BUF_X1 U571 ( .A(n692), .Z(n412) );
  XNOR2_X2 U572 ( .A(n501), .B(G116), .ZN(n554) );
  XNOR2_X2 U573 ( .A(G107), .B(G122), .ZN(n501) );
  NAND2_X1 U574 ( .A1(n414), .A2(n413), .ZN(n647) );
  XNOR2_X2 U575 ( .A(n423), .B(n548), .ZN(n743) );
  NAND2_X1 U576 ( .A1(n433), .A2(n352), .ZN(n432) );
  XNOR2_X2 U577 ( .A(n636), .B(KEYINPUT38), .ZN(n702) );
  NAND2_X1 U578 ( .A1(n641), .A2(n642), .ZN(n416) );
  NOR2_X2 U579 ( .A1(n731), .A2(n742), .ZN(n733) );
  NAND2_X1 U580 ( .A1(n417), .A2(G210), .ZN(n730) );
  XNOR2_X1 U581 ( .A(n436), .B(KEYINPUT67), .ZN(n417) );
  NOR2_X1 U582 ( .A1(n685), .A2(n441), .ZN(n440) );
  XNOR2_X2 U583 ( .A(n502), .B(n353), .ZN(n548) );
  XNOR2_X1 U584 ( .A(n730), .B(n729), .ZN(n731) );
  INV_X1 U585 ( .A(n620), .ZN(n426) );
  NAND2_X1 U586 ( .A1(n513), .A2(n358), .ZN(n428) );
  NAND2_X1 U587 ( .A1(n620), .A2(n358), .ZN(n429) );
  XNOR2_X2 U588 ( .A(n465), .B(n508), .ZN(n620) );
  INV_X1 U589 ( .A(KEYINPUT32), .ZN(n431) );
  NAND2_X1 U590 ( .A1(n433), .A2(n437), .ZN(n436) );
  INV_X1 U591 ( .A(n721), .ZN(n433) );
  NAND2_X1 U592 ( .A1(n721), .A2(KEYINPUT67), .ZN(n435) );
  NAND2_X1 U593 ( .A1(n650), .A2(n438), .ZN(n721) );
  NAND2_X1 U594 ( .A1(n648), .A2(n649), .ZN(n438) );
  NOR2_X1 U595 ( .A1(n351), .A2(n586), .ZN(n439) );
  XNOR2_X1 U596 ( .A(n605), .B(n604), .ZN(n610) );
  NAND2_X1 U597 ( .A1(n726), .A2(n651), .ZN(n506) );
  NAND2_X1 U598 ( .A1(n627), .A2(n672), .ZN(n443) );
  NAND2_X1 U599 ( .A1(n445), .A2(n363), .ZN(n455) );
  NAND2_X1 U600 ( .A1(n447), .A2(n446), .ZN(n445) );
  INV_X1 U601 ( .A(n456), .ZN(n446) );
  INV_X1 U602 ( .A(n457), .ZN(n449) );
  NAND2_X1 U603 ( .A1(n455), .A2(n450), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n451), .A2(n356), .ZN(n450) );
  INV_X1 U605 ( .A(n363), .ZN(n453) );
  XNOR2_X1 U606 ( .A(n467), .B(n466), .ZN(G60) );
  NOR2_X2 U607 ( .A1(n610), .A2(n609), .ZN(n630) );
  XNOR2_X1 U608 ( .A(n574), .B(n573), .ZN(n740) );
  INV_X1 U609 ( .A(n735), .ZN(n478) );
  NAND2_X1 U610 ( .A1(n735), .A2(G469), .ZN(n481) );
  XNOR2_X2 U611 ( .A(n544), .B(n482), .ZN(n759) );
  XNOR2_X2 U612 ( .A(n516), .B(n515), .ZN(n544) );
  INV_X1 U613 ( .A(n588), .ZN(n486) );
  NAND2_X1 U614 ( .A1(n614), .A2(n488), .ZN(n622) );
  NAND2_X1 U615 ( .A1(n489), .A2(n644), .ZN(n650) );
  XNOR2_X2 U616 ( .A(n490), .B(G472), .ZN(n606) );
  XNOR2_X2 U617 ( .A(n492), .B(KEYINPUT22), .ZN(n584) );
  NOR2_X1 U618 ( .A1(n497), .A2(n742), .ZN(G63) );
  XNOR2_X1 U619 ( .A(n500), .B(n498), .ZN(n497) );
  XNOR2_X1 U620 ( .A(n520), .B(n519), .ZN(n521) );
  INV_X1 U621 ( .A(n681), .ZN(n639) );
  XNOR2_X1 U622 ( .A(n568), .B(G134), .ZN(n515) );
  INV_X1 U623 ( .A(KEYINPUT69), .ZN(n514) );
  INV_X1 U624 ( .A(KEYINPUT80), .ZN(n604) );
  XNOR2_X1 U625 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U626 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U627 ( .A(G119), .B(G113), .ZN(n502) );
  NAND2_X1 U628 ( .A1(G224), .A2(n769), .ZN(n503) );
  NAND2_X1 U629 ( .A1(G214), .A2(n507), .ZN(n701) );
  XNOR2_X1 U630 ( .A(n509), .B(KEYINPUT14), .ZN(n510) );
  NAND2_X1 U631 ( .A1(G952), .A2(n510), .ZN(n716) );
  NOR2_X1 U632 ( .A1(G953), .A2(n716), .ZN(n596) );
  NAND2_X1 U633 ( .A1(n510), .A2(G902), .ZN(n511) );
  XOR2_X1 U634 ( .A(n511), .B(KEYINPUT93), .Z(n593) );
  XOR2_X1 U635 ( .A(G898), .B(KEYINPUT92), .Z(n751) );
  NAND2_X1 U636 ( .A1(G953), .A2(n751), .ZN(n747) );
  NOR2_X1 U637 ( .A1(n593), .A2(n747), .ZN(n512) );
  NOR2_X1 U638 ( .A1(n596), .A2(n512), .ZN(n513) );
  XOR2_X1 U639 ( .A(KEYINPUT72), .B(G131), .Z(n568) );
  NAND2_X1 U640 ( .A1(G227), .A2(n769), .ZN(n517) );
  XOR2_X1 U641 ( .A(n518), .B(n517), .Z(n519) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(G119), .Z(n525) );
  XNOR2_X1 U643 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U644 ( .A(n758), .B(n526), .ZN(n533) );
  XOR2_X1 U645 ( .A(KEYINPUT24), .B(n527), .Z(n531) );
  NAND2_X1 U646 ( .A1(n769), .A2(G234), .ZN(n529) );
  XNOR2_X1 U647 ( .A(n529), .B(n528), .ZN(n557) );
  NAND2_X1 U648 ( .A1(G221), .A2(n557), .ZN(n530) );
  XNOR2_X1 U649 ( .A(n531), .B(n530), .ZN(n532) );
  NOR2_X1 U650 ( .A1(G902), .A2(n652), .ZN(n537) );
  NAND2_X1 U651 ( .A1(G234), .A2(n651), .ZN(n534) );
  XNOR2_X1 U652 ( .A(KEYINPUT20), .B(n534), .ZN(n538) );
  NAND2_X1 U653 ( .A1(n538), .A2(G217), .ZN(n535) );
  XOR2_X1 U654 ( .A(KEYINPUT25), .B(n535), .Z(n536) );
  NAND2_X1 U655 ( .A1(n538), .A2(G221), .ZN(n539) );
  XNOR2_X1 U656 ( .A(n539), .B(KEYINPUT21), .ZN(n687) );
  NOR2_X1 U657 ( .A1(n395), .A2(n603), .ZN(n540) );
  XNOR2_X1 U658 ( .A(n540), .B(KEYINPUT94), .ZN(n550) );
  XNOR2_X1 U659 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U660 ( .A1(G210), .A2(n566), .ZN(n545) );
  XNOR2_X1 U661 ( .A(n546), .B(n545), .ZN(n547) );
  INV_X1 U662 ( .A(n606), .ZN(n691) );
  NAND2_X1 U663 ( .A1(n550), .A2(n691), .ZN(n665) );
  NOR2_X1 U664 ( .A1(n691), .A2(n585), .ZN(n698) );
  NAND2_X1 U665 ( .A1(n587), .A2(n698), .ZN(n551) );
  XNOR2_X1 U666 ( .A(n551), .B(KEYINPUT95), .ZN(n552) );
  XNOR2_X1 U667 ( .A(KEYINPUT31), .B(n552), .ZN(n678) );
  NAND2_X1 U668 ( .A1(n665), .A2(n678), .ZN(n577) );
  XOR2_X1 U669 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n556) );
  XNOR2_X1 U670 ( .A(n553), .B(n554), .ZN(n555) );
  XNOR2_X1 U671 ( .A(n556), .B(n555), .ZN(n561) );
  NAND2_X1 U672 ( .A1(G217), .A2(n557), .ZN(n558) );
  XNOR2_X1 U673 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U674 ( .A(n561), .B(n560), .ZN(n741) );
  NOR2_X1 U675 ( .A1(n741), .A2(G902), .ZN(n562) );
  XOR2_X1 U676 ( .A(n562), .B(G478), .Z(n590) );
  XNOR2_X1 U677 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U678 ( .A1(n566), .A2(G214), .ZN(n567) );
  XNOR2_X1 U679 ( .A(n568), .B(G113), .ZN(n572) );
  XNOR2_X1 U680 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U681 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n575) );
  INV_X1 U682 ( .A(n673), .ZN(n676) );
  NAND2_X1 U683 ( .A1(n590), .A2(n576), .ZN(n679) );
  NAND2_X1 U684 ( .A1(n676), .A2(n679), .ZN(n628) );
  NAND2_X1 U685 ( .A1(n577), .A2(n628), .ZN(n581) );
  INV_X1 U686 ( .A(n692), .ZN(n582) );
  NOR2_X1 U687 ( .A1(n589), .A2(n590), .ZN(n615) );
  INV_X1 U688 ( .A(n687), .ZN(n578) );
  NOR2_X1 U689 ( .A1(n586), .A2(n584), .ZN(n579) );
  XOR2_X1 U690 ( .A(KEYINPUT100), .B(n598), .Z(n688) );
  NAND2_X1 U691 ( .A1(n580), .A2(n688), .ZN(n660) );
  INV_X1 U692 ( .A(n586), .ZN(n599) );
  NAND2_X1 U693 ( .A1(n598), .A2(n582), .ZN(n583) );
  XNOR2_X1 U694 ( .A(KEYINPUT76), .B(KEYINPUT34), .ZN(n588) );
  NAND2_X1 U695 ( .A1(n590), .A2(n589), .ZN(n631) );
  OR2_X1 U696 ( .A1(n593), .A2(n769), .ZN(n594) );
  NOR2_X1 U697 ( .A1(G900), .A2(n594), .ZN(n595) );
  NOR2_X1 U698 ( .A1(n596), .A2(n595), .ZN(n602) );
  NOR2_X1 U699 ( .A1(n602), .A2(n687), .ZN(n597) );
  NAND2_X1 U700 ( .A1(n598), .A2(n597), .ZN(n613) );
  XNOR2_X1 U701 ( .A(n600), .B(KEYINPUT43), .ZN(n601) );
  NOR2_X1 U702 ( .A1(n634), .A2(n601), .ZN(n685) );
  XOR2_X1 U703 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n611) );
  NAND2_X1 U704 ( .A1(n701), .A2(n606), .ZN(n607) );
  XNOR2_X1 U705 ( .A(n607), .B(KEYINPUT102), .ZN(n608) );
  XNOR2_X1 U706 ( .A(KEYINPUT30), .B(n608), .ZN(n609) );
  INV_X1 U707 ( .A(n634), .ZN(n636) );
  XOR2_X1 U708 ( .A(KEYINPUT103), .B(n612), .Z(n614) );
  INV_X1 U709 ( .A(n615), .ZN(n704) );
  XNOR2_X1 U710 ( .A(n616), .B(KEYINPUT42), .ZN(n778) );
  XNOR2_X1 U711 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n617) );
  XNOR2_X1 U712 ( .A(n617), .B(KEYINPUT64), .ZN(n618) );
  XNOR2_X1 U713 ( .A(n619), .B(n618), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n628), .A2(n674), .ZN(n623) );
  XNOR2_X1 U715 ( .A(n623), .B(KEYINPUT47), .ZN(n624) );
  INV_X1 U716 ( .A(KEYINPUT84), .ZN(n626) );
  NAND2_X1 U717 ( .A1(KEYINPUT47), .A2(n674), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n626), .A2(n625), .ZN(n627) );
  INV_X1 U719 ( .A(n628), .ZN(n707) );
  NOR2_X1 U720 ( .A1(n707), .A2(KEYINPUT84), .ZN(n629) );
  INV_X1 U721 ( .A(n630), .ZN(n632) );
  NOR2_X1 U722 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n634), .A2(n633), .ZN(n672) );
  XNOR2_X1 U724 ( .A(n637), .B(KEYINPUT36), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n638), .A2(n412), .ZN(n681) );
  NOR2_X1 U726 ( .A1(n640), .A2(n639), .ZN(n641) );
  INV_X1 U727 ( .A(n679), .ZN(n669) );
  NAND2_X1 U728 ( .A1(n643), .A2(n669), .ZN(n684) );
  INV_X1 U729 ( .A(KEYINPUT2), .ZN(n644) );
  XOR2_X1 U730 ( .A(n684), .B(KEYINPUT83), .Z(n645) );
  NAND2_X1 U731 ( .A1(n645), .A2(KEYINPUT2), .ZN(n646) );
  NOR2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X1 U734 ( .A1(G952), .A2(n769), .ZN(n654) );
  NOR2_X2 U735 ( .A1(n655), .A2(n742), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT116), .ZN(G66) );
  XOR2_X1 U737 ( .A(KEYINPUT105), .B(KEYINPUT62), .Z(n657) );
  XNOR2_X1 U738 ( .A(n660), .B(n411), .ZN(G3) );
  NOR2_X1 U739 ( .A1(n676), .A2(n665), .ZN(n662) );
  XNOR2_X1 U740 ( .A(G104), .B(KEYINPUT107), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(G6) );
  XOR2_X1 U742 ( .A(KEYINPUT108), .B(KEYINPUT26), .Z(n664) );
  XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT27), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n664), .B(n663), .ZN(n667) );
  NOR2_X1 U745 ( .A1(n679), .A2(n665), .ZN(n666) );
  XOR2_X1 U746 ( .A(n667), .B(n666), .Z(G9) );
  XNOR2_X1 U747 ( .A(G110), .B(n668), .ZN(G12) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U749 ( .A1(n669), .A2(n674), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(G30) );
  XNOR2_X1 U751 ( .A(G143), .B(n672), .ZN(G45) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U753 ( .A(n675), .B(G146), .ZN(G48) );
  NOR2_X1 U754 ( .A1(n676), .A2(n678), .ZN(n677) );
  XOR2_X1 U755 ( .A(G113), .B(n677), .Z(G15) );
  NOR2_X1 U756 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U757 ( .A(G116), .B(n680), .Z(G18) );
  XNOR2_X1 U758 ( .A(KEYINPUT37), .B(KEYINPUT109), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U760 ( .A(G125), .B(n683), .ZN(G27) );
  XNOR2_X1 U761 ( .A(G134), .B(n684), .ZN(G36) );
  XOR2_X1 U762 ( .A(n685), .B(G140), .Z(n686) );
  XNOR2_X1 U763 ( .A(KEYINPUT110), .B(n686), .ZN(G42) );
  NOR2_X1 U764 ( .A1(n688), .A2(n578), .ZN(n689) );
  XNOR2_X1 U765 ( .A(n689), .B(KEYINPUT49), .ZN(n690) );
  NAND2_X1 U766 ( .A1(n691), .A2(n690), .ZN(n696) );
  NOR2_X1 U767 ( .A1(n693), .A2(n412), .ZN(n694) );
  XNOR2_X1 U768 ( .A(n694), .B(KEYINPUT50), .ZN(n695) );
  NOR2_X1 U769 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U770 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U771 ( .A(KEYINPUT51), .B(n699), .Z(n700) );
  NOR2_X1 U772 ( .A1(n717), .A2(n700), .ZN(n713) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U775 ( .A(KEYINPUT111), .B(n705), .Z(n710) );
  NOR2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U777 ( .A(KEYINPUT112), .B(n708), .ZN(n709) );
  NOR2_X1 U778 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U779 ( .A1(n711), .A2(n718), .ZN(n712) );
  NOR2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U781 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U786 ( .A1(G953), .A2(n723), .ZN(n724) );
  XOR2_X1 U787 ( .A(KEYINPUT53), .B(n724), .Z(n725) );
  XNOR2_X1 U788 ( .A(KEYINPUT113), .B(n725), .ZN(G75) );
  INV_X1 U789 ( .A(n726), .ZN(n728) );
  XOR2_X1 U790 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n727) );
  XOR2_X1 U791 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n732) );
  XNOR2_X1 U792 ( .A(n733), .B(n732), .ZN(G51) );
  XOR2_X1 U793 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n734) );
  XNOR2_X1 U794 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U795 ( .A1(n742), .A2(n738), .ZN(G54) );
  XOR2_X1 U796 ( .A(KEYINPUT114), .B(KEYINPUT59), .Z(n739) );
  XNOR2_X1 U797 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U798 ( .A(n745), .B(KEYINPUT119), .ZN(n746) );
  NAND2_X1 U799 ( .A1(n747), .A2(n746), .ZN(n756) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n748), .B(KEYINPUT117), .ZN(n749) );
  XNOR2_X1 U802 ( .A(n749), .B(KEYINPUT61), .ZN(n750) );
  NOR2_X1 U803 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n648), .A2(n769), .ZN(n752) );
  XOR2_X1 U805 ( .A(KEYINPUT118), .B(n752), .Z(n753) );
  NOR2_X1 U806 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U808 ( .A(KEYINPUT120), .B(n757), .ZN(G69) );
  XOR2_X1 U809 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n761) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n761), .B(n760), .ZN(n766) );
  XNOR2_X1 U812 ( .A(G227), .B(n766), .ZN(n762) );
  NAND2_X1 U813 ( .A1(n762), .A2(G900), .ZN(n763) );
  XOR2_X1 U814 ( .A(KEYINPUT124), .B(n763), .Z(n764) );
  NOR2_X1 U815 ( .A1(n769), .A2(n764), .ZN(n765) );
  XNOR2_X1 U816 ( .A(n765), .B(KEYINPUT125), .ZN(n772) );
  XOR2_X1 U817 ( .A(n766), .B(KEYINPUT123), .Z(n767) );
  XNOR2_X1 U818 ( .A(n768), .B(n767), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U821 ( .A(KEYINPUT126), .B(n773), .ZN(G72) );
  XNOR2_X1 U822 ( .A(n774), .B(G122), .ZN(G24) );
  XNOR2_X1 U823 ( .A(n775), .B(G131), .ZN(n776) );
  XNOR2_X1 U824 ( .A(n776), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U825 ( .A(n777), .B(G119), .ZN(G21) );
  XOR2_X1 U826 ( .A(G137), .B(n778), .Z(G39) );
endmodule

