//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT85), .ZN(new_n203));
  XOR2_X1   g002(.A(G169gat), .B(G197gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT12), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT14), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G50gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(G43gat), .A2(G50gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n218), .B2(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n224), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n226), .A2(new_n215), .A3(new_n221), .A4(new_n222), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT87), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n232), .A3(G1gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G8gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n233), .A2(new_n234), .B1(new_n237), .B2(new_n231), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n236), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT17), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n230), .A2(new_n240), .A3(new_n243), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n228), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT18), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n225), .A2(new_n227), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n240), .A3(new_n243), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n254), .A2(new_n240), .A3(KEYINPUT88), .A4(new_n243), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n247), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n248), .B(KEYINPUT13), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT89), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n253), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n210), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n259), .A2(new_n263), .A3(new_n260), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n263), .B1(new_n259), .B2(new_n260), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT86), .B(new_n209), .C1(new_n270), .C2(new_n253), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT73), .B(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n279), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT27), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT27), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G183gat), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n286), .A2(new_n288), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n296), .A3(KEYINPUT28), .A4(new_n289), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT66), .B1(new_n290), .B2(new_n291), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n290), .A2(KEYINPUT65), .A3(new_n291), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n294), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n307), .A2(KEYINPUT24), .ZN(new_n310));
  XOR2_X1   g109(.A(G183gat), .B(G190gat), .Z(new_n311));
  AOI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(KEYINPUT24), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(KEYINPUT23), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n301), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n312), .A2(KEYINPUT64), .A3(new_n317), .A4(KEYINPUT25), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n313), .A2(new_n319), .A3(new_n315), .A4(new_n301), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT25), .ZN(new_n321));
  INV_X1    g120(.A(new_n310), .ZN(new_n322));
  XNOR2_X1  g121(.A(G183gat), .B(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G226gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n300), .A2(new_n308), .B1(new_n318), .B2(new_n326), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n331), .A2(KEYINPUT29), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n284), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(KEYINPUT29), .B2(new_n331), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n329), .B2(new_n330), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n283), .ZN(new_n339));
  XNOR2_X1  g138(.A(G64gat), .B(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT76), .B(G36gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT75), .B(G8gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n336), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n336), .A2(new_n339), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n344), .B(KEYINPUT77), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n346), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354));
  XNOR2_X1  g153(.A(G141gat), .B(G148gat), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(KEYINPUT2), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n356), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n360), .B(new_n359), .C1(new_n355), .C2(KEYINPUT2), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G127gat), .B(G134gat), .Z(new_n367));
  INV_X1    g166(.A(G113gat), .ZN(new_n368));
  INV_X1    g167(.A(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G113gat), .A2(G120gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n367), .A2(new_n372), .A3(KEYINPUT1), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n375));
  AND2_X1   g174(.A1(G113gat), .A2(G120gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(G113gat), .A2(G120gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n370), .A2(KEYINPUT67), .A3(new_n371), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n381), .A2(KEYINPUT68), .A3(new_n367), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT68), .B1(new_n381), .B2(new_n367), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n366), .B(new_n374), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n354), .B1(new_n384), .B2(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n367), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(KEYINPUT68), .A3(new_n367), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n373), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n390), .A2(KEYINPUT78), .A3(new_n391), .A4(new_n366), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n374), .B1(new_n382), .B2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n366), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  OR3_X1    g201(.A1(new_n390), .A2(KEYINPUT79), .A3(new_n366), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n365), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT79), .A3(new_n384), .ZN(new_n405));
  INV_X1    g204(.A(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(KEYINPUT5), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n366), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n393), .A3(KEYINPUT80), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n384), .A2(new_n412), .A3(KEYINPUT4), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n401), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G57gat), .ZN(new_n417));
  INV_X1    g216(.A(G85gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n408), .A2(new_n414), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n408), .B2(new_n414), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n421), .B(new_n419), .C1(new_n408), .C2(new_n414), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n353), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(G22gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n366), .B2(new_n396), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n283), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT3), .B1(new_n283), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n366), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n431), .B(KEYINPUT81), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n280), .B1(new_n277), .B2(new_n278), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n277), .A2(new_n280), .A3(new_n278), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT82), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n366), .B1(new_n444), .B2(new_n396), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n437), .B1(new_n445), .B2(new_n430), .ZN(new_n446));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT31), .B(G50gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n435), .B2(new_n446), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n428), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n446), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n427), .A3(new_n451), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n333), .B2(new_n390), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n306), .A2(new_n307), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n297), .A2(new_n298), .ZN(new_n462));
  INV_X1    g261(.A(new_n299), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT65), .B1(new_n290), .B2(new_n291), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n318), .A2(new_n326), .ZN(new_n467));
  OAI211_X1 g266(.A(KEYINPUT69), .B(new_n395), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G227gat), .A2(G233gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n333), .A2(new_n390), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n460), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n474), .A3(KEYINPUT34), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT32), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n468), .A3(new_n470), .ZN(new_n479));
  INV_X1    g278(.A(new_n469), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G43gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G71gat), .B(G99gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n481), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  AOI221_X4 g288(.A(new_n478), .B1(new_n489), .B2(new_n483), .C1(new_n479), .C2(new_n480), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n477), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n480), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n482), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n489), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n481), .B1(new_n484), .B2(new_n487), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n474), .B1(new_n471), .B2(KEYINPUT34), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n471), .A2(KEYINPUT34), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n475), .A4(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n458), .A2(new_n491), .A3(new_n500), .A4(KEYINPUT35), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n426), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n491), .A2(new_n500), .A3(KEYINPUT72), .ZN(new_n503));
  INV_X1    g302(.A(new_n477), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n496), .A4(new_n495), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n408), .A2(new_n414), .ZN(new_n508));
  INV_X1    g307(.A(new_n419), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n421), .A3(new_n420), .ZN(new_n511));
  INV_X1    g310(.A(new_n425), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n352), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n513), .A3(new_n458), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n502), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n503), .A2(new_n517), .A3(new_n506), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n491), .A2(new_n500), .A3(KEYINPUT36), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n458), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n426), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n410), .A2(new_n399), .A3(new_n413), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n406), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n403), .A2(new_n405), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n526), .B2(new_n400), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n525), .A3(new_n406), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n419), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT40), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n528), .A2(KEYINPUT40), .A3(new_n419), .A4(new_n529), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n510), .A3(new_n352), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n512), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n348), .A2(KEYINPUT37), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n336), .A2(new_n339), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT38), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n349), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n344), .B1(new_n348), .B2(KEYINPUT37), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n542), .A2(new_n538), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n345), .B(new_n541), .C1(new_n543), .C2(new_n539), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n534), .B(new_n458), .C1(new_n535), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n520), .A2(new_n522), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n273), .B1(new_n516), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G134gat), .B(G162gat), .Z(new_n548));
  AOI21_X1  g347(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT7), .ZN(new_n552));
  XNOR2_X1  g351(.A(G99gat), .B(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(G92gat), .ZN(new_n555));
  AOI22_X1  g354(.A1(KEYINPUT8), .A2(new_n554), .B1(new_n418), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(new_n552), .B2(new_n556), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n230), .A2(new_n244), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n560), .B2(new_n254), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n550), .B1(new_n570), .B2(KEYINPUT94), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n567), .B(new_n568), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(G57gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT92), .B(G57gat), .Z(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n575), .ZN(new_n578));
  XOR2_X1   g377(.A(G71gat), .B(G78gat), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT9), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT90), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n578), .A2(new_n580), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G57gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G64gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n584), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n591), .A2(KEYINPUT91), .A3(new_n579), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT91), .B1(new_n591), .B2(new_n579), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n240), .B(new_n243), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G183gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n595), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G211gat), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n601), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT98), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n594), .A2(new_n560), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n559), .B(new_n587), .C1(new_n593), .C2(new_n592), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n594), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(KEYINPUT95), .A3(new_n559), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G176gat), .ZN(new_n619));
  INV_X1    g418(.A(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n612), .A2(new_n616), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT96), .B(KEYINPUT10), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n611), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT10), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(KEYINPUT97), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n629));
  INV_X1    g428(.A(new_n624), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n612), .B2(new_n616), .ZN(new_n631));
  INV_X1    g430(.A(new_n627), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n622), .B1(new_n634), .B2(new_n613), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n625), .A2(new_n627), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n613), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n621), .B1(new_n637), .B2(new_n617), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n608), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n631), .A2(new_n632), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n617), .B1(new_n640), .B2(new_n614), .ZN(new_n641));
  INV_X1    g440(.A(new_n621), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n614), .B1(new_n628), .B2(new_n633), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n643), .B(KEYINPUT98), .C1(new_n644), .C2(new_n622), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AND4_X1   g446(.A1(new_n547), .A2(new_n574), .A3(new_n607), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n535), .B(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g450(.A1(new_n648), .A2(new_n352), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT16), .B(G8gat), .Z(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n655), .B(new_n656), .C1(new_n242), .C2(new_n652), .ZN(G1325gat));
  AOI21_X1  g456(.A(G15gat), .B1(new_n648), .B2(new_n507), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  INV_X1    g458(.A(new_n520), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n660), .A2(G15gat), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n648), .B2(new_n661), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n648), .A2(new_n521), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n516), .A2(new_n546), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n573), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n573), .A2(new_n668), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n513), .B2(new_n458), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n426), .A2(KEYINPUT105), .A3(new_n521), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n520), .A2(new_n673), .A3(new_n545), .A4(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n516), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n677), .A2(new_n273), .A3(new_n607), .A4(new_n646), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n649), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G29gat), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n647), .A2(new_n573), .A3(new_n606), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n649), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(G29gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n547), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT104), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n680), .A2(new_n689), .A3(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(G36gat), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n683), .A2(new_n547), .A3(new_n692), .A4(new_n352), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT46), .Z(new_n694));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n352), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n696), .B2(new_n692), .ZN(G1329gat));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n660), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G43gat), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n547), .A3(new_n216), .A4(new_n507), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1330gat));
  NAND2_X1  g504(.A1(new_n678), .A2(new_n521), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n217), .A2(KEYINPUT106), .ZN(new_n707));
  NOR4_X1   g506(.A1(new_n682), .A2(KEYINPUT106), .A3(G50gat), .A4(new_n458), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n706), .A2(new_n707), .B1(new_n547), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g509(.A1(new_n574), .A2(new_n607), .A3(new_n273), .A4(new_n646), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n516), .B2(new_n675), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n649), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n577), .ZN(G1332gat));
  XNOR2_X1  g513(.A(new_n352), .B(KEYINPUT107), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  XNOR2_X1  g520(.A(new_n507), .B(KEYINPUT108), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(G71gat), .B1(new_n712), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n660), .A2(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n712), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT109), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n521), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g529(.A1(new_n516), .A2(new_n675), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n607), .A2(new_n272), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n574), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n734), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n647), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n418), .A3(new_n649), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n733), .A2(new_n647), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n670), .B2(new_n676), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n649), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n745), .B2(new_n418), .ZN(G1336gat));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n737), .A2(new_n738), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n647), .A2(new_n715), .A3(G92gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT111), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n716), .B(new_n741), .C1(new_n670), .C2(new_n676), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n753), .B1(new_n752), .B2(new_n755), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n352), .B(new_n741), .C1(new_n670), .C2(new_n676), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G92gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n761), .A2(new_n762), .B1(new_n749), .B2(new_n751), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(KEYINPUT110), .A3(G92gat), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n759), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n747), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n752), .A2(new_n755), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n749), .A2(new_n751), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n772), .A3(new_n764), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n774), .A3(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n766), .A2(new_n775), .ZN(G1337gat));
  INV_X1    g575(.A(G99gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n739), .A2(new_n777), .A3(new_n507), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n742), .B2(new_n520), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n742), .A2(new_n779), .A3(new_n520), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n778), .B1(new_n781), .B2(new_n782), .ZN(G1338gat));
  INV_X1    g582(.A(G106gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n739), .A2(new_n784), .A3(new_n521), .ZN(new_n785));
  OAI21_X1  g584(.A(G106gat), .B1(new_n742), .B2(new_n458), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT53), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n787), .A2(KEYINPUT53), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n789), .B(new_n790), .Z(G1339gat));
  NOR4_X1   g590(.A1(new_n646), .A2(new_n573), .A3(new_n606), .A4(new_n272), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n613), .C1(new_n631), .C2(new_n632), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n642), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT97), .B1(new_n625), .B2(new_n627), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n631), .A2(new_n629), .A3(new_n632), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n613), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n640), .B2(new_n614), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n272), .B1(new_n800), .B2(KEYINPUT55), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n794), .A2(new_n642), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT54), .B1(new_n636), .B2(new_n613), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n644), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n804), .A2(new_n805), .B1(new_n644), .B2(new_n622), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n259), .A2(new_n260), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n248), .B1(new_n245), .B2(new_n247), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n207), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT117), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n210), .A2(new_n265), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n639), .B2(new_n645), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n574), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n635), .B1(new_n800), .B2(KEYINPUT55), .ZN(new_n816));
  INV_X1    g615(.A(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n804), .A2(new_n805), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n573), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n792), .B1(new_n820), .B2(new_n606), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n684), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n458), .A2(new_n491), .A3(new_n500), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n716), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n272), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n649), .A2(new_n715), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n521), .B(new_n827), .C1(new_n506), .C2(new_n503), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n646), .A2(new_n817), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n804), .A2(new_n805), .B1(new_n267), .B2(new_n271), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n816), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n573), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n819), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n606), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n792), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n828), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n368), .A3(new_n273), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n826), .A2(new_n839), .ZN(G1340gat));
  AOI21_X1  g639(.A(new_n369), .B1(new_n837), .B2(new_n646), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT118), .Z(new_n842));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n369), .A3(new_n646), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1341gat));
  INV_X1    g643(.A(G127gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n825), .A2(new_n845), .A3(new_n607), .ZN(new_n846));
  OAI21_X1  g645(.A(G127gat), .B1(new_n838), .B2(new_n606), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1342gat));
  NOR4_X1   g647(.A1(new_n824), .A2(G134gat), .A3(new_n352), .A4(new_n574), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n838), .B2(new_n574), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n646), .A2(new_n817), .B1(new_n816), .B2(new_n830), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n573), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT120), .B(new_n574), .C1(new_n807), .C2(new_n814), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n819), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n792), .B1(new_n859), .B2(new_n606), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n458), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT121), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n833), .B1(new_n815), .B2(new_n855), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n607), .B1(new_n866), .B2(new_n858), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n865), .B(new_n862), .C1(new_n867), .C2(new_n792), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n458), .B1(new_n834), .B2(new_n835), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n861), .C1(new_n821), .C2(new_n458), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n864), .A2(new_n868), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n827), .A2(new_n660), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n272), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G141gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n660), .A2(new_n458), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n822), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n716), .ZN(new_n879));
  INV_X1    g678(.A(G141gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n272), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n876), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n874), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n647), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n869), .B(KEYINPUT57), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(new_n646), .A3(new_n874), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT59), .B1(new_n892), .B2(new_n887), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n887), .A3(new_n646), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n889), .B2(new_n606), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n879), .A2(new_n357), .A3(new_n607), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n889), .B2(new_n574), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n573), .A2(new_n358), .A3(new_n353), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n878), .B2(new_n901), .ZN(G1347gat));
  NAND3_X1  g701(.A1(new_n684), .A2(KEYINPUT122), .A3(new_n352), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n649), .B2(new_n353), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR4_X1   g705(.A1(new_n821), .A2(new_n906), .A3(new_n521), .A4(new_n722), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(G169gat), .A3(new_n272), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n836), .A2(new_n823), .A3(new_n684), .A4(new_n716), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n273), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(G169gat), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT123), .Z(G1348gat));
  INV_X1    g711(.A(new_n907), .ZN(new_n913));
  OAI21_X1  g712(.A(G176gat), .B1(new_n913), .B2(new_n647), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n647), .A2(G176gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n909), .B2(new_n915), .ZN(G1349gat));
  INV_X1    g715(.A(new_n295), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n909), .A2(new_n917), .A3(new_n606), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(new_n919));
  OAI21_X1  g718(.A(G183gat), .B1(new_n913), .B2(new_n606), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g721(.A1(new_n909), .A2(G190gat), .A3(new_n574), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT125), .Z(new_n924));
  OAI21_X1  g723(.A(G190gat), .B1(new_n913), .B2(new_n574), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  AND3_X1   g727(.A1(new_n877), .A2(KEYINPUT126), .A3(new_n716), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT126), .B1(new_n877), .B2(new_n716), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n821), .A4(new_n649), .ZN(new_n931));
  AOI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n272), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n903), .A2(new_n520), .A3(new_n905), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT127), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n891), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n272), .A2(G197gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n620), .A3(new_n646), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  AND3_X1   g738(.A1(new_n891), .A2(new_n646), .A3(new_n934), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n620), .B2(new_n940), .ZN(G1353gat));
  NAND3_X1  g740(.A1(new_n931), .A2(new_n275), .A3(new_n607), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n935), .A2(new_n607), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  AOI21_X1  g745(.A(G218gat), .B1(new_n931), .B2(new_n573), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n574), .A2(new_n276), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n935), .B2(new_n948), .ZN(G1355gat));
endmodule


