//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n217), .A2(new_n209), .B1(KEYINPUT65), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n206), .A2(G50), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n212), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G68), .Z(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  OAI21_X1  g0044(.A(KEYINPUT67), .B1(new_n209), .B2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT67), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n246), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n245), .A2(new_n222), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n245), .A2(KEYINPUT68), .A3(new_n222), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G50), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(G13), .ZN(new_n259));
  OR3_X1    g0059(.A1(KEYINPUT69), .A2(G20), .A3(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT69), .B1(G20), .B2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n244), .A2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(G150), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n258), .B1(G50), .B2(new_n259), .C1(new_n252), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  OAI221_X1 g0075(.A(new_n272), .B1(new_n273), .B2(new_n270), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n277), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n285), .B2(G226), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n269), .B(new_n289), .C1(G179), .C2(new_n287), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n269), .B(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n278), .B2(new_n286), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT10), .B1(new_n293), .B2(KEYINPUT71), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n293), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n291), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n291), .B2(new_n297), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n290), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n265), .A2(G77), .ZN(new_n303));
  INV_X1    g0103(.A(new_n261), .ZN(new_n304));
  NOR3_X1   g0104(.A1(KEYINPUT69), .A2(G20), .A3(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G50), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n303), .B1(new_n223), .B2(G68), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n253), .A2(new_n302), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n303), .B1(new_n223), .B2(G68), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(G50), .B2(new_n262), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT73), .B1(new_n311), .B2(new_n252), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n312), .A3(KEYINPUT11), .ZN(new_n316));
  INV_X1    g0116(.A(new_n248), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n255), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n203), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n321), .B2(new_n320), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n319), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n315), .A2(new_n316), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G33), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n327), .A2(new_n329), .A3(G232), .A4(G1698), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n329), .A3(G226), .A4(new_n271), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G97), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n277), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n281), .B1(new_n285), .B2(G238), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n292), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n340), .A2(KEYINPUT72), .B1(new_n343), .B2(new_n295), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n326), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n334), .A2(new_n338), .A3(new_n335), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n348));
  OAI21_X1  g0148(.A(G169), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(KEYINPUT14), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n343), .A2(new_n354), .A3(G169), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n346), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n349), .A2(KEYINPUT14), .B1(new_n351), .B2(G179), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n345), .B1(new_n360), .B2(new_n326), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n327), .A2(new_n329), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n223), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  AOI211_X1 g0165(.A(new_n365), .B(G20), .C1(new_n327), .C2(new_n329), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G20), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n262), .A2(G159), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(KEYINPUT76), .A3(G20), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n367), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT76), .B1(new_n368), .B2(G20), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n365), .B1(new_n270), .B2(G20), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G68), .B1(G159), .B2(new_n262), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n376), .A2(new_n384), .A3(new_n248), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n327), .A2(new_n329), .A3(G226), .A4(G1698), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n327), .A2(new_n329), .A3(G223), .A4(new_n271), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n277), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G41), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(G1), .A3(G13), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(G232), .A3(new_n279), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n284), .A2(G274), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n390), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n295), .A2(KEYINPUT79), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n295), .A2(KEYINPUT79), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g0203(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n292), .B1(new_n406), .B2(new_n390), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G13), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n255), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n264), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n257), .B2(new_n263), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT80), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n385), .A2(new_n408), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT17), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n288), .B1(new_n406), .B2(new_n390), .ZN(new_n417));
  AND4_X1   g0217(.A1(G179), .A2(new_n390), .A3(new_n396), .A4(new_n398), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT78), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n399), .A2(G169), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT78), .ZN(new_n421));
  INV_X1    g0221(.A(G179), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(new_n422), .C2(new_n399), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n385), .A2(new_n413), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  INV_X1    g0232(.A(G238), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n431), .B1(new_n432), .B2(new_n270), .C1(new_n274), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n277), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n281), .B1(new_n285), .B2(G244), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G179), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n288), .B2(new_n437), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n306), .A2(new_n263), .B1(new_n223), .B2(new_n273), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT70), .ZN(new_n441));
  XOR2_X1   g0241(.A(KEYINPUT15), .B(G87), .Z(new_n442));
  AOI22_X1  g0242(.A1(new_n440), .A2(new_n441), .B1(new_n265), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n441), .B2(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n248), .ZN(new_n445));
  MUX2_X1   g0245(.A(new_n259), .B(new_n318), .S(G77), .Z(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n437), .A2(G200), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n435), .A2(G190), .A3(new_n436), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(new_n445), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n301), .A2(new_n362), .A3(new_n430), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n259), .B1(G1), .B2(new_n244), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n250), .B2(new_n251), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G87), .ZN(new_n457));
  OAI21_X1  g0257(.A(G250), .B1(new_n283), .B2(G1), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n254), .A2(G45), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n277), .A2(new_n458), .B1(new_n280), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n327), .A2(new_n329), .A3(G244), .A4(G1698), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n327), .A2(new_n329), .A3(G238), .A4(new_n271), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G116), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n460), .B1(new_n464), .B2(new_n277), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n292), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(G190), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n259), .A2(new_n442), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT82), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G97), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n265), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT19), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n474), .ZN(new_n478));
  NAND3_X1  g0278(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n223), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT82), .B(G97), .ZN(new_n481));
  INV_X1    g0281(.A(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n432), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n327), .A2(new_n329), .A3(new_n223), .A4(G68), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n477), .A2(new_n478), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  AOI211_X1 g0286(.A(KEYINPUT86), .B(new_n468), .C1(new_n486), .C2(new_n248), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT86), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT19), .B1(new_n481), .B2(new_n265), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n484), .B(new_n485), .C1(new_n489), .C2(KEYINPUT85), .ZN(new_n490));
  INV_X1    g0290(.A(new_n478), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n248), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n468), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n457), .B(new_n467), .C1(new_n487), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n270), .A2(G250), .A3(new_n271), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n497));
  INV_X1    g0297(.A(G294), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(new_n244), .C2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n254), .B(G45), .C1(new_n282), .C2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G41), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n277), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n499), .A2(new_n277), .B1(new_n504), .B2(G264), .ZN(new_n505));
  INV_X1    g0305(.A(new_n502), .ZN(new_n506));
  INV_X1    g0306(.A(new_n459), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(G41), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(G274), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G200), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n327), .A2(new_n329), .A3(new_n223), .A4(G87), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n270), .A2(new_n515), .A3(new_n223), .A4(G87), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n463), .B2(G20), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n223), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n223), .B2(G107), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n432), .A2(KEYINPUT23), .A3(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n512), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n514), .B2(new_n516), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT24), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n529), .A3(new_n248), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n254), .A2(new_n432), .A3(G13), .A4(G20), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n533));
  XOR2_X1   g0333(.A(KEYINPUT88), .B(KEYINPUT25), .Z(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n534), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT89), .A3(new_n531), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n456), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n505), .A2(G190), .A3(new_n509), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n511), .A2(new_n530), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n456), .A2(new_n442), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n483), .B1(new_n470), .B2(new_n472), .ZN(new_n543));
  INV_X1    g0343(.A(new_n480), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n485), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT85), .B1(new_n473), .B2(new_n474), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n317), .B1(new_n547), .B2(new_n478), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT86), .B1(new_n548), .B2(new_n468), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n492), .A2(new_n488), .A3(new_n493), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n465), .A2(G169), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n422), .B2(new_n465), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n495), .B(new_n541), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n456), .A2(G97), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n259), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n470), .A2(new_n472), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT83), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n481), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n223), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n306), .B2(new_n273), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n262), .A2(KEYINPUT81), .A3(G77), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n432), .B1(new_n380), .B2(new_n381), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n556), .B(new_n558), .C1(new_n571), .C2(new_n317), .ZN(new_n572));
  OAI211_X1 g0372(.A(G257), .B(new_n392), .C1(new_n500), .C2(new_n502), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n509), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n327), .A2(new_n329), .A3(G244), .A4(new_n271), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n270), .A2(G250), .A3(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(new_n583), .A3(new_n277), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n582), .B2(new_n277), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n422), .B(new_n575), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n574), .B1(new_n582), .B2(new_n277), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G169), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n572), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n559), .A2(new_n560), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n562), .A2(new_n561), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n564), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n382), .A2(G107), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n567), .A4(new_n568), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n248), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n587), .A2(G190), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(new_n556), .A3(new_n558), .A4(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n590), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n555), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n510), .A2(G169), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n505), .A2(G179), .A3(new_n509), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT90), .ZN(new_n609));
  INV_X1    g0409(.A(new_n529), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n248), .B1(new_n528), .B2(KEYINPUT24), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n539), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n609), .B1(new_n530), .B2(new_n539), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n608), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  OAI21_X1  g0416(.A(G116), .B1(new_n244), .B2(G1), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n410), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n317), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n410), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n470), .A2(new_n472), .A3(new_n244), .ZN(new_n623));
  AOI21_X1  g0423(.A(G20), .B1(G33), .B2(G283), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(G20), .B2(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n248), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(KEYINPUT20), .A3(new_n248), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n622), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n327), .A2(new_n329), .A3(G257), .A4(new_n271), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n327), .A2(new_n329), .A3(G264), .A4(G1698), .ZN(new_n632));
  INV_X1    g0432(.A(G303), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n270), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n277), .ZN(new_n635));
  OAI211_X1 g0435(.A(G270), .B(new_n392), .C1(new_n500), .C2(new_n502), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n509), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G169), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n616), .B1(new_n630), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n629), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT20), .B1(new_n625), .B2(new_n248), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n621), .B(new_n619), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n288), .B1(new_n635), .B2(new_n637), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(KEYINPUT21), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n638), .A2(new_n422), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n640), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n638), .A2(G200), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n630), .B(new_n649), .C1(new_n402), .C2(new_n638), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n615), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n454), .A2(new_n605), .A3(new_n651), .ZN(G372));
  AND3_X1   g0452(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n355), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT75), .B1(new_n358), .B2(new_n355), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n326), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n345), .B2(new_n448), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n416), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n417), .A2(new_n418), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n425), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n428), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n425), .A2(KEYINPUT18), .A3(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n657), .A2(new_n664), .B1(new_n299), .B2(new_n300), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(new_n290), .ZN(new_n666));
  INV_X1    g0466(.A(new_n602), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n557), .B1(new_n599), .B2(new_n248), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n588), .B1(new_n668), .B2(new_n556), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n667), .A2(new_n592), .B1(new_n669), .B2(new_n586), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n549), .A2(new_n550), .B1(G87), .B2(new_n456), .ZN(new_n671));
  INV_X1    g0471(.A(new_n542), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n487), .B2(new_n494), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n671), .A2(new_n467), .B1(new_n673), .B2(new_n553), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n530), .A2(new_n539), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n608), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n648), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n670), .A2(new_n674), .A3(new_n541), .A4(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n495), .B1(new_n551), .B2(new_n554), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT26), .B1(new_n679), .B2(new_n590), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n572), .A2(new_n586), .A3(new_n589), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n553), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .A4(new_n495), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n551), .B2(new_n554), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n673), .A2(KEYINPUT91), .A3(new_n553), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n678), .A2(new_n680), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n666), .B1(new_n454), .B2(new_n690), .ZN(G369));
  NAND2_X1  g0491(.A1(new_n648), .A2(new_n650), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n409), .A2(G20), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n254), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n692), .B1(new_n630), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n648), .A2(new_n643), .A3(new_n699), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G330), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n675), .A2(KEYINPUT90), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n705), .A2(new_n612), .B1(new_n606), .B2(new_n607), .ZN(new_n706));
  INV_X1    g0506(.A(new_n541), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n699), .B1(new_n613), .B2(new_n614), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n640), .A2(new_n645), .A3(new_n647), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n700), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n699), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n704), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n712), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n606), .A2(new_n607), .B1(new_n530), .B2(new_n539), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n708), .A2(new_n716), .B1(new_n717), .B2(new_n700), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(G399));
  NAND2_X1  g0519(.A1(new_n543), .A2(new_n620), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n210), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(G1), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n225), .B2(new_n724), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n706), .A2(new_n711), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n604), .A2(new_n728), .A3(new_n650), .A4(new_n700), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n465), .A2(G179), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT92), .A3(new_n638), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT92), .B1(new_n730), .B2(new_n638), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n591), .B(new_n510), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(new_n646), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n587), .A2(new_n505), .A3(new_n465), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n505), .A2(new_n465), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n646), .A3(KEYINPUT30), .A4(new_n587), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n740), .B2(new_n699), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n684), .A2(new_n688), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n747), .B(new_n680), .C1(new_n605), .C2(new_n728), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n700), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(KEYINPUT93), .A3(new_n700), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n689), .A2(new_n700), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n746), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n745), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n727), .B1(new_n758), .B2(G1), .ZN(G364));
  AOI21_X1  g0559(.A(new_n222), .B1(G20), .B2(new_n288), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n402), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n223), .A2(new_n422), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G58), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G20), .A3(new_n295), .ZN(new_n768));
  INV_X1    g0568(.A(G159), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT32), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(new_n295), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n223), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n295), .A3(G200), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n273), .B1(new_n774), .B2(new_n432), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n223), .A2(new_n422), .A3(new_n292), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G190), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n363), .B(new_n775), .C1(G68), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n223), .B1(new_n767), .B2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n469), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n482), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n777), .A2(new_n402), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n781), .B(new_n783), .C1(new_n784), .C2(G50), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n766), .A2(new_n771), .A3(new_n779), .A4(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n764), .ZN(new_n787));
  INV_X1    g0587(.A(new_n772), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(G322), .B1(G311), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G283), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n774), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n768), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n270), .B(new_n791), .C1(G329), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n782), .ZN(new_n794));
  INV_X1    g0594(.A(new_n780), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n794), .A2(G303), .B1(new_n795), .B2(G294), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G326), .A2(new_n784), .B1(new_n778), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n789), .A2(new_n793), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n761), .B1(new_n786), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n760), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n270), .A2(new_n210), .ZN(new_n806));
  INV_X1    g0606(.A(G355), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n806), .A2(new_n807), .B1(G116), .B2(new_n210), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT94), .Z(new_n809));
  NOR2_X1   g0609(.A1(new_n722), .A2(new_n270), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n226), .B2(new_n283), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n283), .B2(new_n242), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n805), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n254), .B1(new_n693), .B2(G45), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n723), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n800), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n701), .A2(new_n702), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n803), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n703), .A2(new_n818), .ZN(new_n823));
  INV_X1    g0623(.A(G330), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(new_n820), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  AND3_X1   g0627(.A1(new_n439), .A2(new_n447), .A3(new_n700), .ZN(new_n828));
  INV_X1    g0628(.A(new_n447), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n451), .B1(new_n829), .B2(new_n700), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n448), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n680), .A2(new_n684), .A3(new_n688), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n711), .A2(new_n717), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n555), .A2(new_n603), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n700), .B(new_n831), .C1(new_n832), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n689), .A2(new_n837), .A3(new_n700), .A4(new_n831), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n831), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n754), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n817), .B1(new_n842), .B2(new_n745), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n745), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n760), .A2(new_n801), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n818), .B1(new_n847), .B2(new_n273), .ZN(new_n848));
  INV_X1    g0648(.A(new_n774), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n788), .A2(G116), .B1(new_n849), .B2(G87), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n850), .B1(new_n432), .B2(new_n782), .C1(new_n498), .C2(new_n764), .ZN(new_n851));
  INV_X1    g0651(.A(new_n784), .ZN(new_n852));
  INV_X1    g0652(.A(new_n778), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n852), .A2(new_n633), .B1(new_n853), .B2(new_n790), .ZN(new_n854));
  INV_X1    g0654(.A(G311), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n363), .B1(new_n768), .B2(new_n855), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n851), .A2(new_n854), .A3(new_n781), .A4(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n784), .A2(G137), .B1(new_n788), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G150), .ZN(new_n859));
  INV_X1    g0659(.A(new_n765), .ZN(new_n860));
  INV_X1    g0660(.A(G143), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n858), .B1(new_n859), .B2(new_n853), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT34), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n363), .B1(new_n792), .B2(G132), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n202), .B2(new_n780), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n307), .A2(new_n782), .B1(new_n774), .B2(new_n203), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT98), .Z(new_n868));
  AOI21_X1  g0668(.A(new_n857), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n848), .B1(new_n831), .B2(new_n802), .C1(new_n761), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n844), .A2(new_n870), .ZN(G384));
  OAI21_X1  g0671(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n225), .A2(new_n872), .B1(G50), .B2(new_n203), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(G1), .A3(new_n409), .ZN(new_n874));
  OAI211_X1 g0674(.A(G116), .B(new_n224), .C1(new_n596), .C2(KEYINPUT35), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(KEYINPUT35), .B2(new_n596), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n874), .B1(new_n876), .B2(KEYINPUT36), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(KEYINPUT36), .B2(new_n876), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n697), .B(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n663), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n385), .A2(new_n408), .A3(new_n413), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n425), .A2(new_n880), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n884), .A2(new_n426), .A3(KEYINPUT103), .A4(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n419), .A2(new_n423), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(new_n879), .B1(new_n385), .B2(new_n413), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n882), .A2(new_n883), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  INV_X1    g0693(.A(new_n882), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n376), .A2(new_n384), .A3(new_n253), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n658), .B1(new_n895), .B2(new_n413), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n697), .B1(new_n895), .B2(new_n413), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n893), .B1(new_n898), .B2(new_n883), .ZN(new_n899));
  INV_X1    g0699(.A(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n882), .ZN(new_n901));
  OAI211_X1 g0701(.A(KEYINPUT101), .B(KEYINPUT37), .C1(new_n901), .C2(new_n896), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n892), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n430), .A2(new_n897), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n660), .A2(new_n885), .A3(new_n882), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n886), .A2(new_n891), .B1(KEYINPUT37), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n885), .B1(new_n416), .B2(new_n663), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n911), .A2(KEYINPUT39), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n904), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n906), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n905), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT39), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n655), .A2(new_n699), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n881), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n345), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n326), .A2(new_n699), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n655), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n360), .A2(new_n326), .A3(new_n699), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n828), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT100), .B1(new_n839), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT100), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n927), .B(new_n828), .C1(new_n836), .C2(new_n838), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n915), .B(new_n924), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n919), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n752), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT93), .B1(new_n748), .B2(new_n700), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT29), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n453), .A3(new_n755), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n666), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n930), .B(new_n935), .Z(new_n936));
  NOR4_X1   g0736(.A1(new_n651), .A2(new_n555), .A3(new_n603), .A4(new_n699), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n740), .A2(new_n699), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT31), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n831), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n326), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n944), .B(new_n700), .C1(new_n357), .C2(new_n359), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n361), .B2(new_n921), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT104), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n744), .A2(new_n924), .A3(new_n831), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n911), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n949), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n950), .A2(KEYINPUT40), .B1(new_n915), .B2(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n454), .B(new_n952), .C1(new_n729), .C2(new_n743), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n744), .A2(new_n924), .A3(new_n831), .ZN(new_n955));
  AOI22_X1  g0755(.A1(KEYINPUT104), .A2(new_n955), .B1(new_n905), .B2(new_n910), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n956), .B2(new_n949), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n949), .B1(new_n914), .B2(new_n905), .ZN(new_n958));
  OAI21_X1  g0758(.A(G330), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n745), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n453), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n953), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n936), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n254), .B2(new_n693), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n964), .A2(KEYINPUT105), .B1(new_n936), .B2(new_n962), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n964), .A2(KEYINPUT105), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n878), .B1(new_n965), .B2(new_n966), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n572), .A2(new_n699), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n590), .B(new_n968), .C1(new_n593), .C2(new_n602), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n681), .A2(new_n699), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT106), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n969), .A2(new_n970), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT106), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n706), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n590), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n700), .ZN(new_n978));
  XOR2_X1   g0778(.A(KEYINPUT107), .B(KEYINPUT42), .Z(new_n979));
  AND4_X1   g0779(.A1(new_n716), .A2(new_n974), .A3(new_n708), .A4(new_n979), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n706), .A2(new_n712), .A3(new_n707), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n979), .B1(new_n981), .B2(new_n974), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n671), .A2(new_n700), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n679), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n686), .A2(new_n985), .A3(new_n687), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n978), .A2(new_n983), .A3(new_n984), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n984), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n699), .B1(new_n976), .B2(new_n590), .ZN(new_n993));
  INV_X1    g0793(.A(new_n983), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n973), .A2(new_n975), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n715), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n990), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n990), .B2(new_n995), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(KEYINPUT108), .B(new_n997), .C1(new_n990), .C2(new_n995), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n708), .A2(new_n716), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n717), .A2(new_n700), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1004), .B1(new_n1007), .B2(new_n971), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(KEYINPUT44), .A3(new_n971), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n718), .B2(new_n974), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(new_n715), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n710), .A2(new_n713), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n703), .A3(new_n712), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1017), .A2(new_n715), .A3(new_n1005), .ZN(new_n1018));
  AOI221_X4 g0818(.A(new_n960), .B1(new_n1015), .B2(new_n1018), .C1(new_n933), .C2(new_n755), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n723), .B(KEYINPUT41), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n815), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1003), .A2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n235), .A2(new_n810), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n442), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n804), .B1(new_n210), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n817), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n795), .A2(G68), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n202), .B2(new_n782), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n853), .A2(new_n769), .B1(new_n772), .B2(new_n307), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n363), .B1(new_n792), .B2(G137), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n852), .B2(new_n861), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n764), .A2(new_n859), .B1(new_n273), .B2(new_n774), .ZN(new_n1033));
  OR4_X1    g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n782), .A2(new_n620), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n853), .A2(new_n498), .B1(KEYINPUT46), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT46), .B2(new_n1035), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(KEYINPUT109), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n481), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n772), .A2(new_n790), .B1(new_n1040), .B2(new_n774), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n363), .B1(new_n1042), .B2(new_n768), .C1(new_n852), .C2(new_n855), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G107), .C2(new_n795), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1039), .B(new_n1044), .C1(new_n633), .C2(new_n860), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1038), .A2(KEYINPUT109), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1034), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT47), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n761), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1027), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n803), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n988), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1023), .A2(new_n1053), .ZN(G387));
  INV_X1    g0854(.A(new_n231), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n810), .B1(new_n1055), .B2(new_n283), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n721), .B2(new_n806), .ZN(new_n1057));
  AOI21_X1  g0857(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1058));
  OR3_X1    g0858(.A1(new_n263), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT50), .B1(new_n263), .B2(G50), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n721), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1057), .A2(new_n1061), .B1(new_n432), .B2(new_n722), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n817), .B1(new_n1062), .B2(new_n805), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n852), .A2(new_n769), .B1(new_n469), .B2(new_n774), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n853), .A2(new_n263), .B1(new_n273), .B2(new_n782), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n764), .A2(new_n307), .B1(new_n203), .B2(new_n772), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n270), .B1(new_n768), .B2(new_n859), .C1(new_n1025), .C2(new_n780), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT110), .Z(new_n1069));
  AOI21_X1  g0869(.A(new_n270), .B1(new_n792), .B2(G326), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n784), .A2(G322), .B1(new_n788), .B2(G303), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n855), .B2(new_n853), .C1(new_n860), .C2(new_n1042), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT48), .Z(new_n1073));
  OAI22_X1  g0873(.A1(new_n782), .A2(new_n498), .B1(new_n780), .B2(new_n790), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1070), .B1(new_n620), .B2(new_n774), .C1(new_n1075), .C2(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(KEYINPUT49), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1069), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n760), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1016), .A2(new_n803), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1080), .A2(new_n1081), .B1(new_n816), .B2(new_n1018), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n745), .B(new_n1018), .C1(new_n753), .C2(new_n756), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT111), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n723), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n758), .B2(new_n1018), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1084), .B1(new_n1083), .B2(new_n723), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NOR2_X1   g0888(.A1(new_n239), .A2(new_n811), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n805), .B1(new_n722), .B2(new_n481), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n853), .A2(new_n633), .B1(new_n790), .B2(new_n782), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n270), .B1(new_n792), .B2(G322), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n432), .B2(new_n774), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n772), .A2(new_n498), .B1(new_n620), .B2(new_n780), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n852), .A2(new_n1042), .B1(new_n764), .B2(new_n855), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n852), .A2(new_n859), .B1(new_n764), .B2(new_n769), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n853), .A2(new_n307), .B1(new_n273), .B2(new_n780), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n270), .B1(new_n768), .B2(new_n861), .C1(new_n774), .C2(new_n482), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n772), .A2(new_n263), .B1(new_n782), .B2(new_n203), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1096), .A2(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n817), .B1(new_n1089), .B2(new_n1091), .C1(new_n1105), .C2(new_n761), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n996), .B2(new_n803), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n715), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(KEYINPUT112), .A3(new_n1015), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1108), .A2(KEYINPUT112), .A3(new_n1109), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1113), .B2(new_n816), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1083), .A2(new_n1112), .A3(new_n1111), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1010), .A2(new_n715), .A3(new_n1014), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n723), .B1(new_n1083), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(G390));
  NAND3_X1  g0918(.A1(new_n934), .A2(new_n666), .A3(new_n961), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n955), .A2(new_n824), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(KEYINPUT113), .ZN(new_n1121));
  OR3_X1    g0921(.A1(new_n955), .A2(KEYINPUT113), .A3(new_n824), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n946), .B1(new_n745), .B2(new_n840), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n839), .A2(new_n925), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n927), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n839), .A2(KEYINPUT100), .A3(new_n925), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n751), .A2(new_n752), .A3(new_n925), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n830), .A2(new_n448), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1119), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n917), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n946), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n918), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1130), .A2(new_n1131), .A3(new_n924), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n918), .B1(new_n905), .B2(new_n910), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1137), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n924), .B1(new_n926), .B2(new_n928), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n918), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n917), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1143), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n955), .A2(new_n824), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1135), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n918), .B1(new_n1128), .B2(new_n924), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1143), .B(new_n1120), .C1(new_n1152), .C2(new_n917), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1136), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n1134), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1151), .A2(new_n723), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n816), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n817), .B1(new_n846), .B2(new_n264), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n787), .A2(G116), .B1(new_n481), .B2(new_n788), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n270), .B(new_n783), .C1(G294), .C2(new_n792), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G283), .A2(new_n784), .B1(new_n778), .B2(G107), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n849), .A2(G68), .B1(new_n795), .B2(G77), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n787), .A2(G132), .B1(G125), .B2(new_n792), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT54), .B(G143), .Z(new_n1165));
  AOI22_X1  g0965(.A1(new_n784), .A2(G128), .B1(new_n788), .B2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n778), .A2(G137), .B1(G159), .B2(new_n795), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n270), .B1(new_n774), .B2(new_n307), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT114), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n782), .A2(new_n859), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1163), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1158), .B1(new_n1174), .B2(new_n760), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n917), .B2(new_n802), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1157), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1156), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT115), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT115), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1156), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(G378));
  AOI21_X1  g0982(.A(new_n818), .B1(new_n847), .B2(new_n307), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n787), .A2(G128), .B1(G137), .B2(new_n788), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G125), .A2(new_n784), .B1(new_n778), .B2(G132), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n794), .A2(new_n1165), .B1(new_n795), .B2(G150), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n849), .A2(G159), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n774), .A2(new_n202), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n852), .A2(new_n620), .B1(new_n764), .B2(new_n432), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G97), .C2(new_n778), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n363), .A2(new_n282), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G283), .B2(new_n792), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n788), .A2(new_n442), .B1(new_n794), .B2(G77), .ZN(new_n1198));
  AND4_X1   g0998(.A1(new_n1028), .A2(new_n1195), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(KEYINPUT58), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1196), .B(new_n307), .C1(G33), .C2(G41), .ZN(new_n1202));
  AND4_X1   g1002(.A1(new_n1192), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n697), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n269), .A2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n301), .A2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n301), .A2(new_n1207), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1205), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n301), .A2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n301), .A2(new_n1207), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1204), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1183), .B1(new_n761), .B2(new_n1203), .C1(new_n1214), .C2(new_n802), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT116), .Z(new_n1216));
  AND2_X1   g1016(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n952), .B2(new_n824), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1214), .B(G330), .C1(new_n957), .C2(new_n958), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n930), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n919), .A3(new_n1219), .A4(new_n929), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n815), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1216), .A2(new_n1223), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1119), .B(KEYINPUT117), .Z(new_n1225));
  NAND2_X1  g1025(.A1(new_n1155), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n723), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1224), .B1(new_n1230), .B2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n816), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n784), .A2(G294), .B1(G97), .B2(new_n794), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n432), .B2(new_n772), .C1(new_n790), .C2(new_n764), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n363), .B1(new_n768), .B2(new_n633), .C1(new_n774), .C2(new_n273), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n778), .A2(G116), .B1(new_n442), .B2(new_n795), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n765), .A2(G137), .B1(new_n778), .B2(new_n1165), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n784), .A2(G132), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT118), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT119), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n363), .B(new_n1193), .C1(G128), .C2(new_n792), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n782), .A2(new_n769), .B1(new_n780), .B2(new_n307), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G150), .B2(new_n788), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1241), .B1(new_n1246), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(new_n761), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n818), .B(new_n1252), .C1(new_n203), .C2(new_n847), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n946), .A2(new_n801), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1235), .A2(KEYINPUT120), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT120), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n815), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1255), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1129), .A2(new_n1133), .A3(new_n1119), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1135), .A2(new_n1020), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(G381));
  AND2_X1   g1064(.A1(G375), .A2(KEYINPUT121), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(G375), .A2(KEYINPUT121), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1265), .A2(new_n1266), .A3(new_n1178), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n826), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G387), .A2(new_n1268), .A3(G384), .A4(G390), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1261), .A3(new_n1263), .A4(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n698), .A2(G213), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT122), .Z(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1267), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(new_n1274), .A3(G213), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT123), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(G407), .A2(new_n1274), .A3(KEYINPUT123), .A4(G213), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1023), .A2(new_n1053), .A3(G390), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G390), .B1(new_n1023), .B2(new_n1053), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1268), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1285), .B(new_n1280), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT60), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1262), .A2(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1129), .A2(new_n1133), .A3(new_n1119), .A4(KEYINPUT60), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1292), .A2(new_n1135), .A3(new_n723), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT124), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1261), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1295), .A2(KEYINPUT124), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1256), .A2(new_n1260), .B1(new_n1295), .B2(KEYINPUT124), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1298), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1294), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(G2897), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1272), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1299), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1271), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1299), .A2(new_n1302), .B1(G2897), .B2(new_n1307), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  AND4_X1   g1109(.A1(new_n929), .A2(new_n1218), .A3(new_n919), .A4(new_n1219), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1218), .A2(new_n1219), .B1(new_n919), .B2(new_n929), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n816), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1215), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1155), .A2(new_n1225), .B1(new_n1222), .B2(new_n1221), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1313), .B1(new_n1314), .B2(new_n1020), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(new_n1178), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1224), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1226), .A2(new_n1231), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1227), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n724), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1316), .B1(G378), .B2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1309), .B1(new_n1322), .B2(new_n1273), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1229), .B(new_n723), .C1(KEYINPUT57), .C2(new_n1314), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1156), .A2(new_n1180), .A3(new_n1177), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1180), .B1(new_n1156), .B2(new_n1177), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1324), .B(new_n1224), .C1(new_n1325), .C2(new_n1326), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1315), .A2(new_n1178), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1307), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1301), .B1(new_n1300), .B2(new_n1294), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1329), .A2(new_n1333), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1290), .B(new_n1323), .C1(new_n1334), .C2(KEYINPUT62), .ZN(new_n1335));
  AOI211_X1 g1135(.A(new_n1273), .B(new_n1332), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1289), .B1(new_n1335), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1309), .B1(new_n1322), .B2(new_n1307), .ZN(new_n1340));
  AOI22_X1  g1140(.A1(new_n1340), .A2(KEYINPUT63), .B1(new_n1333), .B2(new_n1329), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1342), .A2(KEYINPUT63), .A3(new_n1272), .A4(new_n1333), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1344), .B(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1343), .A2(new_n1346), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1341), .A2(KEYINPUT127), .A3(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT127), .ZN(new_n1349));
  OAI22_X1  g1149(.A1(new_n1330), .A2(new_n1331), .B1(new_n1303), .B2(new_n1271), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1305), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1351), .B1(new_n1342), .B2(new_n1271), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1334), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1344), .B(KEYINPUT126), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1355), .B1(new_n1336), .B2(KEYINPUT63), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1349), .B1(new_n1354), .B2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1339), .B1(new_n1348), .B2(new_n1357), .ZN(G405));
  XOR2_X1   g1158(.A(new_n1332), .B(new_n1289), .Z(new_n1359));
  OAI21_X1  g1159(.A(new_n1327), .B1(new_n1178), .B2(new_n1321), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1359), .B(new_n1360), .ZN(G402));
endmodule


