//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G169gat), .A3(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n214), .B(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT65), .B(G169gat), .Z(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT23), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n207), .A2(new_n209), .B1(KEYINPUT23), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n214), .A2(new_n216), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n218), .A2(new_n219), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n221), .A2(new_n224), .B1(new_n229), .B2(KEYINPUT25), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT68), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n231), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n210), .A2(new_n232), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(G183gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(G183gat), .ZN(new_n243));
  AOI21_X1  g042(.A(G190gat), .B1(new_n243), .B2(KEYINPUT67), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT28), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n238), .A2(KEYINPUT27), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n247), .A2(new_n248), .A3(G190gat), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n217), .B(new_n236), .C1(new_n245), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G120gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n257));
  INV_X1    g056(.A(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G120gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G134gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n230), .A2(new_n250), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n230), .B2(new_n250), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n205), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT32), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT33), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  NAND3_X1  g074(.A1(new_n270), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n275), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n269), .B(KEYINPUT32), .C1(new_n271), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n267), .A2(new_n268), .A3(KEYINPUT34), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n204), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n230), .A2(new_n250), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n257), .A2(new_n265), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT34), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n230), .A2(new_n250), .A3(new_n266), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n204), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n203), .A3(new_n287), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT34), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n282), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n202), .B1(new_n279), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n282), .A2(new_n289), .A3(new_n291), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(KEYINPUT71), .A3(new_n278), .A4(new_n276), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  INV_X1    g097(.A(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G148gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n304), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n303), .A2(new_n307), .B1(new_n310), .B2(new_n301), .ZN(new_n311));
  XNOR2_X1  g110(.A(G197gat), .B(G204gat), .ZN(new_n312));
  INV_X1    g111(.A(G211gat), .ZN(new_n313));
  INV_X1    g112(.A(G218gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(KEYINPUT22), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G211gat), .B(G218gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT73), .B(KEYINPUT29), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n311), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n317), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n316), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n308), .A2(KEYINPUT74), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT2), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n307), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n301), .B1(new_n305), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n322), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OR3_X1    g138(.A1(new_n323), .A2(new_n325), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n318), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n311), .B1(new_n342), .B2(new_n322), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n325), .B1(new_n343), .B2(new_n339), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT31), .B(G50gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT77), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n323), .A2(new_n325), .A3(new_n339), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n322), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n324), .B1(new_n352), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n346), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n356), .B(G22gat), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n348), .A2(new_n354), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n294), .A2(KEYINPUT70), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n292), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n279), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n296), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT83), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n311), .B(new_n284), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT5), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n266), .A2(new_n372), .A3(new_n311), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT4), .B1(new_n351), .B2(new_n284), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT75), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n266), .A2(new_n376), .A3(new_n311), .A4(new_n372), .ZN(new_n377));
  XNOR2_X1  g176(.A(G155gat), .B(G162gat), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n301), .B2(new_n302), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n309), .A2(new_n304), .B1(new_n298), .B2(new_n300), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n284), .A3(new_n336), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(new_n369), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n375), .A2(new_n383), .A3(KEYINPUT76), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n377), .A2(new_n382), .A3(new_n369), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT75), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n371), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT0), .B(G57gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G85gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n374), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(new_n369), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n395), .A2(KEYINPUT5), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n393), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n393), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT76), .B1(new_n375), .B2(new_n383), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n377), .A2(new_n382), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(new_n385), .A3(new_n387), .A4(new_n369), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n370), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n404), .B2(new_n397), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT6), .B(new_n400), .C1(new_n404), .C2(new_n397), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n411), .B1(new_n283), .B2(new_n341), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n410), .B(KEYINPUT72), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n230), .B2(new_n250), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n318), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n283), .A2(new_n411), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n319), .B1(new_n230), .B2(new_n250), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n416), .B(new_n327), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  INV_X1    g220(.A(G64gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G92gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n419), .A3(new_n425), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT30), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n430), .A3(new_n426), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT83), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n296), .A2(new_n434), .A3(new_n361), .A4(new_n365), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n367), .A2(new_n409), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n279), .A2(new_n292), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n296), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n441));
  INV_X1    g240(.A(new_n408), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n407), .B2(KEYINPUT80), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n399), .A2(new_n405), .A3(new_n444), .A4(new_n406), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n441), .B1(new_n446), .B2(new_n433), .ZN(new_n447));
  AOI211_X1 g246(.A(KEYINPUT82), .B(new_n432), .C1(new_n443), .C2(new_n445), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n438), .B(new_n440), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n361), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n437), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n426), .B1(new_n420), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n455), .B2(new_n318), .ZN(new_n456));
  OR3_X1    g255(.A1(new_n412), .A2(new_n318), .A3(new_n414), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT38), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n454), .A2(new_n458), .B1(new_n420), .B2(new_n426), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n452), .A2(new_n408), .A3(new_n445), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT81), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n453), .B2(new_n420), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT38), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT81), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n443), .A2(new_n464), .A3(new_n445), .A4(new_n459), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n369), .B1(new_n394), .B2(new_n382), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT39), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n468), .B1(new_n368), .B2(new_n369), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT79), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n393), .B(new_n469), .C1(new_n471), .C2(new_n467), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n432), .A2(new_n405), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n450), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n466), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT78), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n348), .A2(new_n354), .A3(new_n357), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n357), .B1(new_n348), .B2(new_n354), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n359), .A2(KEYINPUT78), .A3(new_n360), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n409), .B2(new_n433), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n296), .A2(new_n486), .A3(new_n439), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n296), .B2(new_n365), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n478), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n451), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(G43gat), .B(G50gat), .Z(new_n492));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n493));
  INV_X1    g292(.A(G29gat), .ZN(new_n494));
  INV_X1    g293(.A(G36gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n492), .A2(new_n493), .B1(KEYINPUT85), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT14), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n497), .B(new_n499), .C1(KEYINPUT85), .C2(new_n496), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n492), .A2(new_n493), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n509), .B2(new_n508), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G8gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n503), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT13), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n502), .A2(KEYINPUT86), .A3(KEYINPUT17), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT17), .B1(new_n502), .B2(KEYINPUT86), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n503), .A2(new_n512), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n514), .A4(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n522), .A2(new_n523), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(new_n514), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n519), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT12), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n519), .A2(new_n528), .A3(new_n530), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n491), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n491), .A2(KEYINPUT90), .A3(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT9), .B1(new_n550), .B2(KEYINPUT91), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT92), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n548), .B1(new_n547), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n512), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT95), .ZN(new_n564));
  AND2_X1   g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT20), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n561), .A2(new_n562), .ZN(new_n572));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT94), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT19), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n572), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n569), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n571), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n571), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G190gat), .B(G218gat), .Z(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT98), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT8), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT97), .B(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n586), .B(new_n588), .C1(new_n590), .C2(G85gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n584), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n597), .A2(new_n502), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n520), .B2(new_n521), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n582), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT96), .B(G134gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G162gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n604), .B(new_n605), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n600), .A3(new_n582), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n608), .B1(new_n601), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT100), .A4(new_n582), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n610), .B1(new_n614), .B2(new_n606), .ZN(new_n615));
  AOI211_X1 g414(.A(KEYINPUT101), .B(new_n607), .C1(new_n612), .C2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n581), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT105), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G120gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n297), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n554), .A2(new_n560), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n584), .B(KEYINPUT102), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n591), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n594), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n596), .A2(new_n561), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT103), .B(KEYINPUT10), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G230gat), .A2(G233gat), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n624), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  AOI211_X1 g435(.A(KEYINPUT106), .B(new_n636), .C1(new_n631), .C2(new_n632), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n634), .B1(new_n628), .B2(new_n629), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n623), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n631), .A2(new_n642), .A3(new_n632), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n631), .B2(new_n632), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n634), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n645), .A2(new_n640), .A3(new_n623), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n546), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n409), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n509), .ZN(G1324gat));
  NOR2_X1   g450(.A1(new_n649), .A2(new_n433), .ZN(new_n652));
  NAND2_X1  g451(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n653));
  INV_X1    g452(.A(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n505), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n658), .B(new_n659), .C1(new_n654), .C2(new_n652), .ZN(G1325gat));
  NOR2_X1   g459(.A1(new_n487), .A2(new_n488), .ZN(new_n661));
  OAI21_X1  g460(.A(G15gat), .B1(new_n649), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(G15gat), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n546), .A2(new_n663), .A3(new_n440), .A4(new_n648), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT107), .Z(G1326gat));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n484), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  XNOR2_X1  g468(.A(new_n647), .B(KEYINPUT109), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n541), .A3(new_n580), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n490), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n478), .A2(KEYINPUT110), .A3(new_n489), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n451), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n617), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT111), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n676), .A2(KEYINPUT111), .A3(new_n677), .A4(new_n617), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n677), .B1(new_n491), .B2(new_n617), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n672), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n409), .ZN(new_n687));
  INV_X1    g486(.A(new_n647), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n580), .A2(new_n617), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT108), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n544), .B2(new_n545), .ZN(new_n691));
  INV_X1    g490(.A(new_n409), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n494), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n687), .A2(new_n694), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n432), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(G36gat), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n691), .A2(KEYINPUT112), .A3(new_n495), .A4(new_n432), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(KEYINPUT113), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(G36gat), .B1(new_n686), .B2(new_n433), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n702), .B(new_n703), .C1(new_n700), .C2(new_n704), .ZN(G1329gat));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n706));
  INV_X1    g505(.A(new_n661), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n685), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n683), .B1(new_n680), .B2(new_n681), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n709), .A2(KEYINPUT114), .A3(new_n661), .A4(new_n672), .ZN(new_n710));
  INV_X1    g509(.A(G43gat), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n440), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT47), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(G43gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n685), .A2(new_n707), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  OAI22_X1  g516(.A1(new_n712), .A2(new_n714), .B1(new_n717), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g517(.A(G50gat), .B1(new_n686), .B2(new_n361), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n484), .A2(G50gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT115), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n691), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(KEYINPUT48), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n484), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n685), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n725), .A2(G50gat), .B1(new_n691), .B2(new_n721), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n676), .A2(new_n670), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n619), .A2(new_n541), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n692), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n432), .B1(new_n734), .B2(new_n422), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT116), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n422), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n731), .A2(new_n740), .A3(new_n440), .ZN(new_n741));
  OAI21_X1  g540(.A(G71gat), .B1(new_n730), .B2(new_n661), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g543(.A1(new_n730), .A2(new_n484), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT117), .B(G78gat), .Z(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1335gat));
  INV_X1    g546(.A(new_n541), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n580), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n688), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n682), .B2(new_n684), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n409), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n676), .A2(new_n617), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  OR3_X1    g555(.A1(new_n755), .A2(new_n756), .A3(new_n749), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n749), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n688), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n760), .A3(new_n692), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n761), .ZN(G1336gat));
  NAND2_X1  g561(.A1(new_n682), .A2(new_n684), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n432), .A3(new_n750), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n590), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n757), .A2(new_n758), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n433), .A2(G92gat), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n670), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n765), .A2(KEYINPUT118), .A3(KEYINPUT52), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g568(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n770));
  NAND2_X1  g569(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n589), .B1(new_n752), .B2(new_n432), .ZN(new_n772));
  INV_X1    g571(.A(new_n767), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n671), .B(new_n773), .C1(new_n757), .C2(new_n758), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n769), .A2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n753), .B2(new_n661), .ZN(new_n777));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n778), .A3(new_n440), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1338gat));
  AOI211_X1 g579(.A(G106gat), .B(new_n671), .C1(new_n757), .C2(new_n758), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n781), .B2(new_n450), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT119), .B(G106gat), .Z(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n753), .B2(new_n361), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n752), .A2(new_n724), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n787), .A2(new_n783), .B1(new_n781), .B2(new_n450), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n631), .A2(new_n636), .A3(new_n632), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n645), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n623), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n635), .B2(new_n637), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n792), .A4(new_n794), .ZN(new_n798));
  INV_X1    g597(.A(new_n646), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n797), .A2(new_n541), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n529), .A2(new_n514), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n513), .A2(new_n516), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n536), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n540), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n647), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n617), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n797), .A2(new_n799), .A3(new_n798), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n617), .A2(new_n804), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n580), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n581), .A2(new_n618), .A3(new_n748), .A4(new_n688), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n367), .A2(new_n435), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n409), .A2(new_n432), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n260), .A3(new_n541), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n812), .A2(new_n440), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n484), .A3(new_n814), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n819), .A2(KEYINPUT120), .A3(new_n484), .A4(new_n814), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n541), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n825), .B2(new_n260), .ZN(G1340gat));
  NAND4_X1  g625(.A1(new_n822), .A2(G120gat), .A3(new_n670), .A4(new_n823), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n258), .B1(new_n816), .B2(new_n688), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n827), .A2(KEYINPUT121), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n817), .B2(new_n581), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n580), .A2(new_n253), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n824), .B2(new_n835), .ZN(G1342gat));
  NOR3_X1   g635(.A1(new_n816), .A2(G134gat), .A3(new_n618), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT56), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n824), .A2(new_n617), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n251), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n661), .A2(new_n814), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n361), .B1(new_n810), .B2(new_n811), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n806), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT122), .B(new_n617), .C1(new_n800), .C2(new_n805), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n809), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n581), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n811), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n724), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n845), .B1(new_n853), .B2(KEYINPUT57), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n299), .B1(new_n854), .B2(new_n541), .ZN(new_n855));
  INV_X1    g654(.A(new_n841), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n842), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(G141gat), .A3(new_n748), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT58), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n806), .A2(new_n846), .ZN(new_n860));
  INV_X1    g659(.A(new_n848), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n850), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n580), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n484), .B1(new_n863), .B2(new_n811), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n844), .B1(new_n864), .B2(new_n843), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n748), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867));
  INV_X1    g666(.A(new_n858), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n859), .A2(new_n869), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n812), .A2(new_n450), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n484), .A2(KEYINPUT57), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n871), .A2(KEYINPUT57), .B1(new_n812), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(new_n647), .A3(new_n856), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n874), .B2(new_n297), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n865), .B2(new_n688), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n297), .ZN(new_n878));
  INV_X1    g677(.A(new_n857), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n297), .A3(new_n647), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1345gat));
  AOI21_X1  g680(.A(G155gat), .B1(new_n879), .B2(new_n581), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n865), .A2(new_n580), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g683(.A(G162gat), .B1(new_n879), .B2(new_n617), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n618), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(G162gat), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n813), .A2(new_n432), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n692), .B1(new_n888), .B2(KEYINPUT123), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n812), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n222), .A3(new_n541), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT124), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n692), .A2(new_n433), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n819), .A2(new_n484), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n748), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n892), .B2(new_n647), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n896), .A2(new_n223), .A3(new_n671), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  OAI21_X1  g700(.A(G183gat), .B1(new_n896), .B2(new_n580), .ZN(new_n902));
  INV_X1    g701(.A(new_n247), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n890), .A2(new_n903), .A3(new_n581), .A4(new_n891), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(KEYINPUT125), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT60), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(new_n902), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1350gat));
  INV_X1    g710(.A(G190gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n912), .A3(new_n617), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n896), .A2(new_n618), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G1351gat));
  NAND2_X1  g717(.A1(new_n812), .A2(new_n872), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n661), .A2(new_n895), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n919), .B(new_n921), .C1(new_n843), .C2(new_n842), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT126), .B1(new_n922), .B2(new_n748), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n873), .A2(new_n924), .A3(new_n541), .A4(new_n921), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n925), .A3(G197gat), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n842), .A2(new_n921), .ZN(new_n927));
  OR3_X1    g726(.A1(new_n927), .A2(G197gat), .A3(new_n748), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(KEYINPUT127), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1352gat));
  NOR3_X1   g732(.A1(new_n927), .A2(G204gat), .A3(new_n688), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  OAI21_X1  g734(.A(G204gat), .B1(new_n922), .B2(new_n671), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n873), .A2(new_n581), .A3(new_n921), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n581), .A2(new_n313), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n940), .A2(new_n941), .B1(new_n927), .B2(new_n942), .ZN(G1354gat));
  OAI21_X1  g742(.A(G218gat), .B1(new_n922), .B2(new_n618), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n617), .A2(new_n314), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n927), .B2(new_n945), .ZN(G1355gat));
endmodule


