//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085;
  AND2_X1   g000(.A1(KEYINPUT68), .A2(G953), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT68), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XOR2_X1   g004(.A(G110), .B(G140), .Z(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT65), .B1(new_n196), .B2(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(new_n198), .C1(new_n194), .C2(G137), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n199), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n194), .B2(G137), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n201), .A4(new_n195), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n203), .A2(KEYINPUT66), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(G131), .C1(new_n199), .C2(new_n202), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n208), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT67), .B1(new_n208), .B2(new_n210), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n214));
  XNOR2_X1  g028(.A(G104), .B(G107), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT76), .B(G101), .ZN(new_n218));
  INV_X1    g032(.A(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(new_n219), .B2(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(G107), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G104), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n218), .A2(new_n220), .A3(new_n221), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(G104), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n221), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT77), .A3(G101), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n217), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT10), .ZN(new_n230));
  INV_X1    g044(.A(G143), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n231), .B2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(G146), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  OAI211_X1 g049(.A(G128), .B(new_n232), .C1(new_n233), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(G143), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(G146), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(new_n238), .C1(KEYINPUT1), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n229), .A2(new_n230), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n217), .A2(new_n225), .A3(new_n228), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT10), .B1(new_n244), .B2(new_n241), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n220), .A2(new_n224), .A3(new_n221), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G101), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT75), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n247), .A2(new_n250), .A3(G101), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n225), .A4(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(new_n253), .A3(G101), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT0), .A3(G128), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT0), .B(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n246), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n193), .B1(new_n213), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n196), .A2(G134), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n204), .B2(KEYINPUT11), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n206), .B1(new_n267), .B2(new_n201), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n210), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n208), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n243), .A2(new_n245), .B1(new_n252), .B2(new_n260), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n263), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n229), .A2(new_n242), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n244), .A2(new_n241), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT12), .B1(new_n213), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n278), .B2(new_n279), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n269), .A2(new_n270), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n276), .B1(new_n286), .B2(new_n192), .ZN(new_n287));
  OAI21_X1  g101(.A(G469), .B1(new_n287), .B2(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n271), .A2(new_n280), .A3(new_n272), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n289), .A2(new_n282), .B1(new_n284), .B2(new_n283), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT78), .B1(new_n290), .B2(new_n263), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n192), .B1(new_n273), .B2(new_n274), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n293), .C1(new_n281), .C2(new_n285), .ZN(new_n294));
  INV_X1    g108(.A(new_n277), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n192), .B1(new_n295), .B2(new_n275), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  OAI21_X1  g116(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G110), .B(G122), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G116), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G113), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n317), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n254), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n249), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n311), .A2(G119), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n314), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT5), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n328), .A2(new_n329), .B1(new_n320), .B2(new_n319), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n225), .A3(new_n228), .A4(new_n217), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n308), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n249), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n251), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n307), .C1(new_n336), .C2(new_n323), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n259), .A2(G125), .ZN(new_n339));
  INV_X1    g153(.A(G125), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT79), .B1(new_n241), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n342), .B(G125), .C1(new_n236), .C2(new_n240), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G953), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G224), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n344), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n308), .C1(new_n325), .C2(new_n332), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n338), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n299), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n307), .B(KEYINPUT8), .ZN(new_n353));
  INV_X1    g167(.A(new_n330), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n244), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n331), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT80), .B1(new_n229), .B2(new_n330), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n241), .A2(new_n340), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n342), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n241), .A2(KEYINPUT79), .A3(new_n340), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n339), .A4(new_n346), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n364), .A3(new_n337), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(KEYINPUT81), .A3(new_n362), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n341), .B2(new_n343), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n368), .A3(new_n339), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT7), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n347), .B1(KEYINPUT82), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(KEYINPUT82), .B2(new_n370), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(KEYINPUT83), .A3(new_n372), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n365), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n306), .B1(new_n352), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n359), .A2(new_n364), .A3(new_n337), .ZN(new_n380));
  INV_X1    g194(.A(new_n376), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT83), .B1(new_n369), .B2(new_n372), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(new_n299), .A3(new_n351), .A4(new_n305), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G214), .B1(G237), .B2(G902), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n352), .A2(new_n377), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT84), .A3(new_n305), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n304), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n259), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n271), .A2(new_n391), .A3(new_n272), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n194), .A2(G137), .ZN(new_n393));
  OAI21_X1  g207(.A(G131), .B1(new_n393), .B2(new_n266), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n242), .A2(new_n207), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n322), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n392), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT28), .B1(new_n392), .B2(new_n397), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n189), .A2(G210), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT27), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT26), .B(G101), .Z(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n208), .A2(new_n391), .A3(new_n210), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n395), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n322), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n398), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n416), .A2(new_n402), .A3(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n395), .A2(KEYINPUT30), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n392), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n396), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n420), .A2(new_n422), .B1(new_n392), .B2(new_n397), .ZN(new_n423));
  INV_X1    g237(.A(new_n408), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n409), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n411), .B(new_n299), .C1(new_n417), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G472), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n408), .B1(new_n416), .B2(new_n402), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n408), .B1(new_n392), .B2(new_n397), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n418), .B1(new_n213), .B2(new_n391), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n414), .A2(new_n421), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n322), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT31), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n420), .A2(new_n422), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT69), .B(KEYINPUT31), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n439));
  NOR2_X1   g253(.A1(G472), .A2(G902), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n427), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G137), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n340), .A2(G140), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(KEYINPUT16), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT16), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT71), .B1(new_n448), .B2(KEYINPUT16), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G146), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n234), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n239), .A2(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n309), .A2(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT24), .B(G110), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NOR2_X1   g280(.A1(KEYINPUT70), .A2(KEYINPUT23), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n459), .B(new_n465), .C1(new_n468), .C2(new_n458), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n462), .B1(new_n469), .B2(G110), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n460), .A2(new_n461), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n469), .B2(G110), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n448), .A2(new_n449), .A3(new_n234), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n455), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT72), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n471), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n471), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n446), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n446), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n471), .A2(new_n475), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(KEYINPUT72), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n299), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n479), .A2(new_n299), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G217), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G234), .B2(new_n299), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n491), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n479), .A2(new_n299), .A3(new_n493), .A4(new_n482), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT74), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT20), .ZN(new_n498));
  XNOR2_X1  g312(.A(G113), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n219), .ZN(new_n500));
  OR2_X1    g314(.A1(KEYINPUT68), .A2(G953), .ZN(new_n501));
  NAND2_X1  g315(.A1(KEYINPUT68), .A2(G953), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n501), .A2(G214), .A3(new_n404), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n231), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n189), .A2(G143), .A3(G214), .A4(new_n404), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n206), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT85), .A4(new_n206), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G131), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n448), .A2(new_n449), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT19), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n455), .C1(G146), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(G146), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n474), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT18), .A2(G131), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n504), .B2(new_n505), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n500), .B1(new_n515), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n526), .B(new_n206), .C1(new_n504), .C2(new_n505), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n457), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n508), .A2(new_n511), .A3(new_n526), .A4(new_n509), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT86), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(new_n500), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n530), .B2(new_n500), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n525), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G475), .A2(G902), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n498), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n528), .A2(new_n529), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n500), .A3(new_n523), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n531), .A3(new_n500), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n524), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(KEYINPUT87), .B2(KEYINPUT20), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n540), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n537), .A2(new_n523), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n500), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n530), .A2(KEYINPUT88), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G475), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n536), .A2(new_n546), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G478), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(KEYINPUT92), .B2(KEYINPUT15), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n231), .A2(G128), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n239), .A2(G143), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n194), .ZN(new_n561));
  INV_X1    g375(.A(G122), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G116), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n311), .A2(G122), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(new_n223), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n223), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT13), .B1(new_n231), .B2(G128), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n231), .A2(G128), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n231), .A2(KEYINPUT13), .A3(G128), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n194), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT89), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n311), .A2(G122), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n562), .A2(G116), .ZN(new_n575));
  OAI21_X1  g389(.A(G107), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n563), .A2(new_n564), .A3(new_n223), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n239), .B2(G143), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n571), .A3(new_n560), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G134), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT89), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n578), .A2(new_n582), .A3(new_n583), .A4(new_n561), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n239), .A2(G143), .ZN(new_n585));
  OAI21_X1  g399(.A(G134), .B1(new_n585), .B2(new_n569), .ZN(new_n586));
  XNOR2_X1  g400(.A(G116), .B(G122), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n586), .A2(new_n561), .B1(new_n223), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT14), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n311), .B2(G122), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT90), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n564), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT14), .B1(new_n562), .B2(G116), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n575), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT90), .B1(new_n564), .B2(KEYINPUT14), .ZN(new_n595));
  OAI211_X1 g409(.A(G107), .B(new_n592), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n302), .A2(new_n490), .A3(G953), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n573), .A2(new_n584), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT91), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n578), .A2(new_n582), .A3(new_n561), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n601), .A2(KEYINPUT89), .B1(new_n596), .B2(new_n588), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n602), .A2(new_n603), .A3(new_n584), .A4(new_n598), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n573), .A2(new_n584), .A3(new_n597), .ZN(new_n605));
  INV_X1    g419(.A(new_n598), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n299), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT93), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(KEYINPUT93), .A3(new_n299), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n558), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n558), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n345), .A2(G952), .ZN(new_n617));
  INV_X1    g431(.A(G234), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n404), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n299), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n556), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n390), .A2(new_n443), .A3(new_n497), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(new_n218), .Z(G3));
  INV_X1    g442(.A(G472), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n438), .B2(new_n299), .ZN(new_n630));
  INV_X1    g444(.A(new_n440), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT31), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n435), .B2(new_n429), .ZN(new_n633));
  INV_X1    g447(.A(new_n433), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n436), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n635), .B2(new_n428), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n496), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n386), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n378), .B2(new_n384), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n607), .A2(KEYINPUT33), .A3(new_n599), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n640), .A2(KEYINPUT95), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT94), .B(KEYINPUT33), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n608), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(KEYINPUT95), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G478), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(G902), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n645), .A2(new_n647), .B1(new_n646), .B2(new_n609), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n556), .A2(new_n639), .A3(new_n649), .A4(new_n624), .ZN(new_n650));
  INV_X1    g464(.A(new_n303), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n288), .B2(new_n300), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n637), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  AND2_X1   g469(.A1(new_n639), .A2(new_n624), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n657));
  INV_X1    g471(.A(new_n535), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n541), .A2(KEYINPUT20), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(new_n659), .B2(new_n536), .ZN(new_n660));
  OAI21_X1  g474(.A(KEYINPUT20), .B1(new_n541), .B2(new_n658), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n534), .A2(new_n498), .A3(new_n535), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT96), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  OAI22_X1  g478(.A1(new_n554), .A2(new_n555), .B1(new_n613), .B2(new_n615), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n656), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n630), .A2(new_n636), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n667), .A2(new_n669), .A3(new_n496), .A4(new_n304), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT35), .B(G107), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NOR2_X1   g486(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n481), .B(new_n673), .Z(new_n674));
  NOR3_X1   g488(.A1(new_n674), .A2(G902), .A3(new_n491), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n489), .B2(new_n491), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n390), .A2(new_n626), .A3(new_n668), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT97), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT97), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n683), .A2(new_n619), .A3(new_n684), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n685), .B(new_n665), .C1(new_n660), .C2(new_n663), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n301), .A2(new_n303), .A3(new_n639), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n443), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  AND2_X1   g503(.A1(new_n392), .A2(new_n395), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n398), .B1(new_n690), .B2(new_n396), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n299), .B1(new_n691), .B2(new_n424), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n423), .A2(new_n408), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n441), .B2(new_n442), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n556), .ZN(new_n697));
  INV_X1    g511(.A(new_n558), .ZN(new_n698));
  INV_X1    g512(.A(new_n612), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT93), .B1(new_n608), .B2(new_n299), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n614), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n676), .A2(new_n702), .A3(new_n386), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n696), .A2(new_n697), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n385), .A2(new_n388), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT38), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n685), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n652), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n704), .A2(new_n709), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  INV_X1    g529(.A(new_n685), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n556), .A2(new_n649), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n687), .A2(new_n718), .A3(new_n443), .A4(new_n677), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(new_n297), .A2(new_n299), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(new_n303), .A3(new_n300), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n650), .A2(new_n443), .A3(new_n497), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(KEYINPUT41), .B(G113), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND2_X1  g540(.A1(new_n438), .A2(new_n440), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT32), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n496), .B1(new_n730), .B2(new_n427), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n664), .A2(new_n666), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n733), .A3(new_n656), .A4(new_n723), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT98), .B(G116), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G18));
  AND4_X1   g550(.A1(new_n303), .A2(new_n639), .A3(new_n722), .A4(new_n300), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n443), .A3(new_n626), .A4(new_n677), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  NAND2_X1  g553(.A1(new_n722), .A2(new_n300), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n623), .A3(new_n651), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n378), .A2(new_n384), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n702), .A3(new_n386), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT101), .B1(new_n743), .B2(new_n556), .ZN(new_n744));
  AND4_X1   g558(.A1(KEYINPUT101), .A2(new_n556), .A3(new_n639), .A4(new_n702), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n402), .B1(new_n691), .B2(KEYINPUT28), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT99), .B(new_n434), .C1(new_n747), .C2(new_n424), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT99), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n424), .B1(new_n401), .B2(new_n403), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n749), .B1(new_n750), .B2(new_n633), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n751), .A3(new_n437), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n440), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n630), .A2(KEYINPUT100), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n630), .A2(KEYINPUT100), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n753), .B(new_n497), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n746), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n562), .ZN(G24));
  OAI211_X1 g573(.A(new_n753), .B(new_n677), .C1(new_n755), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n717), .A2(KEYINPUT102), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n534), .A2(new_n544), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n661), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n500), .B1(new_n548), .B2(new_n549), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n552), .A2(new_n764), .B1(new_n539), .B2(new_n540), .ZN(new_n765));
  OAI21_X1  g579(.A(G475), .B1(new_n765), .B2(G902), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n648), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT102), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n716), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n737), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n760), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT103), .B(G125), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G27));
  AOI21_X1  g588(.A(new_n638), .B1(new_n385), .B2(new_n388), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n761), .A2(new_n769), .A3(new_n652), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n443), .A2(new_n497), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n770), .ZN(new_n779));
  INV_X1    g593(.A(new_n775), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n304), .ZN(new_n781));
  OAI21_X1  g595(.A(KEYINPUT104), .B1(new_n441), .B2(new_n442), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n728), .A2(new_n783), .A3(new_n729), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n784), .A3(new_n427), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n497), .A3(new_n781), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n778), .B1(KEYINPUT42), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G131), .ZN(G33));
  NAND3_X1  g602(.A1(new_n443), .A2(new_n497), .A3(new_n775), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT105), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n664), .A2(new_n652), .A3(new_n666), .A4(new_n716), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT105), .B1(new_n789), .B2(new_n792), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  INV_X1    g611(.A(new_n300), .ZN(new_n798));
  NAND2_X1  g612(.A1(G469), .A2(G902), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n293), .B1(new_n273), .B2(new_n274), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n290), .A2(new_n295), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n193), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n298), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n287), .A2(KEYINPUT45), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n804), .A2(KEYINPUT106), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT106), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n799), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n798), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n807), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(KEYINPUT106), .A3(new_n805), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT46), .A4(new_n799), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT46), .B(new_n799), .C1(new_n806), .C2(new_n807), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT107), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n303), .A3(new_n710), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT108), .Z(new_n820));
  OR3_X1    g634(.A1(new_n556), .A2(KEYINPUT43), .A3(new_n648), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT43), .B1(new_n556), .B2(new_n648), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n669), .A2(new_n821), .A3(new_n677), .A4(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT44), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n825), .A2(new_n826), .A3(new_n780), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  NAND2_X1  g643(.A1(new_n818), .A2(new_n303), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT47), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n818), .A2(KEYINPUT47), .A3(new_n303), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n443), .A2(new_n780), .A3(new_n717), .A4(new_n497), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT109), .Z(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n385), .A2(new_n388), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n626), .A2(new_n840), .A3(new_n386), .A4(new_n652), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n668), .A2(new_n677), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n777), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n757), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n723), .A2(new_n624), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n639), .A2(new_n702), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n697), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n743), .A2(KEYINPUT101), .A3(new_n556), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n443), .A2(new_n497), .A3(new_n723), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n724), .B1(new_n667), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n556), .A2(new_n649), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT112), .B1(new_n613), .B2(new_n615), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n701), .A2(new_n856), .A3(new_n614), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n763), .A2(new_n855), .A3(new_n766), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n624), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n637), .A2(new_n859), .A3(new_n860), .A4(new_n652), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n738), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n766), .A2(new_n716), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n855), .B2(new_n857), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n443), .A2(new_n664), .A3(new_n865), .A4(new_n677), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n760), .B2(new_n770), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(new_n781), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n851), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n785), .A2(new_n497), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT42), .B1(new_n870), .B2(new_n776), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n777), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n796), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n744), .A2(new_n745), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT113), .B1(new_n676), .B2(new_n716), .ZN(new_n877));
  INV_X1    g691(.A(new_n488), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n483), .B2(new_n484), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n493), .B1(new_n879), .B2(new_n487), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT113), .ZN(new_n881));
  NOR4_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n675), .A4(new_n685), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n695), .B(new_n652), .C1(new_n877), .C2(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n688), .B(new_n719), .C1(new_n876), .C2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n875), .B1(new_n884), .B2(new_n772), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT100), .ZN(new_n886));
  AOI21_X1  g700(.A(G902), .B1(new_n635), .B2(new_n428), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n629), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n754), .B1(new_n440), .B2(new_n752), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n779), .A2(new_n677), .A3(new_n737), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n848), .A2(new_n849), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n877), .A2(new_n882), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n892), .A3(new_n652), .A4(new_n695), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n676), .B1(new_n730), .B2(new_n427), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n687), .C1(new_n686), .C2(new_n718), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT52), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n885), .A2(new_n896), .A3(KEYINPUT114), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT114), .B1(new_n885), .B2(new_n896), .ZN(new_n898));
  OAI211_X1 g712(.A(KEYINPUT53), .B(new_n874), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n900));
  NAND4_X1  g714(.A1(new_n734), .A2(new_n724), .A3(new_n738), .A4(new_n861), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n627), .B(new_n678), .C1(new_n746), .C2(new_n757), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n787), .A3(new_n796), .A4(new_n868), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n885), .A2(new_n896), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n899), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n874), .B1(new_n897), .B2(new_n898), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n904), .A2(new_n905), .ZN(new_n911));
  INV_X1    g725(.A(new_n900), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n909), .A2(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n821), .A2(new_n822), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n757), .A2(new_n915), .A3(new_n619), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n737), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n723), .A2(new_n775), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n918), .A2(new_n695), .A3(new_n496), .A4(new_n619), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n767), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n617), .A3(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n870), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n915), .A2(new_n918), .A3(new_n619), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n924), .A2(KEYINPUT48), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(KEYINPUT48), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n923), .A2(new_n677), .A3(new_n889), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n919), .A2(new_n697), .A3(new_n648), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n723), .A2(new_n638), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT117), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n723), .A2(new_n935), .A3(new_n638), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n936), .A3(new_n708), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n916), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n940));
  AOI21_X1  g754(.A(KEYINPUT119), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n821), .A2(new_n822), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n497), .A3(new_n620), .A4(new_n889), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT119), .B(new_n940), .C1(new_n943), .C2(new_n937), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n916), .A3(KEYINPUT50), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT51), .B(new_n932), .C1(new_n941), .C2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n740), .A2(new_n303), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n832), .A2(new_n833), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n943), .A2(new_n780), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n928), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT116), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n932), .B1(new_n941), .B2(new_n946), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(KEYINPUT51), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n839), .B1(new_n914), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n951), .A2(new_n952), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n927), .B1(new_n962), .B2(new_n947), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n953), .A2(KEYINPUT116), .ZN(new_n964));
  INV_X1    g778(.A(new_n958), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT51), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n911), .A2(new_n912), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n885), .A2(new_n896), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT114), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n885), .A2(new_n896), .A3(KEYINPUT114), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n904), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n970), .B1(KEYINPUT53), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT54), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n969), .A2(new_n977), .A3(KEYINPUT120), .A4(new_n908), .ZN(new_n978));
  NOR2_X1   g792(.A1(G952), .A2(G953), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT121), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n961), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n497), .A2(new_n386), .A3(new_n303), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n982), .A2(new_n556), .A3(new_n648), .ZN(new_n983));
  AOI22_X1  g797(.A1(new_n983), .A2(KEYINPUT110), .B1(KEYINPUT49), .B2(new_n740), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(KEYINPUT110), .B2(new_n983), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT111), .Z(new_n986));
  OR2_X1    g800(.A1(new_n740), .A2(KEYINPUT49), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n986), .A2(new_n708), .A3(new_n696), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n981), .A2(new_n988), .ZN(G75));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n912), .B1(new_n874), .B2(new_n971), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n975), .B2(KEYINPUT53), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n992), .B2(new_n299), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n899), .A2(new_n906), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(KEYINPUT122), .A3(G902), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n993), .A2(new_n306), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n338), .A2(new_n350), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(new_n348), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT55), .ZN(new_n999));
  XNOR2_X1  g813(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n996), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n189), .A2(G952), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n994), .A2(G210), .A3(G902), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT56), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1003), .B1(new_n1006), .B2(new_n999), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1002), .A2(new_n1007), .ZN(G51));
  INV_X1    g822(.A(new_n908), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n907), .B1(new_n899), .B2(new_n906), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n799), .B(KEYINPUT57), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n297), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n993), .A2(new_n811), .A3(new_n812), .A4(new_n995), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1003), .B1(new_n1013), .B2(new_n1014), .ZN(G54));
  AND2_X1   g829(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n993), .A2(new_n995), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n541), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1003), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n993), .A2(new_n534), .A3(new_n995), .A4(new_n1016), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(G60));
  INV_X1    g835(.A(KEYINPUT124), .ZN(new_n1022));
  INV_X1    g836(.A(new_n645), .ZN(new_n1023));
  NAND2_X1  g837(.A1(G478), .A2(G902), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1024), .B(KEYINPUT59), .Z(new_n1025));
  NOR2_X1   g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n994), .A2(KEYINPUT54), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(new_n908), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1022), .B1(new_n1029), .B2(new_n1003), .ZN(new_n1030));
  OAI211_X1 g844(.A(KEYINPUT124), .B(new_n1019), .C1(new_n1011), .C2(new_n1027), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1025), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n914), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1023), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(G63));
  NAND2_X1  g849(.A1(G217), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT60), .Z(new_n1037));
  NAND2_X1  g851(.A1(new_n994), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n479), .A2(new_n482), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n674), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n994), .A2(new_n1041), .A3(new_n1037), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1040), .A2(new_n1019), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(KEYINPUT61), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1043), .B(new_n1044), .ZN(G66));
  INV_X1    g859(.A(new_n622), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n345), .B1(new_n1046), .B2(G224), .ZN(new_n1047));
  INV_X1    g861(.A(new_n903), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1047), .B1(new_n1048), .B2(new_n189), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n997), .B1(G898), .B2(new_n189), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1049), .B(new_n1050), .Z(G69));
  AND2_X1   g865(.A1(new_n890), .A2(new_n895), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(new_n714), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT62), .ZN(new_n1054));
  XNOR2_X1  g868(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n790), .A2(new_n652), .A3(new_n710), .A4(new_n859), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n828), .A2(new_n1055), .A3(new_n837), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n189), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n420), .A2(new_n431), .ZN(new_n1059));
  XNOR2_X1  g873(.A(new_n514), .B(KEYINPUT125), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  AND4_X1   g876(.A1(new_n787), .A2(new_n837), .A3(new_n796), .A4(new_n1052), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n820), .A2(new_n891), .A3(new_n922), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n1063), .A2(new_n189), .A3(new_n1064), .A4(new_n828), .ZN(new_n1065));
  INV_X1    g879(.A(new_n189), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1061), .B1(G900), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g882(.A(KEYINPUT126), .ZN(new_n1069));
  NAND3_X1  g883(.A1(new_n1062), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g886(.A(new_n1071), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n1062), .A2(new_n1068), .A3(new_n1069), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g888(.A1(new_n1072), .A2(new_n1074), .ZN(G72));
  OAI21_X1  g889(.A(new_n433), .B1(new_n423), .B2(new_n424), .ZN(new_n1076));
  XNOR2_X1  g890(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g891(.A1(G472), .A2(G902), .ZN(new_n1078));
  XNOR2_X1  g892(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  NAND2_X1  g893(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g894(.A(new_n1019), .B1(new_n913), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g895(.A1(new_n423), .A2(new_n408), .ZN(new_n1082));
  NAND4_X1  g896(.A1(new_n1063), .A2(new_n828), .A3(new_n1064), .A4(new_n903), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n1082), .B1(new_n1083), .B2(new_n1079), .ZN(new_n1084));
  OAI21_X1  g898(.A(new_n1079), .B1(new_n1057), .B2(new_n1048), .ZN(new_n1085));
  AOI211_X1 g899(.A(new_n1081), .B(new_n1084), .C1(new_n1085), .C2(new_n693), .ZN(G57));
endmodule


