//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1120, new_n1121;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n458), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n463), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(G136), .B2(new_n477), .ZN(G162));
  NAND2_X1  g053(.A1(new_n472), .A2(G126), .ZN(new_n479));
  MUX2_X1   g054(.A(G102), .B(G114), .S(G2105), .Z(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n477), .A2(G138), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(KEYINPUT65), .A3(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT65), .A2(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n477), .A2(G138), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n482), .B1(new_n484), .B2(new_n486), .ZN(G164));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G543), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n490));
  INV_X1    g065(.A(G543), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(KEYINPUT66), .A3(G543), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(G88), .B1(G50), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n494), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(G166));
  AND2_X1   g081(.A1(new_n496), .A2(G89), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n494), .A2(G63), .A3(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT7), .ZN(new_n510));
  INV_X1    g085(.A(G51), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n508), .B(new_n510), .C1(new_n497), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G168));
  XOR2_X1   g088(.A(KEYINPUT70), .B(G90), .Z(new_n514));
  AOI22_X1  g089(.A1(new_n496), .A2(new_n514), .B1(G52), .B2(new_n498), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G77), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n494), .B2(G64), .ZN(new_n519));
  OAI21_X1  g094(.A(G651), .B1(new_n519), .B2(KEYINPUT68), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n521));
  AOI211_X1 g096(.A(new_n521), .B(new_n518), .C1(new_n494), .C2(G64), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT69), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n491), .A2(KEYINPUT5), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n488), .A2(KEYINPUT66), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(KEYINPUT66), .B1(new_n488), .B2(G543), .ZN(new_n526));
  OAI211_X1 g101(.A(G64), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n517), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n500), .B1(new_n528), .B2(new_n521), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n519), .A2(KEYINPUT68), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n516), .B1(new_n523), .B2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n494), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n535), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(G651), .A3(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n496), .A2(G81), .B1(G43), .B2(new_n498), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G860), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT72), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n495), .A2(G53), .A3(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G91), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n494), .A2(new_n495), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n494), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n500), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n550), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g134(.A1(new_n555), .A2(new_n550), .A3(new_n557), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n559), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NOR2_X1   g137(.A1(G171), .A2(new_n562), .ZN(new_n563));
  AOI211_X1 g138(.A(KEYINPUT75), .B(new_n516), .C1(new_n523), .C2(new_n532), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n498), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n494), .B2(G74), .ZN(new_n569));
  INV_X1    g144(.A(G87), .ZN(new_n570));
  OAI211_X1 g145(.A(new_n568), .B(new_n569), .C1(new_n570), .C2(new_n554), .ZN(G288));
  AOI22_X1  g146(.A1(new_n496), .A2(G86), .B1(G48), .B2(new_n498), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT76), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n572), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n494), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n500), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT77), .B(G47), .Z(new_n583));
  OAI22_X1  g158(.A1(new_n554), .A2(new_n582), .B1(new_n497), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n496), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n575), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G54), .B2(new_n498), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n595), .B2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n587), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT78), .B2(new_n587), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(KEYINPUT78), .B2(new_n587), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G860), .ZN(G148));
  NOR2_X1   g180(.A1(new_n540), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n590), .A2(new_n594), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n606), .B1(new_n608), .B2(G868), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n477), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  MUX2_X1   g190(.A(G99), .B(G111), .S(G2105), .Z(new_n616));
  AOI22_X1  g191(.A1(new_n472), .A2(G123), .B1(G2104), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n465), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT80), .ZN(new_n620));
  INV_X1    g195(.A(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n615), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(new_n638), .A3(KEYINPUT14), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n632), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n632), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(G14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n647), .B2(new_n644), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(KEYINPUT85), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(KEYINPUT85), .B2(new_n651), .ZN(new_n653));
  INV_X1    g228(.A(new_n644), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n654), .A2(new_n646), .A3(new_n649), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n621), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  INV_X1    g244(.A(new_n664), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n662), .A2(new_n663), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XOR2_X1   g253(.A(G1981), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G229));
  NOR2_X1   g256(.A1(G6), .A2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G305), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(G16), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT91), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT32), .B(G1981), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT92), .B(G1971), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n688), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT33), .B(G1976), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  NOR4_X1   g274(.A1(new_n687), .A2(new_n693), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n477), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n472), .A2(G119), .ZN(new_n705));
  MUX2_X1   g280(.A(G95), .B(G107), .S(G2105), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2104), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT88), .B(G29), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n708), .S(new_n710), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n688), .A2(G24), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT89), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n585), .B2(new_n688), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n717), .A2(G1986), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(G1986), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n714), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n702), .A2(new_n703), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT24), .B(G34), .ZN(new_n723));
  AOI22_X1  g298(.A1(G160), .A2(G29), .B1(new_n709), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G2084), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G11), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT94), .B(G28), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT30), .ZN(new_n728));
  AOI22_X1  g303(.A1(G129), .A2(new_n472), .B1(new_n477), .B2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n459), .A2(G105), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND3_X1  g307(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G32), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n726), .B1(G29), .B2(new_n728), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n735), .A2(G33), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT25), .B1(new_n459), .B2(G103), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n464), .A2(G127), .ZN(new_n744));
  NAND2_X1  g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n458), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n743), .B(new_n746), .C1(G139), .C2(new_n477), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n735), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n725), .B(new_n739), .C1(G2072), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n709), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n472), .A2(G128), .ZN(new_n753));
  MUX2_X1   g328(.A(G104), .B(G116), .S(G2105), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2104), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(new_n757), .B2(new_n735), .ZN(new_n758));
  INV_X1    g333(.A(G2067), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n724), .A2(G2084), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT93), .Z(new_n762));
  OAI22_X1  g337(.A1(new_n748), .A2(G2072), .B1(new_n620), .B2(new_n709), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n737), .B2(new_n738), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n749), .A2(new_n760), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G19), .ZN(new_n766));
  INV_X1    g341(.A(new_n540), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n710), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n710), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G2090), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n710), .A2(G27), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G164), .B2(new_n710), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT96), .B(G2078), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n774), .A2(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n688), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n688), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n775), .A2(new_n779), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n765), .A2(new_n769), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G5), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G171), .B2(G16), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT95), .Z(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n688), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n601), .B2(new_n688), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT98), .B(G1956), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n595), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1348), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n789), .A2(G1961), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n786), .A2(new_n790), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n722), .A2(new_n802), .ZN(G311));
  INV_X1    g378(.A(G311), .ZN(G150));
  AOI22_X1  g379(.A1(new_n494), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n500), .ZN(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n554), .A2(new_n807), .B1(new_n808), .B2(new_n497), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n541), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT37), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n540), .B(new_n810), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT38), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n607), .A2(new_n604), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n541), .B1(new_n817), .B2(KEYINPUT39), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n812), .B1(new_n818), .B2(new_n819), .ZN(G145));
  XNOR2_X1  g395(.A(new_n482), .B(KEYINPUT101), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n484), .A2(KEYINPUT100), .A3(new_n486), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n484), .A2(new_n486), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n756), .ZN(new_n827));
  MUX2_X1   g402(.A(G106), .B(G118), .S(G2105), .Z(new_n828));
  AOI22_X1  g403(.A1(new_n472), .A2(G130), .B1(G2104), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G142), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n465), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n708), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n613), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n827), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n747), .B(new_n734), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(G162), .B(G160), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n620), .ZN(new_n838));
  AOI21_X1  g413(.A(G37), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n836), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g416(.A(new_n810), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(G868), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n696), .B(new_n585), .ZN(new_n844));
  NAND2_X1  g419(.A1(G166), .A2(G305), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n504), .A2(new_n505), .A3(new_n683), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n844), .A3(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n595), .B1(new_n560), .B2(new_n559), .ZN(new_n851));
  INV_X1    g426(.A(new_n560), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n852), .A3(new_n558), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n813), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n608), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n813), .B1(G559), .B2(new_n607), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  AND3_X1   g435(.A1(new_n851), .A2(new_n860), .A3(new_n853), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n851), .B2(new_n853), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(new_n857), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n859), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n850), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n871));
  INV_X1    g446(.A(new_n850), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n843), .B1(new_n875), .B2(G868), .ZN(G295));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n877));
  XNOR2_X1  g452(.A(G295), .B(new_n877), .ZN(G331));
  NAND2_X1  g453(.A1(new_n850), .A2(KEYINPUT105), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n848), .A2(new_n880), .A3(new_n849), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n861), .A2(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n851), .A2(new_n860), .A3(new_n853), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT107), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT104), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n520), .A2(KEYINPUT69), .A3(new_n522), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n515), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT75), .ZN(new_n891));
  NAND2_X1  g466(.A1(G171), .A2(new_n562), .ZN(new_n892));
  AOI21_X1  g467(.A(G286), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(G171), .A2(G168), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(G168), .B1(new_n563), .B2(new_n564), .ZN(new_n896));
  INV_X1    g471(.A(new_n894), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(KEYINPUT104), .A3(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n895), .A2(new_n855), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n855), .B1(new_n895), .B2(new_n898), .ZN(new_n900));
  OAI221_X1 g475(.A(new_n883), .B1(new_n862), .B2(new_n886), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n893), .A2(new_n887), .A3(new_n894), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT104), .B1(new_n896), .B2(new_n897), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n813), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n895), .A2(new_n855), .A3(new_n898), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n854), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n882), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n863), .B1(new_n899), .B2(new_n900), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n850), .A3(new_n906), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n908), .A2(new_n906), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n910), .B(new_n909), .C1(new_n916), .C2(new_n882), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(KEYINPUT44), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n882), .B1(new_n908), .B2(new_n906), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n921), .B(KEYINPUT43), .C1(new_n911), .C2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n882), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n883), .B1(new_n862), .B2(new_n886), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n905), .B2(new_n904), .ZN(new_n926));
  INV_X1    g501(.A(new_n906), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n910), .A4(new_n909), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n921), .B1(new_n917), .B2(KEYINPUT43), .ZN(new_n932));
  OAI211_X1 g507(.A(KEYINPUT108), .B(new_n920), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n911), .B2(new_n922), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n923), .A3(new_n930), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT108), .B1(new_n937), .B2(new_n920), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n919), .B1(new_n934), .B2(new_n938), .ZN(G397));
  INV_X1    g514(.A(G1384), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT45), .B1(new_n826), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G160), .A2(G40), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(G1996), .A3(new_n733), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT110), .Z(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(G1996), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n756), .B(G2067), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n948), .A2(new_n734), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n708), .A2(new_n713), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n708), .A2(new_n713), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n944), .A2(G1986), .A3(G290), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT48), .Z(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n951), .A2(new_n953), .B1(new_n759), .B2(new_n757), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(new_n944), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT127), .Z(new_n962));
  NOR2_X1   g537(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT126), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n949), .A2(new_n733), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n962), .B(new_n964), .C1(new_n944), .C2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  NOR2_X1   g542(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n826), .A2(new_n940), .A3(new_n943), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT113), .B(G8), .Z(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n578), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(G305), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n972), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n977), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n979), .A2(KEYINPUT115), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(KEYINPUT115), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1976), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n972), .B1(new_n989), .B2(G288), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n696), .A2(G1976), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n990), .A2(KEYINPUT52), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(KEYINPUT52), .B2(new_n990), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n988), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(G164), .A2(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NOR2_X1   g572(.A1(G164), .A2(G1384), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n826), .A2(new_n940), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1001), .B(new_n943), .C1(KEYINPUT50), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(G2084), .ZN(new_n1004));
  OR3_X1    g579(.A1(new_n941), .A2(KEYINPUT120), .A3(new_n942), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT120), .B1(new_n941), .B2(new_n942), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(new_n783), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(G286), .A3(new_n971), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n826), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n942), .B1(new_n995), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1971), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT112), .B(G2090), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1003), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT55), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n994), .A2(new_n1010), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT63), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n696), .A2(new_n989), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n987), .A2(new_n1026), .B1(G1981), .B2(G305), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n972), .B(KEYINPUT118), .Z(new_n1028));
  AOI22_X1  g603(.A1(new_n994), .A2(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n971), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G286), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1009), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1032), .B1(new_n1009), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n1032), .C1(new_n1009), .C2(new_n971), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2078), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1041), .B1(new_n1014), .B2(G2078), .ZN(new_n1044));
  INV_X1    g619(.A(G1961), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1003), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G301), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1047), .A2(KEYINPUT62), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1040), .A2(new_n1049), .B1(new_n1050), .B2(new_n1010), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(KEYINPUT62), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT121), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1011), .A2(new_n1013), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n555), .A2(new_n557), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT57), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n826), .A2(KEYINPUT50), .A3(new_n940), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n995), .A2(new_n999), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n942), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1056), .B(new_n1058), .C1(new_n1061), .C2(G1956), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT122), .ZN(new_n1063));
  INV_X1    g638(.A(G1348), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1003), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n969), .A2(G2067), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n607), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1056), .B1(new_n1061), .B2(G1956), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1058), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1063), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  AOI211_X1 g648(.A(new_n595), .B(new_n1066), .C1(new_n1003), .C2(new_n1064), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT60), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT58), .B(G1341), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1014), .A2(G1996), .B1(new_n970), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n767), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT59), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1080), .A3(new_n767), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1071), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n607), .A2(KEYINPUT60), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1065), .A2(new_n1067), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(new_n1082), .A3(new_n1083), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1071), .A2(KEYINPUT123), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1069), .A2(new_n1088), .A3(new_n1070), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1063), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1073), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n941), .A2(new_n942), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1011), .A3(new_n1042), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1046), .A2(new_n1044), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n1095), .B2(new_n1048), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1094), .A2(new_n1044), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(G301), .A4(new_n1046), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1052), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1095), .B2(G171), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1053), .B1(new_n1092), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1051), .B1(new_n1105), .B2(new_n1040), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n988), .A2(new_n993), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1061), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1016), .B1(new_n1110), .B2(new_n1017), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1031), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1025), .B1(new_n1021), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1108), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1030), .B1(new_n1106), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n585), .B(G1986), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n955), .B1(new_n944), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n968), .B1(new_n1115), .B2(new_n1117), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g693(.A(G319), .ZN(new_n1120));
  NOR4_X1   g694(.A1(G401), .A2(new_n1120), .A3(G229), .A4(G227), .ZN(new_n1121));
  NAND3_X1  g695(.A1(new_n937), .A2(new_n840), .A3(new_n1121), .ZN(G225));
  INV_X1    g696(.A(G225), .ZN(G308));
endmodule


