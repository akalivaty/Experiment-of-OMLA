

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n540), .B(n539), .ZN(G164) );
  INV_X1 U556 ( .A(G2105), .ZN(n530) );
  BUF_X1 U557 ( .A(n898), .Z(n524) );
  XNOR2_X1 U558 ( .A(n531), .B(KEYINPUT17), .ZN(n898) );
  AND2_X1 U559 ( .A1(n719), .A2(n807), .ZN(n721) );
  INV_X1 U560 ( .A(KEYINPUT26), .ZN(n720) );
  XNOR2_X1 U561 ( .A(n546), .B(n545), .ZN(n548) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n545) );
  XNOR2_X1 U563 ( .A(n721), .B(n720), .ZN(n726) );
  XNOR2_X1 U564 ( .A(n755), .B(n754), .ZN(n760) );
  INV_X1 U565 ( .A(KEYINPUT94), .ZN(n539) );
  XNOR2_X1 U566 ( .A(n552), .B(KEYINPUT66), .ZN(G160) );
  NAND2_X1 U567 ( .A1(G303), .A2(n759), .ZN(n525) );
  OR2_X1 U568 ( .A1(G1971), .A2(G303), .ZN(n526) );
  AND2_X1 U569 ( .A1(n726), .A2(n725), .ZN(n527) );
  INV_X1 U570 ( .A(n983), .ZN(n723) );
  AND2_X1 U571 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U572 ( .A1(n707), .A2(n765), .ZN(n708) );
  INV_X1 U573 ( .A(KEYINPUT29), .ZN(n747) );
  INV_X1 U574 ( .A(KEYINPUT105), .ZN(n754) );
  NAND2_X1 U575 ( .A1(n779), .A2(n526), .ZN(n780) );
  OR2_X2 U576 ( .A1(n781), .A2(n780), .ZN(n822) );
  INV_X1 U577 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n530), .ZN(n901) );
  NOR2_X1 U579 ( .A1(G651), .A2(n653), .ZN(n668) );
  NAND2_X1 U580 ( .A1(n530), .A2(G2104), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT67), .ZN(n637) );
  NAND2_X1 U582 ( .A1(G102), .A2(n637), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U584 ( .A1(G138), .A2(n898), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U586 ( .A(n534), .B(KEYINPUT93), .ZN(n538) );
  NAND2_X1 U587 ( .A1(G126), .A2(n901), .ZN(n536) );
  AND2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n902) );
  NAND2_X1 U589 ( .A1(G114), .A2(n902), .ZN(n535) );
  AND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n902), .A2(G113), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT69), .B(n541), .Z(n543) );
  NAND2_X1 U594 ( .A1(n898), .A2(G137), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U596 ( .A(KEYINPUT70), .B(n544), .ZN(n551) );
  NAND2_X1 U597 ( .A1(n637), .A2(G101), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n901), .A2(G125), .ZN(n547) );
  NAND2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U600 ( .A(n549), .B(KEYINPUT68), .ZN(n550) );
  NOR2_X1 U601 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U602 ( .A(G2438), .B(G2454), .Z(n554) );
  XNOR2_X1 U603 ( .A(G2435), .B(G2430), .ZN(n553) );
  XNOR2_X1 U604 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U605 ( .A(n555), .B(G2427), .Z(n557) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n556) );
  XNOR2_X1 U607 ( .A(n557), .B(n556), .ZN(n561) );
  XOR2_X1 U608 ( .A(G2443), .B(G2446), .Z(n559) );
  XNOR2_X1 U609 ( .A(KEYINPUT108), .B(G2451), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U611 ( .A(n561), .B(n560), .Z(n562) );
  AND2_X1 U612 ( .A1(G14), .A2(n562), .ZN(G401) );
  XOR2_X1 U613 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  NAND2_X1 U614 ( .A1(G52), .A2(n668), .ZN(n565) );
  INV_X1 U615 ( .A(G651), .ZN(n566) );
  NOR2_X1 U616 ( .A1(G543), .A2(n566), .ZN(n563) );
  XOR2_X1 U617 ( .A(KEYINPUT1), .B(n563), .Z(n669) );
  NAND2_X1 U618 ( .A1(G64), .A2(n669), .ZN(n564) );
  NAND2_X1 U619 ( .A1(n565), .A2(n564), .ZN(n571) );
  NOR2_X1 U620 ( .A1(G651), .A2(G543), .ZN(n676) );
  NAND2_X1 U621 ( .A1(G90), .A2(n676), .ZN(n568) );
  NOR2_X1 U622 ( .A1(n653), .A2(n566), .ZN(n673) );
  NAND2_X1 U623 ( .A1(G77), .A2(n673), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U626 ( .A1(n571), .A2(n570), .ZN(G171) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G132), .ZN(G219) );
  INV_X1 U630 ( .A(G82), .ZN(G220) );
  NAND2_X1 U631 ( .A1(G88), .A2(n676), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G75), .A2(n673), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G50), .A2(n668), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G62), .A2(n669), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U637 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U638 ( .A(G166), .ZN(G303) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT10), .ZN(n579) );
  XNOR2_X1 U641 ( .A(KEYINPUT74), .B(n579), .ZN(G223) );
  XNOR2_X1 U642 ( .A(KEYINPUT75), .B(G223), .ZN(n849) );
  NAND2_X1 U643 ( .A1(n849), .A2(G567), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  XNOR2_X1 U645 ( .A(KEYINPUT77), .B(KEYINPUT13), .ZN(n586) );
  NAND2_X1 U646 ( .A1(G81), .A2(n676), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT12), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT76), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G68), .A2(n673), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n669), .A2(G56), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n587), .Z(n588) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n668), .A2(G43), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n983) );
  NAND2_X1 U657 ( .A1(n723), .A2(G860), .ZN(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U660 ( .A1(G92), .A2(n676), .ZN(n593) );
  NAND2_X1 U661 ( .A1(G79), .A2(n673), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G54), .A2(n668), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G66), .A2(n669), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT15), .B(n598), .Z(n985) );
  OR2_X1 U668 ( .A1(n985), .A2(G868), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U670 ( .A1(n668), .A2(G51), .ZN(n601) );
  XNOR2_X1 U671 ( .A(KEYINPUT81), .B(n601), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n669), .A2(G63), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT80), .B(n602), .Z(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(KEYINPUT6), .B(n605), .ZN(n613) );
  NAND2_X1 U676 ( .A1(G89), .A2(n676), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT78), .ZN(n607) );
  XNOR2_X1 U678 ( .A(n607), .B(KEYINPUT4), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G76), .A2(n673), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n611) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n610) );
  XNOR2_X1 U682 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n614), .B(KEYINPUT7), .ZN(n615) );
  XNOR2_X1 U685 ( .A(KEYINPUT82), .B(n615), .ZN(G168) );
  XOR2_X1 U686 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U687 ( .A1(G91), .A2(n676), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G78), .A2(n673), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G65), .A2(n669), .ZN(n618) );
  XNOR2_X1 U691 ( .A(KEYINPUT73), .B(n618), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n668), .A2(G53), .ZN(n621) );
  NAND2_X1 U694 ( .A1(n622), .A2(n621), .ZN(G299) );
  XNOR2_X1 U695 ( .A(KEYINPUT83), .B(G868), .ZN(n623) );
  NOR2_X1 U696 ( .A1(G286), .A2(n623), .ZN(n626) );
  NOR2_X1 U697 ( .A1(G868), .A2(G299), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n624), .B(KEYINPUT84), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n626), .A2(n625), .ZN(G297) );
  INV_X1 U700 ( .A(G559), .ZN(n627) );
  NOR2_X1 U701 ( .A1(G860), .A2(n627), .ZN(n628) );
  XNOR2_X1 U702 ( .A(KEYINPUT85), .B(n628), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n629), .A2(n985), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U705 ( .A1(G868), .A2(n983), .ZN(n631) );
  XNOR2_X1 U706 ( .A(KEYINPUT86), .B(n631), .ZN(n634) );
  NAND2_X1 U707 ( .A1(G868), .A2(n985), .ZN(n632) );
  NOR2_X1 U708 ( .A1(G559), .A2(n632), .ZN(n633) );
  NOR2_X1 U709 ( .A1(n634), .A2(n633), .ZN(G282) );
  NAND2_X1 U710 ( .A1(G123), .A2(n901), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT18), .B(n635), .Z(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(KEYINPUT87), .ZN(n639) );
  BUF_X1 U713 ( .A(n637), .Z(n897) );
  NAND2_X1 U714 ( .A1(G99), .A2(n897), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G111), .A2(n902), .ZN(n641) );
  NAND2_X1 U717 ( .A1(G135), .A2(n524), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n937) );
  XNOR2_X1 U720 ( .A(n937), .B(G2096), .ZN(n645) );
  INV_X1 U721 ( .A(G2100), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G156) );
  NAND2_X1 U723 ( .A1(G86), .A2(n676), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G61), .A2(n669), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n673), .A2(G73), .ZN(n648) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n668), .A2(G48), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n668), .ZN(n655) );
  NAND2_X1 U732 ( .A1(G87), .A2(n653), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n669), .A2(n656), .ZN(n659) );
  NAND2_X1 U735 ( .A1(G74), .A2(G651), .ZN(n657) );
  XOR2_X1 U736 ( .A(KEYINPUT91), .B(n657), .Z(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(G288) );
  NAND2_X1 U738 ( .A1(G47), .A2(n668), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT72), .B(n660), .Z(n665) );
  NAND2_X1 U740 ( .A1(G85), .A2(n676), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G72), .A2(n673), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U743 ( .A(KEYINPUT71), .B(n663), .Z(n664) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n669), .A2(G60), .ZN(n666) );
  NAND2_X1 U746 ( .A1(n667), .A2(n666), .ZN(G290) );
  INV_X1 U747 ( .A(G868), .ZN(n681) );
  NAND2_X1 U748 ( .A1(G55), .A2(n668), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G67), .A2(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(KEYINPUT89), .ZN(n675) );
  NAND2_X1 U752 ( .A1(G80), .A2(n673), .ZN(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U754 ( .A1(n676), .A2(G93), .ZN(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT88), .B(n677), .Z(n678) );
  NOR2_X1 U756 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U757 ( .A(KEYINPUT90), .B(n680), .Z(n856) );
  NAND2_X1 U758 ( .A1(n681), .A2(n856), .ZN(n682) );
  XNOR2_X1 U759 ( .A(n682), .B(KEYINPUT92), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n856), .B(G305), .ZN(n683) );
  XNOR2_X1 U761 ( .A(n683), .B(G288), .ZN(n684) );
  XOR2_X1 U762 ( .A(n684), .B(KEYINPUT19), .Z(n686) );
  INV_X1 U763 ( .A(G299), .ZN(n990) );
  XNOR2_X1 U764 ( .A(n990), .B(G166), .ZN(n685) );
  XNOR2_X1 U765 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U766 ( .A(n687), .B(G290), .ZN(n920) );
  NAND2_X1 U767 ( .A1(G559), .A2(n985), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n688), .B(n983), .ZN(n854) );
  XNOR2_X1 U769 ( .A(n920), .B(n854), .ZN(n689) );
  NAND2_X1 U770 ( .A1(G868), .A2(n689), .ZN(n690) );
  NAND2_X1 U771 ( .A1(n691), .A2(n690), .ZN(G295) );
  NAND2_X1 U772 ( .A1(G2078), .A2(G2084), .ZN(n692) );
  XOR2_X1 U773 ( .A(KEYINPUT20), .B(n692), .Z(n693) );
  NAND2_X1 U774 ( .A1(G2090), .A2(n693), .ZN(n694) );
  XNOR2_X1 U775 ( .A(KEYINPUT21), .B(n694), .ZN(n695) );
  NAND2_X1 U776 ( .A1(n695), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U777 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U778 ( .A1(G220), .A2(G219), .ZN(n696) );
  XOR2_X1 U779 ( .A(KEYINPUT22), .B(n696), .Z(n697) );
  NOR2_X1 U780 ( .A1(G218), .A2(n697), .ZN(n698) );
  NAND2_X1 U781 ( .A1(G96), .A2(n698), .ZN(n857) );
  NAND2_X1 U782 ( .A1(n857), .A2(G2106), .ZN(n702) );
  NAND2_X1 U783 ( .A1(G69), .A2(G120), .ZN(n699) );
  NOR2_X1 U784 ( .A1(G237), .A2(n699), .ZN(n700) );
  NAND2_X1 U785 ( .A1(G108), .A2(n700), .ZN(n858) );
  NAND2_X1 U786 ( .A1(n858), .A2(G567), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n702), .A2(n701), .ZN(n931) );
  NAND2_X1 U788 ( .A1(G661), .A2(G483), .ZN(n703) );
  NOR2_X1 U789 ( .A1(n931), .A2(n703), .ZN(n853) );
  NAND2_X1 U790 ( .A1(n853), .A2(G36), .ZN(G176) );
  NAND2_X1 U791 ( .A1(G40), .A2(G160), .ZN(n806) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n705) );
  INV_X1 U793 ( .A(KEYINPUT64), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n705), .B(n704), .ZN(n718) );
  NOR2_X1 U795 ( .A1(n806), .A2(n718), .ZN(n722) );
  INV_X1 U796 ( .A(n722), .ZN(n756) );
  NOR2_X1 U797 ( .A1(n756), .A2(G2084), .ZN(n706) );
  XNOR2_X1 U798 ( .A(n706), .B(KEYINPUT97), .ZN(n766) );
  NAND2_X1 U799 ( .A1(G8), .A2(n766), .ZN(n707) );
  NAND2_X1 U800 ( .A1(G8), .A2(n756), .ZN(n783) );
  NOR2_X1 U801 ( .A1(G1966), .A2(n783), .ZN(n765) );
  XOR2_X1 U802 ( .A(KEYINPUT30), .B(n708), .Z(n709) );
  NOR2_X1 U803 ( .A1(G168), .A2(n709), .ZN(n715) );
  BUF_X1 U804 ( .A(n722), .Z(n738) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n967) );
  NAND2_X1 U806 ( .A1(n738), .A2(n967), .ZN(n710) );
  XNOR2_X1 U807 ( .A(n710), .B(KEYINPUT99), .ZN(n712) );
  XNOR2_X1 U808 ( .A(G1961), .B(KEYINPUT98), .ZN(n1017) );
  NOR2_X1 U809 ( .A1(n1017), .A2(n738), .ZN(n711) );
  NOR2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U811 ( .A(KEYINPUT100), .B(n713), .Z(n749) );
  NOR2_X1 U812 ( .A1(G171), .A2(n749), .ZN(n714) );
  NOR2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U814 ( .A(n716), .B(KEYINPUT103), .ZN(n717) );
  XNOR2_X1 U815 ( .A(n717), .B(KEYINPUT31), .ZN(n753) );
  INV_X1 U816 ( .A(G1996), .ZN(n968) );
  NOR2_X1 U817 ( .A1(n806), .A2(n968), .ZN(n719) );
  INV_X1 U818 ( .A(n718), .ZN(n807) );
  NAND2_X1 U819 ( .A1(n756), .A2(G1341), .ZN(n724) );
  INV_X1 U820 ( .A(KEYINPUT65), .ZN(n727) );
  XNOR2_X1 U821 ( .A(n527), .B(n727), .ZN(n729) );
  NOR2_X1 U822 ( .A1(n729), .A2(n985), .ZN(n728) );
  XNOR2_X1 U823 ( .A(n728), .B(KEYINPUT101), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n729), .A2(n985), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n738), .A2(G1348), .ZN(n731) );
  NOR2_X1 U826 ( .A1(G2067), .A2(n756), .ZN(n730) );
  NOR2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U830 ( .A(n736), .B(KEYINPUT102), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n738), .A2(G2072), .ZN(n737) );
  XNOR2_X1 U832 ( .A(n737), .B(KEYINPUT27), .ZN(n740) );
  INV_X1 U833 ( .A(G1956), .ZN(n1018) );
  NOR2_X1 U834 ( .A1(n1018), .A2(n738), .ZN(n739) );
  NOR2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n743), .A2(n990), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n743), .A2(n990), .ZN(n744) );
  XOR2_X1 U839 ( .A(n744), .B(KEYINPUT28), .Z(n745) );
  NAND2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U841 ( .A(n748), .B(n747), .ZN(n751) );
  NAND2_X1 U842 ( .A1(G171), .A2(n749), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n763) );
  NAND2_X1 U845 ( .A1(n763), .A2(G286), .ZN(n755) );
  NOR2_X1 U846 ( .A1(G1971), .A2(n783), .ZN(n758) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n525), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n761), .A2(G8), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(KEYINPUT32), .ZN(n772) );
  INV_X1 U852 ( .A(n763), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n769) );
  INV_X1 U854 ( .A(n766), .ZN(n767) );
  NAND2_X1 U855 ( .A1(G8), .A2(n767), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U857 ( .A(KEYINPUT104), .B(n770), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n825) );
  INV_X1 U859 ( .A(n825), .ZN(n781) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n773) );
  XOR2_X1 U861 ( .A(KEYINPUT106), .B(n773), .Z(n993) );
  INV_X1 U862 ( .A(KEYINPUT33), .ZN(n774) );
  AND2_X1 U863 ( .A1(n993), .A2(n774), .ZN(n778) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U865 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  NOR2_X1 U866 ( .A1(n783), .A2(n776), .ZN(n789) );
  INV_X1 U867 ( .A(n789), .ZN(n777) );
  AND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  INV_X1 U869 ( .A(n783), .ZN(n826) );
  NAND2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n994) );
  AND2_X1 U871 ( .A1(n826), .A2(n994), .ZN(n782) );
  NOR2_X1 U872 ( .A1(KEYINPUT33), .A2(n782), .ZN(n787) );
  XOR2_X1 U873 ( .A(G1981), .B(G305), .Z(n1001) );
  NOR2_X1 U874 ( .A1(n783), .A2(n993), .ZN(n784) );
  NAND2_X1 U875 ( .A1(KEYINPUT33), .A2(n784), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n1001), .A2(n785), .ZN(n786) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  OR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n820) );
  NAND2_X1 U879 ( .A1(G95), .A2(n897), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G131), .A2(n524), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G119), .A2(n901), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G107), .A2(n902), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n893) );
  INV_X1 U886 ( .A(G1991), .ZN(n963) );
  NOR2_X1 U887 ( .A1(n893), .A2(n963), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G105), .A2(n897), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT38), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G129), .A2(n901), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G117), .A2(n902), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G141), .A2(n524), .ZN(n799) );
  XNOR2_X1 U894 ( .A(KEYINPUT95), .B(n799), .ZN(n800) );
  NOR2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n908) );
  AND2_X1 U897 ( .A1(n908), .A2(G1996), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n940) );
  NOR2_X1 U899 ( .A1(n806), .A2(n807), .ZN(n844) );
  XOR2_X1 U900 ( .A(n844), .B(KEYINPUT96), .Z(n808) );
  NOR2_X1 U901 ( .A1(n940), .A2(n808), .ZN(n837) );
  INV_X1 U902 ( .A(n837), .ZN(n818) );
  NAND2_X1 U903 ( .A1(G104), .A2(n897), .ZN(n810) );
  NAND2_X1 U904 ( .A1(G140), .A2(n524), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT34), .B(n811), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G128), .A2(n901), .ZN(n813) );
  NAND2_X1 U908 ( .A1(G116), .A2(n902), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U910 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT36), .B(n817), .ZN(n917) );
  XNOR2_X1 U913 ( .A(KEYINPUT37), .B(G2067), .ZN(n842) );
  NOR2_X1 U914 ( .A1(n917), .A2(n842), .ZN(n942) );
  NAND2_X1 U915 ( .A1(n844), .A2(n942), .ZN(n840) );
  NAND2_X1 U916 ( .A1(n818), .A2(n840), .ZN(n827) );
  INV_X1 U917 ( .A(n827), .ZN(n819) );
  AND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n831) );
  NOR2_X1 U920 ( .A1(G2090), .A2(G303), .ZN(n823) );
  NAND2_X1 U921 ( .A1(G8), .A2(n823), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U926 ( .A(G1986), .B(G290), .ZN(n989) );
  NAND2_X1 U927 ( .A1(n989), .A2(n844), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n847) );
  NOR2_X1 U929 ( .A1(G1996), .A2(n908), .ZN(n951) );
  AND2_X1 U930 ( .A1(n963), .A2(n893), .ZN(n834) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(n834), .Z(n938) );
  NOR2_X1 U932 ( .A1(G1986), .A2(G290), .ZN(n835) );
  NOR2_X1 U933 ( .A1(n938), .A2(n835), .ZN(n836) );
  NOR2_X1 U934 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U935 ( .A1(n951), .A2(n838), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT39), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n917), .A2(n842), .ZN(n943) );
  NAND2_X1 U939 ( .A1(n843), .A2(n943), .ZN(n845) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U941 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U942 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n851) );
  XOR2_X1 U947 ( .A(KEYINPUT109), .B(n851), .Z(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(G188) );
  NOR2_X1 U950 ( .A1(G860), .A2(n854), .ZN(n855) );
  XOR2_X1 U951 ( .A(n856), .B(n855), .Z(G145) );
  INV_X1 U952 ( .A(G120), .ZN(G236) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  XOR2_X1 U957 ( .A(KEYINPUT111), .B(G1971), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1961), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n861), .B(KEYINPUT110), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U963 ( .A(G1976), .B(G1981), .Z(n865) );
  XNOR2_X1 U964 ( .A(G1966), .B(G1956), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U967 ( .A(G2474), .B(KEYINPUT41), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(G229) );
  XOR2_X1 U969 ( .A(G2100), .B(G2096), .Z(n871) );
  XNOR2_X1 U970 ( .A(KEYINPUT42), .B(G2678), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U972 ( .A(KEYINPUT43), .B(G2090), .Z(n873) );
  XNOR2_X1 U973 ( .A(G2067), .B(G2072), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U976 ( .A(G2078), .B(G2084), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(G227) );
  NAND2_X1 U978 ( .A1(G100), .A2(n897), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G112), .A2(n902), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT112), .B(n880), .ZN(n885) );
  NAND2_X1 U982 ( .A1(n901), .A2(G124), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n881), .B(KEYINPUT44), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G136), .A2(n524), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  NOR2_X1 U986 ( .A1(n885), .A2(n884), .ZN(G162) );
  NAND2_X1 U987 ( .A1(G130), .A2(n901), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G118), .A2(n902), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G106), .A2(n897), .ZN(n889) );
  NAND2_X1 U991 ( .A1(G142), .A2(n524), .ZN(n888) );
  NAND2_X1 U992 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U993 ( .A(KEYINPUT45), .B(n890), .Z(n891) );
  NOR2_X1 U994 ( .A1(n892), .A2(n891), .ZN(n912) );
  XOR2_X1 U995 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n895) );
  XNOR2_X1 U996 ( .A(n893), .B(KEYINPUT46), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U998 ( .A(n896), .B(n937), .Z(n910) );
  NAND2_X1 U999 ( .A1(G103), .A2(n897), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(G139), .A2(n524), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G127), .A2(n901), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G115), .A2(n902), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n932) );
  XOR2_X1 U1007 ( .A(n908), .B(n932), .Z(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(G160), .B(G162), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(G164), .B(n915), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G395) );
  XNOR2_X1 U1015 ( .A(n985), .B(n983), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(G286), .ZN(n922) );
  XOR2_X1 U1017 ( .A(G171), .B(n920), .Z(n921) );
  XNOR2_X1 U1018 ( .A(n922), .B(n921), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n923), .ZN(G397) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n924), .B(KEYINPUT49), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT115), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(G401), .A2(n931), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT114), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(n931), .ZN(G319) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n958) );
  XOR2_X1 U1032 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT50), .B(n935), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(n936), .B(KEYINPUT118), .ZN(n949) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1041 ( .A(G2084), .B(G160), .Z(n945) );
  XNOR2_X1 U1042 ( .A(KEYINPUT116), .B(n945), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1047 ( .A(KEYINPUT117), .B(n952), .Z(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(KEYINPUT51), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n956), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(G29), .ZN(n1043) );
  XOR2_X1 U1053 ( .A(G2090), .B(G35), .Z(n962) );
  XOR2_X1 U1054 ( .A(G34), .B(KEYINPUT54), .Z(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(G2084), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n978) );
  XNOR2_X1 U1057 ( .A(G25), .B(n963), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G28), .ZN(n974) );
  XNOR2_X1 U1059 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(G33), .B(G2072), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n972) );
  XOR2_X1 U1062 ( .A(n967), .B(G27), .Z(n970) );
  XOR2_X1 U1063 ( .A(n968), .B(G32), .Z(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1067 ( .A(KEYINPUT53), .B(n975), .Z(n976) );
  XNOR2_X1 U1068 ( .A(n976), .B(KEYINPUT119), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1070 ( .A(KEYINPUT55), .B(n979), .Z(n980) );
  NOR2_X1 U1071 ( .A1(G29), .A2(n980), .ZN(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT120), .B(n981), .Z(n982) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n982), .ZN(n1041) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  XNOR2_X1 U1075 ( .A(G1341), .B(KEYINPUT124), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n984), .B(n983), .ZN(n987) );
  XOR2_X1 U1077 ( .A(G1348), .B(n985), .Z(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n1008) );
  XNOR2_X1 U1079 ( .A(G1961), .B(G301), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n1000) );
  XNOR2_X1 U1081 ( .A(G166), .B(G1971), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n990), .B(G1956), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(KEYINPUT122), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(n998), .Z(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT57), .B(n1003), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(KEYINPUT121), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1039) );
  INV_X1 U1096 ( .A(G16), .ZN(n1037) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1976), .B(G23), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1016), .ZN(n1033) );
  XNOR2_X1 U1104 ( .A(n1017), .B(G5), .ZN(n1031) );
  XNOR2_X1 U1105 ( .A(G20), .B(n1018), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G19), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G1981), .B(G6), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT59), .B(G1348), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(G4), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(KEYINPUT60), .B(n1026), .Z(n1028) );
  XNOR2_X1 U1114 ( .A(G1966), .B(G21), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(KEYINPUT125), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(n1034), .B(KEYINPUT127), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1035), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1123 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1124 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1044), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

