//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT93), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G1gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n204), .A2(KEYINPUT94), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G8gat), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n204), .A2(new_n210), .A3(KEYINPUT94), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n216));
  OR3_X1    g015(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n217), .A2(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT91), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n222), .A2(KEYINPUT15), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT92), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n225));
  NOR3_X1   g024(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n222), .B2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n219), .ZN(new_n228));
  OAI22_X1  g027(.A1(new_n221), .A2(new_n223), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n229), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n229), .B(new_n215), .Z(new_n237));
  XOR2_X1   g036(.A(new_n231), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  INV_X1    g040(.A(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT11), .B(G169gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n235), .A2(new_n236), .A3(new_n239), .A4(new_n246), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G85gat), .A2(G92gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT7), .ZN(new_n253));
  OR2_X1    g052(.A1(G99gat), .A2(G106gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G85gat), .ZN(new_n258));
  INV_X1    g057(.A(G92gat), .ZN(new_n259));
  AOI22_X1  g058(.A1(KEYINPUT8), .A2(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT96), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n261), .B(new_n263), .Z(new_n264));
  OR2_X1    g063(.A1(G57gat), .A2(G64gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G57gat), .A2(G64gat), .ZN(new_n266));
  AND2_X1   g065(.A1(G71gat), .A2(G78gat), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(KEYINPUT9), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT95), .B1(G71gat), .B2(G78gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G71gat), .A2(G78gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n272), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n261), .B(new_n263), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT10), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n264), .A2(KEYINPUT10), .A3(new_n275), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G230gat), .A2(G233gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n279), .ZN(new_n286));
  INV_X1    g085(.A(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G120gat), .B(G148gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G176gat), .B(G204gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n285), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n251), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n299), .B(new_n229), .Z(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G232gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT41), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n300), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n300), .A2(new_n304), .ZN(new_n306));
  XOR2_X1   g105(.A(G134gat), .B(G162gat), .Z(new_n307));
  XNOR2_X1  g106(.A(G190gat), .B(G218gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OR3_X1    g109(.A1(new_n305), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n305), .B2(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n215), .B1(new_n275), .B2(KEYINPUT21), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT21), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n275), .B(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n316), .B2(new_n215), .ZN(new_n317));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G211gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n317), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G155gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n322), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G106gat), .ZN(new_n329));
  XOR2_X1   g128(.A(G50gat), .B(G78gat), .Z(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(KEYINPUT86), .B2(G22gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(G22gat), .B2(new_n331), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT73), .ZN(new_n338));
  XNOR2_X1  g137(.A(G197gat), .B(G204gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT22), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G218gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n336), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n339), .A2(new_n343), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(new_n336), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n344), .A2(new_n337), .A3(KEYINPUT74), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  AND2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G141gat), .B(G148gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT2), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n360), .A2(G141gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(G141gat), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(G148gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n364), .B2(new_n356), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n354), .B(new_n359), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT78), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  INV_X1    g167(.A(G162gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n368), .B2(new_n369), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n360), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n371), .B1(new_n374), .B2(new_n361), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n354), .A4(new_n359), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n367), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n353), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT83), .B(KEYINPUT29), .C1(new_n367), .C2(new_n377), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n335), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  AND2_X1   g182(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n385));
  OAI21_X1  g184(.A(G148gat), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n361), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n360), .A2(G141gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n364), .B1(new_n361), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n388), .A2(new_n371), .B1(new_n390), .B2(new_n357), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n376), .B1(new_n391), .B2(new_n354), .ZN(new_n392));
  AND4_X1   g191(.A1(new_n376), .A2(new_n375), .A3(new_n354), .A4(new_n359), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n383), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n379), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(KEYINPUT84), .A3(new_n396), .A4(new_n353), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n352), .B2(new_n383), .ZN(new_n398));
  OAI211_X1 g197(.A(G228gat), .B(G233gat), .C1(new_n398), .C2(new_n391), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n382), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n382), .A2(new_n397), .A3(new_n400), .A4(KEYINPUT85), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n350), .A2(new_n351), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n349), .A2(new_n336), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n383), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n354), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n375), .A2(new_n359), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n353), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n334), .B1(new_n405), .B2(new_n416), .ZN(new_n417));
  AOI211_X1 g216(.A(new_n333), .B(new_n415), .C1(new_n403), .C2(new_n404), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G169gat), .ZN(new_n422));
  INV_X1    g221(.A(G176gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT26), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT26), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G169gat), .B2(G176gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n427), .A2(new_n428), .B1(G183gat), .B2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  INV_X1    g229(.A(G190gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n319), .B2(KEYINPUT27), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435));
  AOI21_X1  g234(.A(G190gat), .B1(new_n435), .B2(G183gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n319), .A2(KEYINPUT27), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n436), .A2(new_n433), .A3(new_n430), .A4(new_n437), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n429), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n443));
  AND3_X1   g242(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT23), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT23), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(G169gat), .B2(G176gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n428), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n428), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n450), .A3(KEYINPUT25), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n447), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n452), .A2(KEYINPUT66), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n443), .C1(new_n447), .C2(new_n451), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n442), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(KEYINPUT69), .A2(G134gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G113gat), .B(G120gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(KEYINPUT1), .ZN(new_n465));
  INV_X1    g264(.A(G120gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(G113gat), .ZN(new_n467));
  INV_X1    g266(.A(G113gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G120gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT1), .ZN(new_n471));
  INV_X1    g270(.A(G134gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G127gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n465), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n465), .B2(new_n473), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n452), .A2(KEYINPUT66), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n456), .A2(new_n457), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n460), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n441), .ZN(new_n483));
  INV_X1    g282(.A(new_n478), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n421), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT71), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT71), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n479), .A2(new_n485), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n420), .B(KEYINPUT64), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT34), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(G15gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(G43gat), .ZN(new_n499));
  XOR2_X1   g298(.A(G71gat), .B(G99gat), .Z(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n479), .A2(new_n485), .A3(new_n494), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(KEYINPUT32), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n502), .B(KEYINPUT32), .C1(new_n503), .C2(new_n501), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n488), .A2(KEYINPUT71), .B1(new_n492), .B2(new_n495), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(new_n491), .A3(new_n507), .A4(new_n506), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n514));
  XNOR2_X1  g313(.A(G1gat), .B(G29gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G57gat), .B(G85gat), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n516), .B(new_n517), .Z(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n410), .A2(KEYINPUT3), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n478), .B(new_n520), .C1(new_n392), .C2(new_n393), .ZN(new_n521));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n465), .A2(new_n473), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G127gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n410), .B1(new_n524), .B2(new_n475), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT4), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n526), .B(new_n391), .C1(new_n476), .C2(new_n477), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n521), .B(new_n522), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n522), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n476), .A2(new_n391), .A3(new_n477), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n525), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT5), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n530), .A2(new_n534), .A3(KEYINPUT79), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n530), .B2(KEYINPUT79), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n519), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(KEYINPUT79), .ZN(new_n538));
  INV_X1    g337(.A(new_n534), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n530), .A2(new_n534), .A3(KEYINPUT79), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n518), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n535), .A2(new_n536), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT81), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT6), .A4(new_n518), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n540), .A2(KEYINPUT6), .A3(new_n541), .A4(new_n518), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT81), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n544), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n419), .A2(new_n513), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G226gat), .A2(G233gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n461), .B2(KEYINPUT29), .ZN(new_n554));
  INV_X1    g353(.A(new_n553), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT75), .B1(new_n483), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557));
  AOI211_X1 g356(.A(new_n557), .B(new_n553), .C1(new_n482), .C2(new_n441), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n352), .B(new_n554), .C1(new_n556), .C2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n555), .B1(new_n483), .B2(new_n383), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n461), .A2(new_n553), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n353), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G8gat), .B(G36gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G64gat), .B(G92gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n559), .A2(new_n562), .A3(KEYINPUT30), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n483), .A2(new_n555), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n352), .B1(new_n554), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n557), .B1(new_n461), .B2(new_n553), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n483), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n560), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(new_n352), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n567), .B1(new_n573), .B2(new_n566), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n562), .A3(new_n566), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n575), .A3(new_n577), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT87), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n566), .B1(new_n559), .B2(new_n562), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n559), .A2(new_n562), .A3(new_n566), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(KEYINPUT30), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n586));
  AND4_X1   g385(.A1(KEYINPUT87), .A2(new_n584), .A3(new_n586), .A4(new_n580), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n552), .A2(new_n588), .A3(KEYINPUT90), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n419), .A2(new_n513), .ZN(new_n591));
  INV_X1    g390(.A(new_n580), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n592), .A2(new_n574), .A3(new_n578), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n550), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT35), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n584), .A2(new_n586), .A3(new_n580), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT87), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n579), .A2(KEYINPUT87), .A3(new_n580), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n589), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n596), .B1(new_n551), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n590), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n509), .A2(new_n511), .A3(new_n604), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n509), .A2(new_n511), .B1(KEYINPUT72), .B2(KEYINPUT36), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n395), .A2(new_n353), .A3(new_n396), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n399), .B1(new_n608), .B2(new_n335), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT85), .B1(new_n609), .B2(new_n397), .ZN(new_n610));
  AND4_X1   g409(.A1(KEYINPUT85), .A2(new_n382), .A3(new_n397), .A4(new_n400), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n416), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n333), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n405), .A2(new_n416), .A3(new_n334), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND4_X1   g414(.A1(new_n544), .A2(new_n547), .A3(new_n549), .A4(new_n576), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT89), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT37), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n559), .A2(new_n618), .A3(new_n562), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n565), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n353), .B(new_n554), .C1(new_n556), .C2(new_n558), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n352), .B1(new_n560), .B2(new_n561), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT37), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT38), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n617), .B1(new_n620), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n554), .A2(new_n568), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n618), .B1(new_n627), .B2(new_n352), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT38), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n629), .A2(KEYINPUT89), .A3(new_n565), .A4(new_n619), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n618), .B1(new_n559), .B2(new_n562), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT38), .B1(new_n620), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n626), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n615), .B1(new_n616), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n521), .B1(new_n527), .B2(new_n529), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n531), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n532), .A2(new_n525), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n522), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n637), .A3(new_n531), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n519), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT40), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n542), .B1(new_n642), .B2(new_n644), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n643), .B1(new_n642), .B2(new_n644), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n649), .B1(new_n581), .B2(new_n587), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n607), .B1(new_n634), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n594), .A2(new_n615), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n298), .B(new_n327), .C1(new_n603), .C2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n550), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  INV_X1    g456(.A(new_n588), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(KEYINPUT97), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n659), .A2(new_n213), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT97), .B2(new_n663), .ZN(G1325gat));
  AOI21_X1  g467(.A(G15gat), .B1(new_n654), .B2(new_n513), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n607), .A2(G15gat), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n654), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n615), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  AOI21_X1  g473(.A(new_n313), .B1(new_n603), .B2(new_n653), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n652), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n594), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n605), .A2(new_n606), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n642), .A2(new_n644), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n642), .A2(new_n644), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n542), .A4(new_n645), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n599), .B2(new_n600), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n544), .A2(new_n547), .A3(new_n549), .A4(new_n576), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n626), .A2(new_n632), .A3(new_n630), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n419), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n682), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n681), .A2(new_n691), .A3(KEYINPUT99), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n594), .A2(KEYINPUT98), .A3(new_n615), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT98), .B1(new_n594), .B2(new_n615), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n693), .B1(new_n696), .B2(new_n651), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n603), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n313), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n676), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n677), .B1(new_n700), .B2(KEYINPUT100), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT99), .B1(new_n681), .B2(new_n691), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n651), .A3(new_n693), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n313), .B1(new_n705), .B2(new_n603), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n702), .B1(new_n706), .B2(new_n676), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n298), .A2(new_n326), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n655), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G29gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n675), .A2(new_n709), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(G29gat), .A3(new_n550), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT45), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(G1328gat));
  OAI211_X1 g514(.A(new_n658), .B(new_n709), .C1(new_n701), .C2(new_n707), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G36gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n588), .A2(G36gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n675), .A2(new_n709), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n675), .A2(new_n723), .A3(new_n709), .A4(new_n719), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(new_n724), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(KEYINPUT46), .ZN(new_n728));
  AOI211_X1 g527(.A(KEYINPUT102), .B(new_n722), .C1(new_n721), .C2(new_n724), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT103), .B1(new_n718), .B2(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n732), .A2(new_n733), .A3(new_n717), .A4(new_n725), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(G1329gat));
  OAI211_X1 g534(.A(new_n607), .B(new_n709), .C1(new_n701), .C2(new_n707), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n712), .A2(G43gat), .A3(new_n512), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(KEYINPUT47), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1330gat));
  OR3_X1    g542(.A1(new_n712), .A2(G50gat), .A3(new_n419), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n744), .A2(KEYINPUT48), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n615), .B(new_n709), .C1(new_n701), .C2(new_n707), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n747));
  OAI21_X1  g546(.A(G50gat), .B1(new_n746), .B2(KEYINPUT104), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(G50gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n744), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(G1331gat));
  NAND2_X1  g553(.A1(new_n251), .A2(new_n296), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n327), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT105), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n705), .B2(new_n603), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n655), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT106), .B(G57gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1332gat));
  AOI21_X1  g560(.A(new_n588), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT107), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n764), .B(new_n765), .Z(G1333gat));
  AOI21_X1  g565(.A(G71gat), .B1(new_n758), .B2(new_n513), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n607), .A2(G71gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n767), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n615), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n326), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n708), .A2(new_n655), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G85gat), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n250), .A2(new_n326), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n698), .A2(new_n699), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n698), .A2(KEYINPUT51), .A3(new_n699), .A4(new_n776), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(KEYINPUT108), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n780), .A2(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n296), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n655), .A2(new_n258), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n775), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  INV_X1    g588(.A(new_n296), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n588), .A2(G92gat), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n781), .A2(new_n782), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT110), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n781), .A2(new_n782), .A3(new_n794), .A4(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n658), .B(new_n773), .C1(new_n701), .C2(new_n707), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(new_n797), .B2(G92gat), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(G92gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n780), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n791), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n803), .ZN(G1337gat));
  OAI211_X1 g603(.A(new_n607), .B(new_n773), .C1(new_n701), .C2(new_n707), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(KEYINPUT111), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(G99gat), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n512), .A2(G99gat), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n785), .A2(new_n296), .A3(new_n786), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1338gat));
  OAI211_X1 g610(.A(new_n615), .B(new_n773), .C1(new_n701), .C2(new_n707), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n419), .A2(G106gat), .A3(new_n790), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n783), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n815), .B(KEYINPUT112), .Z(new_n818));
  AOI22_X1  g617(.A1(new_n812), .A2(G106gat), .B1(new_n801), .B2(new_n818), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n813), .A2(new_n817), .B1(new_n819), .B2(new_n814), .ZN(G1339gat));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n237), .A2(new_n238), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n245), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT114), .B(new_n245), .C1(new_n822), .C2(new_n823), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n249), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n821), .B1(new_n828), .B2(new_n790), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n296), .A3(KEYINPUT115), .A4(new_n249), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n281), .A2(new_n282), .A3(new_n287), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n281), .A2(new_n835), .A3(new_n282), .A4(new_n287), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n834), .A2(new_n285), .A3(KEYINPUT54), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n287), .B1(new_n281), .B2(new_n282), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n294), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n837), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n295), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n251), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n313), .B1(new_n832), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n313), .A2(new_n845), .A3(new_n828), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n326), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n251), .A2(new_n313), .A3(new_n790), .A4(new_n326), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n588), .A2(new_n655), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n591), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n250), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n468), .A2(KEYINPUT116), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n468), .A2(KEYINPUT116), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n856), .B2(new_n857), .ZN(G1340gat));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n296), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n326), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT69), .B(G127gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1342gat));
  NAND3_X1  g664(.A1(new_n855), .A2(new_n472), .A3(new_n699), .ZN(new_n866));
  AND2_X1   g665(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n867));
  NOR2_X1   g666(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n855), .A2(new_n699), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G134gat), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n869), .B(new_n871), .C1(new_n866), .C2(new_n867), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n607), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(new_n853), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n615), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n844), .A2(new_n295), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT55), .B1(new_n837), .B2(new_n840), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n843), .A2(KEYINPUT119), .A3(new_n295), .A4(new_n844), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n250), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n830), .A2(new_n249), .A3(new_n296), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n699), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(KEYINPUT120), .A3(new_n884), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n848), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n851), .B1(new_n889), .B2(new_n326), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(KEYINPUT57), .A3(new_n615), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n877), .B1(new_n891), .B2(KEYINPUT121), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT57), .A4(new_n615), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n874), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n362), .B1(new_n895), .B2(new_n250), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n853), .A2(new_n419), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n873), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(G141gat), .A3(new_n251), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT58), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  INV_X1    g700(.A(new_n899), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n251), .B(new_n874), .C1(new_n892), .C2(new_n894), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n362), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(new_n898), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n360), .A3(new_n296), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n615), .B(new_n875), .C1(new_n850), .C2(new_n852), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT122), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT57), .B1(new_n890), .B2(new_n615), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n296), .B(new_n873), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT123), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n360), .B1(new_n912), .B2(KEYINPUT123), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT59), .B(new_n360), .C1(new_n895), .C2(new_n296), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n906), .B2(new_n326), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n326), .A2(G155gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n895), .B2(new_n919), .ZN(G1346gat));
  NAND3_X1  g719(.A1(new_n906), .A2(new_n369), .A3(new_n699), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n895), .A2(new_n922), .A3(new_n699), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G162gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n895), .B2(new_n699), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1347gat));
  NOR3_X1   g725(.A1(new_n853), .A2(new_n551), .A3(new_n588), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n250), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n296), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g730(.A(new_n319), .B1(new_n927), .B2(new_n326), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(KEYINPUT60), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n435), .A2(G183gat), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n927), .A2(new_n935), .A3(new_n437), .A4(new_n326), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n933), .A2(KEYINPUT60), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n937), .B(new_n938), .Z(G1350gat));
  NAND2_X1  g738(.A1(new_n927), .A2(new_n699), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G190gat), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(KEYINPUT61), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n945), .A2(new_n946), .B1(G190gat), .B2(new_n940), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n588), .A2(new_n607), .A3(new_n655), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n897), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT127), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n242), .A3(new_n250), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n910), .A2(new_n911), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(new_n948), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(new_n250), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n954), .B2(new_n242), .ZN(G1352gat));
  INV_X1    g754(.A(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n956), .A3(new_n296), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  AND3_X1   g757(.A1(new_n952), .A2(new_n296), .A3(new_n948), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n956), .B2(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n950), .A2(new_n341), .A3(new_n326), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n326), .A3(new_n948), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n950), .B2(new_n699), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n313), .A2(new_n342), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n953), .B2(new_n967), .ZN(G1355gat));
endmodule


