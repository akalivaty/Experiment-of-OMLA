//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G128), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(new_n196), .C1(G119), .C2(new_n195), .ZN(new_n197));
  XNOR2_X1  g011(.A(G119), .B(G128), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  AOI22_X1  g013(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT77), .B(G125), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n201), .A2(KEYINPUT16), .A3(G140), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  NOR2_X1   g017(.A1(G125), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT77), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n204), .B1(new_n209), .B2(G140), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n204), .ZN(new_n213));
  INV_X1    g027(.A(G140), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n201), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT78), .A3(KEYINPUT16), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n202), .B1(new_n212), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  AOI211_X1 g033(.A(new_n219), .B(new_n202), .C1(new_n212), .C2(new_n216), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n200), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G146), .ZN(new_n222));
  XOR2_X1   g036(.A(G125), .B(G140), .Z(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT79), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT65), .A2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT65), .A2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n197), .A2(G110), .B1(new_n198), .B2(new_n199), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n222), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G953), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(KEYINPUT80), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G137), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n231), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n221), .A2(new_n230), .A3(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n191), .B1(new_n240), .B2(new_n188), .ZN(new_n241));
  AOI211_X1 g055(.A(G902), .B(new_n190), .C1(new_n238), .C2(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n189), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n189), .A2(G902), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n244), .B(KEYINPUT82), .Z(new_n245));
  NAND2_X1  g059(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n252), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n219), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT65), .A2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G143), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n219), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(KEYINPUT0), .A3(G128), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n219), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n261), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g087(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n265), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT66), .B1(new_n258), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n251), .A2(KEYINPUT67), .A3(G134), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n249), .B2(G137), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n251), .A2(G134), .ZN(new_n281));
  OAI211_X1 g095(.A(G131), .B(new_n278), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n257), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n262), .A2(new_n264), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n195), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n288), .B2(new_n270), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n283), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n266), .B1(new_n227), .B2(G143), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n273), .A2(new_n274), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n271), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n255), .A2(new_n257), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .A4(new_n265), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n277), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT69), .A2(G116), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT69), .A2(G116), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n302), .A2(new_n303), .A3(new_n193), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G119), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n301), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n301), .ZN(new_n308));
  OR2_X1    g122(.A1(KEYINPUT69), .A2(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT69), .A2(G116), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(G119), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n306), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n315), .B(new_n301), .C1(new_n304), .C2(new_n306), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n278), .A2(G131), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n251), .A2(G134), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n253), .A3(new_n279), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT68), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT71), .B1(new_n284), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n320), .A2(KEYINPUT68), .A3(G131), .A4(new_n278), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n290), .A2(new_n323), .A3(new_n324), .A4(new_n257), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n325), .A3(new_n289), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n294), .A2(new_n295), .A3(new_n265), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n300), .A2(new_n317), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n314), .A2(new_n316), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n232), .A3(G210), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(KEYINPUT27), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT31), .ZN(new_n339));
  INV_X1    g153(.A(new_n336), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n298), .A2(new_n317), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(new_n331), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n331), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n340), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT31), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n329), .A2(new_n337), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT72), .B1(new_n338), .B2(KEYINPUT31), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G472), .A2(G902), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT74), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT32), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n352), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n284), .A2(new_n321), .ZN(new_n359));
  AOI22_X1  g173(.A1(KEYINPUT66), .A2(new_n327), .B1(new_n359), .B2(new_n289), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n330), .B1(new_n360), .B2(new_n297), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n326), .A2(new_n330), .A3(new_n327), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n341), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n346), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(new_n340), .B1(KEYINPUT31), .B2(new_n338), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT32), .ZN(new_n367));
  INV_X1    g181(.A(new_n356), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n357), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n330), .B1(new_n326), .B2(new_n327), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT28), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n340), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n346), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n188), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT76), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT76), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n378), .A3(new_n188), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n363), .A2(new_n336), .A3(new_n346), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n373), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n329), .A2(new_n331), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT75), .B1(new_n383), .B2(new_n340), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n385), .B(new_n336), .C1(new_n329), .C2(new_n331), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n382), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G472), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n247), .B1(new_n370), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G214), .B1(G237), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(G234), .A2(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G952), .A3(new_n232), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(G902), .A3(G953), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT21), .B(G898), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  INV_X1    g215(.A(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G107), .ZN(new_n403));
  INV_X1    g217(.A(G107), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n405), .B2(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT3), .B1(new_n402), .B2(G107), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(KEYINPUT83), .B(KEYINPUT3), .C1(new_n402), .C2(G107), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G101), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n401), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  OAI21_X1  g228(.A(G101), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n402), .A2(KEYINPUT3), .A3(G107), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n404), .A2(G104), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT83), .B1(new_n405), .B2(KEYINPUT3), .ZN(new_n419));
  INV_X1    g233(.A(new_n410), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n418), .B(new_n414), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n413), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n317), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n412), .B1(new_n425), .B2(KEYINPUT84), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n401), .A4(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(KEYINPUT84), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n429), .A2(new_n401), .A3(G101), .A4(new_n421), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT85), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n424), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT86), .B1(new_n404), .B2(G104), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT86), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n402), .A3(G107), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n435), .A3(new_n405), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G101), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n418), .B(new_n412), .C1(new_n419), .C2(new_n420), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(KEYINPUT87), .A3(G101), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n311), .A2(KEYINPUT5), .A3(new_n312), .ZN(new_n443));
  INV_X1    g257(.A(G113), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT5), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n306), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(new_n313), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n400), .B1(new_n432), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n431), .A2(new_n428), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n426), .A2(new_n421), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n330), .B1(new_n453), .B2(new_n413), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n399), .A3(new_n449), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n289), .A2(new_n201), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n276), .B2(new_n201), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n232), .A2(G224), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n399), .B1(new_n455), .B2(new_n449), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n466));
  NOR4_X1   g280(.A1(new_n466), .A2(KEYINPUT91), .A3(KEYINPUT6), .A4(new_n399), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n457), .B(new_n461), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT92), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n443), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n311), .A2(KEYINPUT92), .A3(KEYINPUT5), .A4(new_n312), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n446), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n439), .A2(new_n440), .A3(new_n313), .A4(new_n441), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT93), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n442), .A2(new_n476), .A3(new_n472), .A4(new_n313), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n477), .C1(new_n448), .C2(new_n442), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n399), .B(KEYINPUT8), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n459), .B(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n456), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT94), .A3(new_n188), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT94), .B1(new_n483), .B2(new_n188), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n468), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n468), .B(new_n488), .C1(new_n485), .C2(new_n486), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n391), .B(new_n398), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n309), .A2(G122), .A3(new_n310), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n302), .A2(new_n303), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT97), .A3(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n305), .A2(G122), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n404), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n498), .A2(new_n404), .A3(new_n500), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(G107), .B(new_n499), .C1(new_n495), .C2(new_n497), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT98), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT13), .B1(new_n195), .B2(G143), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(new_n249), .ZN(new_n509));
  XNOR2_X1  g323(.A(G128), .B(G143), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n499), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n495), .A2(new_n497), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n404), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT99), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n510), .B(new_n249), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n504), .A2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT97), .B1(new_n496), .B2(G122), .ZN(new_n521));
  INV_X1    g335(.A(G122), .ZN(new_n522));
  NOR4_X1   g336(.A1(new_n302), .A2(new_n303), .A3(new_n494), .A4(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT14), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n515), .A3(new_n500), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G107), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n504), .A2(new_n518), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT99), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n512), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT9), .B(G234), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n530), .A2(new_n187), .A3(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n512), .B(new_n531), .C1(new_n520), .C2(new_n528), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n188), .ZN(new_n536));
  INV_X1    g350(.A(G478), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT15), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n535), .B(new_n188), .C1(KEYINPUT15), .C2(new_n537), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n402), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n224), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n227), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n332), .A2(new_n232), .A3(G214), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(G143), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n550), .B2(new_n256), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n269), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT95), .A3(G131), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n256), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n222), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n210), .A2(G146), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n228), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n550), .B1(new_n559), .B2(new_n256), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(KEYINPUT18), .A3(G131), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n543), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n218), .A2(new_n220), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n551), .A2(new_n553), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n551), .A2(new_n553), .A3(new_n568), .A4(new_n554), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n564), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n563), .B1(new_n571), .B2(new_n543), .ZN(new_n572));
  NOR2_X1   g386(.A1(G475), .A2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT20), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n563), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n212), .A2(new_n216), .ZN(new_n577));
  INV_X1    g391(.A(new_n202), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n219), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(new_n222), .A3(new_n567), .A4(new_n569), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n543), .A3(new_n562), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n573), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n571), .A2(new_n543), .ZN(new_n587));
  INV_X1    g401(.A(new_n582), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n188), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G475), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n541), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G221), .B1(new_n530), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G469), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n188), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n225), .A2(new_n226), .A3(new_n269), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT1), .ZN(new_n599));
  OAI21_X1  g413(.A(G128), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n263), .B1(new_n227), .B2(G143), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n600), .A2(new_n292), .B1(new_n601), .B2(new_n286), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n195), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n287), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n605), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n295), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT89), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT12), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n258), .B1(new_n603), .B2(new_n606), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT89), .B1(new_n612), .B2(KEYINPUT12), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(KEYINPUT12), .A3(new_n295), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT88), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(KEYINPUT88), .A3(KEYINPUT12), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n276), .B1(new_n453), .B2(new_n413), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n452), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n440), .A2(new_n441), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n289), .A4(new_n439), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n606), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n622), .A2(new_n258), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(G110), .B(G140), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n232), .A2(G227), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT90), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n627), .B1(new_n452), .B2(new_n621), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n258), .ZN(new_n636));
  INV_X1    g450(.A(new_n276), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n423), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n428), .B2(new_n431), .ZN(new_n639));
  OAI211_X1 g453(.A(KEYINPUT90), .B(new_n295), .C1(new_n639), .C2(new_n627), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n633), .B1(new_n635), .B2(new_n258), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n630), .A2(new_n633), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n596), .B1(new_n643), .B2(G469), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n620), .A2(new_n642), .ZN(new_n645));
  INV_X1    g459(.A(new_n629), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n636), .B2(new_n640), .ZN(new_n647));
  INV_X1    g461(.A(new_n633), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n595), .A3(new_n188), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n594), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n389), .A2(new_n492), .A3(new_n592), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  INV_X1    g467(.A(new_n591), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n529), .B2(new_n532), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n517), .B1(new_n516), .B2(new_n519), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT99), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(KEYINPUT100), .A3(new_n512), .A4(new_n531), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n534), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n656), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT101), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n656), .A2(new_n662), .A3(new_n665), .A4(new_n660), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT33), .B1(new_n533), .B2(new_n534), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n537), .A2(G902), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n536), .A2(new_n537), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n654), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n358), .B2(new_n365), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  OAI22_X1  g489(.A1(new_n674), .A2(new_n675), .B1(new_n354), .B2(new_n356), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n247), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n492), .A2(new_n651), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  INV_X1    g495(.A(new_n398), .ZN(new_n682));
  INV_X1    g496(.A(new_n491), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n483), .A2(new_n188), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT94), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n484), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n488), .B1(new_n687), .B2(new_n468), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n390), .B(new_n682), .C1(new_n683), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n584), .B1(new_n583), .B2(new_n573), .ZN(new_n690));
  AOI211_X1 g504(.A(KEYINPUT20), .B(new_n574), .C1(new_n576), .C2(new_n582), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n575), .A2(new_n693), .A3(new_n585), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n590), .A3(new_n541), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n681), .B1(new_n689), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n391), .B1(new_n490), .B2(new_n491), .ZN(new_n698));
  INV_X1    g512(.A(new_n696), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT103), .A4(new_n682), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n651), .A3(new_n677), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  INV_X1    g518(.A(new_n239), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n236), .B1(new_n221), .B2(new_n230), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n188), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n190), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n240), .A2(new_n188), .A3(new_n191), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n231), .B(new_n711), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n710), .A2(new_n189), .B1(new_n245), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n676), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n492), .A2(new_n592), .A3(new_n651), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT37), .B(G110), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G12));
  AOI21_X1  g531(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n718));
  AOI211_X1 g532(.A(KEYINPUT32), .B(new_n356), .C1(new_n358), .C2(new_n365), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n388), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n713), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n651), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT104), .B(G900), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n394), .B1(new_n396), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n695), .A2(new_n590), .A3(new_n541), .A4(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n698), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(new_n727), .B2(new_n698), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n722), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G128), .ZN(G30));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n724), .B(new_n734), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n651), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n490), .A2(new_n491), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT38), .ZN(new_n740));
  INV_X1    g554(.A(new_n383), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n340), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n362), .A2(new_n371), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n188), .B1(new_n743), .B2(new_n336), .ZN(new_n744));
  OAI21_X1  g558(.A(G472), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT106), .B(G472), .C1(new_n742), .C2(new_n744), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n718), .B2(new_n719), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n541), .A2(new_n591), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n390), .A2(new_n750), .A3(new_n713), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n738), .A2(new_n740), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G143), .ZN(G45));
  NAND2_X1  g569(.A1(new_n739), .A2(new_n390), .ZN(new_n756));
  INV_X1    g570(.A(new_n670), .ZN(new_n757));
  AOI211_X1 g571(.A(new_n668), .B(new_n757), .C1(new_n664), .C2(new_n666), .ZN(new_n758));
  INV_X1    g572(.A(new_n672), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n591), .B(new_n725), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n722), .A3(KEYINPUT108), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n698), .A2(new_n673), .A3(new_n725), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n720), .A2(new_n651), .A3(new_n721), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G146), .ZN(G48));
  AOI22_X1  g582(.A1(new_n613), .A2(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n629), .A2(new_n648), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n622), .A2(new_n628), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT90), .B1(new_n772), .B2(new_n295), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n634), .B(new_n258), .C1(new_n622), .C2(new_n628), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n629), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n775), .B2(new_n633), .ZN(new_n776));
  OAI21_X1  g590(.A(G469), .B1(new_n776), .B2(G902), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n593), .A3(new_n650), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT109), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n780), .A3(new_n593), .A4(new_n650), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n389), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n492), .A2(new_n673), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g598(.A(KEYINPUT41), .B(G113), .Z(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G15));
  AND3_X1   g600(.A1(new_n389), .A2(new_n779), .A3(new_n781), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n701), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G116), .ZN(G18));
  AOI21_X1  g603(.A(new_n713), .B1(new_n370), .B2(new_n388), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n649), .A2(new_n595), .A3(new_n188), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n595), .B1(new_n649), .B2(new_n188), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n594), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n541), .A2(new_n591), .A3(new_n398), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n790), .A2(new_n698), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G119), .ZN(G21));
  XOR2_X1   g610(.A(KEYINPUT110), .B(G472), .Z(new_n797));
  NOR2_X1   g611(.A1(new_n674), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n336), .B1(new_n372), .B2(new_n346), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(KEYINPUT31), .B2(new_n338), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n356), .B1(new_n800), .B2(new_n358), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n798), .A2(new_n247), .A3(new_n398), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n779), .A2(new_n802), .A3(new_n781), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n698), .A2(new_n804), .A3(new_n751), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n739), .A2(new_n390), .A3(new_n751), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n522), .ZN(G24));
  NOR3_X1   g623(.A1(new_n798), .A2(new_n713), .A3(new_n801), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n673), .A3(new_n725), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n793), .A2(new_n698), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n205), .ZN(G27));
  INV_X1    g628(.A(KEYINPUT42), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n490), .A2(new_n390), .A3(new_n491), .ZN(new_n816));
  INV_X1    g630(.A(new_n247), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n720), .A3(new_n817), .A4(new_n651), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n815), .B1(new_n818), .B2(new_n760), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n683), .A2(new_n688), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n820), .A2(new_n651), .A3(new_n390), .ZN(new_n821));
  INV_X1    g635(.A(new_n760), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n821), .A2(KEYINPUT42), .A3(new_n389), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G131), .ZN(G33));
  INV_X1    g639(.A(KEYINPUT112), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n818), .B2(new_n726), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n821), .A2(KEYINPUT112), .A3(new_n389), .A4(new_n727), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G134), .ZN(G36));
  INV_X1    g644(.A(new_n596), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n641), .A2(new_n642), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n633), .B1(new_n769), .B2(new_n646), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT45), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n595), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n643), .B2(KEYINPUT45), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n838), .A2(new_n833), .A3(new_n834), .A4(KEYINPUT45), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n832), .B(new_n837), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT113), .B1(new_n835), .B2(new_n836), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n643), .A2(new_n838), .A3(KEYINPUT45), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n832), .B1(new_n845), .B2(new_n837), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n831), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT46), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT46), .B(new_n831), .C1(new_n842), .C2(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n650), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n593), .A3(new_n736), .ZN(new_n852));
  INV_X1    g666(.A(new_n816), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n654), .B1(new_n758), .B2(new_n759), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT43), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(KEYINPUT43), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n721), .A2(new_n676), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT44), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(new_n251), .ZN(G39));
  OAI21_X1  g677(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT114), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n596), .B1(new_n865), .B2(new_n841), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n650), .B1(new_n866), .B2(KEYINPUT46), .ZN(new_n867));
  INV_X1    g681(.A(new_n850), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n593), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT115), .B(KEYINPUT47), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n851), .A2(new_n593), .A3(new_n870), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n853), .A2(new_n760), .A3(new_n720), .A4(new_n817), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(G140), .ZN(G42));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT122), .Z(new_n878));
  AND2_X1   g692(.A1(new_n855), .A2(new_n856), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n853), .A2(new_n393), .A3(new_n778), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n389), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT48), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n370), .A2(new_n817), .A3(new_n749), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n673), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n886), .A2(G952), .A3(new_n232), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n798), .A2(new_n247), .A3(new_n393), .A4(new_n801), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n879), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n883), .B(new_n887), .C1(new_n812), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n853), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n791), .B1(new_n847), .B2(new_n848), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n594), .B(new_n871), .C1(new_n892), .C2(new_n850), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n870), .B1(new_n851), .B2(new_n593), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n791), .A2(new_n792), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n593), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n891), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n793), .A2(new_n391), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n740), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n793), .A2(KEYINPUT120), .A3(new_n391), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT50), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n904), .A2(new_n905), .A3(new_n889), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n904), .B2(new_n889), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n758), .A2(new_n591), .A3(new_n759), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n880), .A2(new_n885), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n912), .A2(new_n913), .B1(new_n810), .B2(new_n881), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT51), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n890), .B1(new_n899), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n898), .B1(new_n872), .B2(new_n873), .ZN(new_n917));
  INV_X1    g731(.A(new_n891), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT119), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n908), .A3(new_n914), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n899), .A2(KEYINPUT119), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n922), .B2(KEYINPUT51), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n807), .A2(new_n805), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n651), .A2(new_n750), .A3(new_n713), .A4(new_n725), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n762), .A2(new_n766), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT105), .B1(new_n756), .B2(new_n726), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n729), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n813), .B1(new_n929), .B2(new_n722), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n927), .A2(KEYINPUT52), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT52), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n720), .A2(new_n721), .A3(new_n794), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n812), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n673), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n689), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n787), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n779), .A2(new_n781), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n925), .A2(new_n939), .A3(new_n802), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n938), .A2(new_n788), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n541), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n591), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n492), .A2(new_n651), .A3(new_n677), .A4(new_n943), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n652), .A2(new_n678), .A3(new_n715), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n816), .A2(new_n651), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT116), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT102), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n693), .B1(new_n575), .B2(new_n585), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n590), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n539), .A2(new_n540), .A3(new_n725), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n539), .A2(new_n540), .A3(new_n725), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(KEYINPUT116), .A3(new_n695), .A4(new_n590), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n952), .A2(new_n720), .A3(new_n721), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n946), .B1(new_n955), .B2(new_n811), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n827), .B2(new_n828), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n941), .A2(new_n824), .A3(new_n945), .A4(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n924), .B1(new_n933), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT54), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT52), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n925), .A2(new_n926), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n767), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n813), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n732), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n927), .A2(KEYINPUT52), .A3(new_n930), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n957), .A2(KEYINPUT53), .A3(new_n945), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n824), .A2(new_n938), .A3(new_n788), .A4(new_n940), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT117), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n795), .B1(new_n782), .B2(new_n783), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n808), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT117), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n788), .A4(new_n824), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n959), .A2(new_n960), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT118), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n933), .A2(new_n958), .A3(new_n924), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n957), .A2(new_n945), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT53), .B1(new_n968), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT54), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT118), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n959), .A2(new_n976), .A3(new_n984), .A4(new_n960), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n978), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n878), .B1(new_n923), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n817), .A2(new_n390), .A3(new_n593), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n740), .A2(new_n750), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n854), .B1(new_n897), .B2(KEYINPUT49), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n989), .B(new_n990), .C1(KEYINPUT49), .C2(new_n897), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(G75));
  OAI21_X1  g806(.A(new_n969), .B1(new_n931), .B2(new_n932), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n971), .A2(new_n975), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(G210), .B(G902), .C1(new_n995), .C2(new_n982), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT56), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n457), .B1(new_n465), .B2(new_n467), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n461), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT55), .Z(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n996), .A2(new_n997), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n996), .B2(new_n997), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n232), .A2(G952), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(G51));
  OAI21_X1  g819(.A(KEYINPUT54), .B1(new_n995), .B2(new_n982), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT123), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n1007), .A3(new_n977), .ZN(new_n1008));
  OAI211_X1 g822(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n995), .C2(new_n982), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n596), .B(KEYINPUT57), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n649), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n995), .A2(new_n982), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(new_n188), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(new_n841), .A3(new_n865), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1004), .B1(new_n1012), .B2(new_n1015), .ZN(G54));
  AND2_X1   g830(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n1014), .A2(new_n583), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n583), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n1018), .A2(new_n1019), .A3(new_n1004), .ZN(G60));
  AOI21_X1  g834(.A(new_n668), .B1(new_n664), .B2(new_n666), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G478), .A2(G902), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT59), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1008), .A2(new_n1021), .A3(new_n1009), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1004), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1021), .B1(new_n986), .B2(new_n1023), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1026), .A2(new_n1027), .ZN(G63));
  INV_X1    g842(.A(KEYINPUT61), .ZN(new_n1029));
  NAND2_X1  g843(.A1(G217), .A2(G902), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT60), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n239), .B(new_n238), .C1(new_n1013), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n1025), .ZN(new_n1033));
  INV_X1    g847(.A(new_n712), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1013), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1029), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1035), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n1037), .A2(KEYINPUT61), .A3(new_n1025), .A4(new_n1032), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1036), .A2(new_n1038), .ZN(G66));
  INV_X1    g853(.A(G224), .ZN(new_n1040));
  OAI21_X1  g854(.A(G953), .B1(new_n397), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n941), .A2(new_n945), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1041), .B1(new_n1043), .B2(G953), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n998), .B1(G898), .B2(new_n232), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1044), .B(new_n1045), .ZN(G69));
  INV_X1    g860(.A(KEYINPUT125), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n925), .A2(new_n389), .ZN(new_n1048));
  NAND4_X1  g862(.A1(new_n851), .A2(new_n593), .A3(new_n1048), .A4(new_n736), .ZN(new_n1049));
  AND2_X1   g863(.A1(new_n930), .A2(new_n767), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n824), .A2(new_n829), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OR2_X1    g866(.A1(new_n852), .A2(new_n861), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1052), .A2(new_n1053), .A3(new_n232), .A4(new_n875), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n300), .A2(new_n328), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n545), .A2(new_n546), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1058), .B1(G900), .B2(G953), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n862), .B1(new_n895), .B2(new_n874), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n930), .A2(new_n754), .A3(new_n767), .ZN(new_n1062));
  INV_X1    g876(.A(KEYINPUT62), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g878(.A1(new_n930), .A2(KEYINPUT62), .A3(new_n754), .A4(new_n767), .ZN(new_n1065));
  INV_X1    g879(.A(new_n818), .ZN(new_n1066));
  INV_X1    g880(.A(new_n943), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n735), .B1(new_n936), .B2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g882(.A1(new_n1064), .A2(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(G953), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g884(.A(new_n1057), .B(KEYINPUT124), .ZN(new_n1071));
  INV_X1    g885(.A(new_n1071), .ZN(new_n1072));
  OAI211_X1 g886(.A(new_n1047), .B(new_n1060), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g887(.A(KEYINPUT126), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n232), .B1(G227), .B2(G900), .ZN(new_n1075));
  INV_X1    g889(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1078));
  NAND2_X1  g892(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1079));
  NAND4_X1  g893(.A1(new_n1053), .A2(new_n1078), .A3(new_n875), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g894(.A1(new_n1080), .A2(new_n232), .ZN(new_n1081));
  AOI22_X1  g895(.A1(new_n1081), .A2(new_n1071), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1082));
  AOI21_X1  g896(.A(KEYINPUT126), .B1(new_n1082), .B2(new_n1047), .ZN(new_n1083));
  OAI211_X1 g897(.A(KEYINPUT126), .B(new_n1060), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1084));
  NAND2_X1  g898(.A1(new_n1084), .A2(new_n1075), .ZN(new_n1085));
  OAI21_X1  g899(.A(new_n1077), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g900(.A(new_n1086), .ZN(G72));
  NAND2_X1  g901(.A1(G472), .A2(G902), .ZN(new_n1088));
  XOR2_X1   g902(.A(new_n1088), .B(KEYINPUT63), .Z(new_n1089));
  OAI21_X1  g903(.A(new_n1089), .B1(new_n1080), .B2(new_n1042), .ZN(new_n1090));
  INV_X1    g904(.A(KEYINPUT127), .ZN(new_n1091));
  OAI21_X1  g905(.A(new_n742), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g906(.A(new_n1092), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  AND3_X1   g907(.A1(new_n1061), .A2(new_n1043), .A3(new_n1052), .ZN(new_n1094));
  INV_X1    g908(.A(new_n1089), .ZN(new_n1095));
  OAI211_X1 g909(.A(new_n340), .B(new_n741), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g910(.A1(new_n384), .A2(new_n386), .ZN(new_n1097));
  AOI21_X1  g911(.A(new_n1095), .B1(new_n1097), .B2(new_n338), .ZN(new_n1098));
  OAI21_X1  g912(.A(new_n1098), .B1(new_n979), .B2(new_n982), .ZN(new_n1099));
  NAND3_X1  g913(.A1(new_n1096), .A2(new_n1025), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g914(.A1(new_n1093), .A2(new_n1100), .ZN(G57));
endmodule


