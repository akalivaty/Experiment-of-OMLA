//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1175, new_n1176,
    new_n1178, new_n1179, new_n1180, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1259, new_n1260;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n206), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G97), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n201), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n219), .B2(new_n220), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n228), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n217), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n252), .A2(G274), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  NOR3_X1   g0057(.A1(new_n256), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n264), .A2(G223), .B1(G77), .B2(new_n262), .ZN(new_n265));
  INV_X1    g0065(.A(G222), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI211_X1 g0069(.A(new_n255), .B(new_n258), .C1(new_n269), .C2(new_n256), .ZN(new_n270));
  INV_X1    g0070(.A(G200), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(KEYINPUT66), .B1(G190), .B2(new_n270), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n274));
  XOR2_X1   g0074(.A(KEYINPUT8), .B(G58), .Z(new_n275));
  NAND2_X1  g0075(.A1(new_n210), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n275), .A2(new_n277), .B1(G150), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n217), .B1(new_n211), .B2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G13), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n284), .A2(new_n210), .A3(G1), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n209), .A2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n283), .B1(G50), .B2(new_n286), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT9), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n273), .B(new_n291), .C1(KEYINPUT66), .C2(new_n272), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n270), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n290), .C1(G169), .C2(new_n270), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT16), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G20), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n250), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT69), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT69), .A2(G33), .ZN(new_n306));
  OAI211_X1 g0106(.A(KEYINPUT73), .B(new_n260), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  OR2_X1    g0108(.A1(KEYINPUT69), .A2(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(KEYINPUT69), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT73), .B1(new_n311), .B2(new_n260), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n300), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT72), .ZN(new_n314));
  AOI21_X1  g0114(.A(G20), .B1(new_n259), .B2(new_n261), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(KEYINPUT7), .ZN(new_n316));
  OAI211_X1 g0116(.A(KEYINPUT72), .B(new_n299), .C1(new_n267), .C2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n202), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G58), .A2(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n203), .A2(new_n205), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G20), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(KEYINPUT71), .A3(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n278), .A2(G159), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n298), .B1(new_n319), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT74), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n309), .A2(KEYINPUT3), .A3(new_n310), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT7), .B1(new_n333), .B2(G20), .ZN(new_n334));
  AOI21_X1  g0134(.A(G20), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n202), .B1(new_n335), .B2(new_n299), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n327), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n281), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(new_n298), .C1(new_n319), .C2(new_n327), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n329), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n287), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n275), .A2(new_n288), .ZN(new_n343));
  INV_X1    g0143(.A(new_n275), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n342), .A2(new_n343), .B1(new_n285), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT76), .Z(new_n351));
  NAND2_X1  g0151(.A1(new_n331), .A2(new_n332), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n257), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G223), .B2(G1698), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n256), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n256), .A2(new_n254), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n255), .B1(G232), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n294), .B2(new_n359), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n348), .A2(new_n349), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT18), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT78), .B1(new_n359), .B2(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n359), .A2(new_n271), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT78), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n356), .A2(new_n358), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n345), .A4(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT17), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n348), .A2(new_n363), .A3(new_n374), .A4(new_n349), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n365), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n278), .A2(G50), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n377), .B1(new_n210), .B2(G68), .C1(new_n222), .C2(new_n276), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n282), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT11), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(KEYINPUT67), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(KEYINPUT67), .ZN(new_n382));
  OR3_X1    g0182(.A1(new_n286), .A2(KEYINPUT12), .A3(G68), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT12), .B1(new_n286), .B2(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n383), .A2(new_n384), .B1(new_n342), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n381), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n255), .B1(G238), .B2(new_n357), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n268), .B2(new_n257), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(G232), .B2(new_n264), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n252), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n393), .A2(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(KEYINPUT13), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(KEYINPUT68), .A2(KEYINPUT14), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n393), .B(KEYINPUT13), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n396), .A2(new_n397), .B1(new_n294), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(G169), .A3(new_n397), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n387), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n398), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n387), .B1(new_n403), .B2(G190), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n271), .B2(new_n403), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NOR3_X1   g0206(.A1(new_n256), .A2(new_n254), .A3(new_n223), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n264), .A2(G238), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n224), .B2(new_n267), .C1(new_n228), .C2(new_n268), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n255), .B(new_n407), .C1(new_n409), .C2(new_n256), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(new_n294), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n285), .A2(new_n222), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n288), .A2(G77), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n414), .A2(new_n276), .B1(new_n210), .B2(new_n222), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n275), .B2(new_n278), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n412), .B1(new_n287), .B2(new_n413), .C1(new_n416), .C2(new_n281), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n410), .B2(G169), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n417), .B1(new_n410), .B2(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n271), .B2(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n297), .A2(new_n376), .A3(new_n406), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n286), .A2(new_n229), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n281), .B(new_n286), .C1(G1), .C2(new_n250), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(new_n229), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT81), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n313), .A2(new_n318), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n430), .A2(KEYINPUT80), .A3(new_n224), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT80), .B1(new_n430), .B2(new_n224), .ZN(new_n432));
  XOR2_X1   g0232(.A(G97), .B(G107), .Z(new_n433));
  NAND2_X1  g0233(.A1(KEYINPUT6), .A2(G97), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n433), .A2(KEYINPUT6), .B1(G107), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n431), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n429), .B1(new_n437), .B2(new_n282), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n252), .A2(G274), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT5), .B(G41), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n253), .A2(G1), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT82), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n256), .B1(new_n441), .B2(new_n440), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G257), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n445), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(G250), .B2(new_n264), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT4), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n263), .A2(G244), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n352), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n256), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n388), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n252), .B1(new_n454), .B2(new_n457), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n462), .A2(new_n448), .A3(new_n449), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n294), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n438), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n460), .A2(new_n369), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n463), .A2(new_n271), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n438), .ZN(new_n470));
  XOR2_X1   g0270(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n471));
  INV_X1    g0271(.A(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(G87), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n352), .A2(new_n472), .A3(G20), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n267), .A2(new_n210), .A3(G87), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT23), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n210), .B2(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n224), .A2(KEYINPUT23), .A3(G20), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n475), .A2(new_n472), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n311), .A2(new_n210), .A3(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n471), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n333), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n483));
  INV_X1    g0283(.A(new_n471), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(new_n480), .A4(new_n479), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n281), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT25), .B1(new_n285), .B2(new_n224), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n285), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n426), .A2(new_n224), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(G250), .A2(G1698), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n230), .B2(G1698), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n333), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n311), .A2(G294), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n252), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n446), .A2(G264), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n444), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n490), .B(new_n500), .C1(new_n369), .C2(new_n499), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n466), .A2(new_n470), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n285), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n427), .A2(G116), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n210), .A2(G116), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n282), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT85), .B1(new_n281), .B2(new_n507), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n452), .B(new_n210), .C1(G33), .C2(new_n229), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT20), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n504), .B(new_n505), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G257), .A2(G1698), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n225), .B2(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n333), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n262), .A2(G303), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n252), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n446), .A2(G270), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n444), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G169), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n505), .A2(new_n504), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n511), .A2(new_n512), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n531), .B2(new_n513), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n532), .B2(new_n524), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n521), .A2(new_n523), .A3(new_n294), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n516), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G200), .B1(new_n521), .B2(new_n523), .ZN(new_n536));
  INV_X1    g0336(.A(new_n521), .ZN(new_n537));
  INV_X1    g0337(.A(new_n523), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(G190), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AND4_X1   g0340(.A1(new_n526), .A2(new_n533), .A3(new_n535), .A4(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G238), .A2(G1698), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n223), .B2(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n331), .A2(new_n332), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n311), .A2(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT84), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n256), .ZN(new_n548));
  INV_X1    g0348(.A(new_n441), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n252), .A2(G250), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT83), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n252), .A2(G274), .A3(new_n441), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n548), .A2(new_n294), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n333), .A2(new_n210), .A3(G68), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n277), .A2(new_n557), .A3(G97), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n473), .B1(new_n390), .B2(new_n210), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n281), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n414), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n286), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n414), .B2(new_n426), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n553), .B1(new_n547), .B2(new_n256), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n555), .B(new_n566), .C1(G169), .C2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n548), .A2(G190), .A3(new_n554), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n426), .A2(new_n473), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n562), .A2(new_n570), .A3(new_n564), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n571), .C1(new_n271), .C2(new_n567), .ZN(new_n572));
  INV_X1    g0372(.A(new_n495), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n573), .A2(new_n294), .A3(new_n444), .A4(new_n496), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n495), .A2(new_n443), .A3(new_n497), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G169), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n576), .A2(new_n490), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n541), .A2(new_n568), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n502), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n424), .A2(new_n579), .ZN(G372));
  NAND2_X1  g0380(.A1(new_n405), .A2(new_n419), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n402), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n582), .A2(new_n373), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n346), .A2(new_n361), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n584), .B(new_n374), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n293), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n296), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n568), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n568), .A2(new_n572), .A3(KEYINPUT87), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n526), .A2(new_n533), .A3(new_n535), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n576), .A2(new_n490), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT87), .B1(new_n568), .B2(new_n572), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n466), .A2(new_n470), .A3(new_n501), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n590), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n568), .A2(new_n572), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n438), .A2(new_n465), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n591), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT26), .B1(new_n466), .B2(new_n600), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n424), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n608), .ZN(G369));
  NAND3_X1  g0409(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n610), .A2(KEYINPUT27), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(KEYINPUT27), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(G213), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G343), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n615), .B1(new_n486), .B2(new_n489), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT88), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT88), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n619), .A2(new_n501), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n617), .B1(new_n621), .B2(new_n594), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n593), .A2(new_n616), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n617), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n532), .A2(new_n616), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n593), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n526), .A2(new_n533), .A3(new_n535), .A4(new_n540), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(G330), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0435(.A(new_n213), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G41), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n559), .A2(new_n473), .A3(new_n503), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n637), .A2(new_n638), .A3(new_n209), .ZN(new_n639));
  INV_X1    g0439(.A(new_n220), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(new_n637), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT28), .Z(new_n642));
  NAND4_X1  g0442(.A1(new_n534), .A2(new_n450), .A3(new_n459), .A4(new_n498), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n548), .A2(new_n554), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT90), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT30), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT30), .ZN(new_n647));
  OAI211_X1 g0447(.A(KEYINPUT90), .B(new_n647), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n294), .B1(new_n521), .B2(new_n523), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n463), .A2(new_n575), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n644), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n646), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n615), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT31), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT91), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(KEYINPUT31), .A3(new_n615), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n645), .A2(KEYINPUT30), .B1(new_n650), .B2(new_n644), .ZN(new_n659));
  AOI211_X1 g0459(.A(new_n654), .B(new_n616), .C1(new_n659), .C2(new_n648), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT31), .B1(new_n652), .B2(new_n615), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT91), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n604), .B1(new_n438), .B2(new_n469), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n600), .A2(new_n629), .A3(new_n594), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n501), .A4(new_n616), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n658), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT29), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n577), .A2(new_n526), .A3(new_n533), .A4(new_n535), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n602), .A2(new_n669), .A3(new_n591), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n568), .B1(new_n670), .B2(new_n502), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n605), .A2(new_n606), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n668), .B(new_n616), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NOR4_X1   g0473(.A1(new_n600), .A2(new_n438), .A3(KEYINPUT26), .A4(new_n465), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n602), .A2(new_n604), .A3(new_n591), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n615), .B1(new_n599), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n673), .B1(new_n677), .B2(new_n668), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n667), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n642), .B1(new_n679), .B2(G1), .ZN(G364));
  XOR2_X1   g0480(.A(new_n631), .B(KEYINPUT92), .Z(new_n681));
  NOR2_X1   g0481(.A1(new_n284), .A2(G20), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n209), .B1(new_n682), .B2(G45), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n637), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n681), .B(new_n686), .C1(G330), .C2(new_n630), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n216), .B1(G20), .B2(new_n388), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT93), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n210), .A2(new_n294), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G200), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n369), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G50), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n210), .A2(G179), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(new_n369), .A3(G200), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n696), .A2(new_n697), .B1(new_n699), .B2(new_n224), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(G190), .A3(G200), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n700), .B1(G87), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G190), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n267), .B1(new_n705), .B2(new_n222), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n693), .A2(G190), .A3(new_n271), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n706), .B1(G58), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n210), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n694), .A2(G190), .ZN(new_n713));
  AOI22_X1  g0513(.A1(G97), .A2(new_n712), .B1(new_n713), .B2(G68), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n698), .A2(new_n704), .ZN(new_n715));
  INV_X1    g0515(.A(G159), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT32), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n703), .A2(new_n709), .A3(new_n714), .A4(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G311), .ZN(new_n720));
  INV_X1    g0520(.A(G329), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n705), .A2(new_n720), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n267), .B(new_n722), .C1(G322), .C2(new_n708), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n701), .B(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G303), .ZN(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT94), .B(G326), .Z(new_n726));
  INV_X1    g0526(.A(new_n699), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n695), .A2(new_n726), .B1(new_n727), .B2(G283), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT33), .B(G317), .ZN(new_n729));
  AOI22_X1  g0529(.A1(G294), .A2(new_n712), .B1(new_n713), .B2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n723), .A2(new_n725), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n692), .B1(new_n719), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G13), .A2(G33), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G20), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n691), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n333), .A2(new_n636), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n640), .A2(new_n253), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(new_n253), .C2(new_n248), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n636), .A2(new_n262), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n741), .A2(G355), .B1(new_n503), .B2(new_n636), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n737), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n732), .A2(new_n743), .A3(new_n686), .ZN(new_n744));
  INV_X1    g0544(.A(new_n735), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n630), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n687), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(G396));
  NOR2_X1   g0548(.A1(new_n691), .A2(new_n733), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n686), .B1(new_n749), .B2(new_n222), .ZN(new_n750));
  INV_X1    g0550(.A(new_n715), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n267), .B1(new_n751), .B2(G311), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n752), .B1(new_n503), .B2(new_n705), .C1(new_n753), .C2(new_n707), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n699), .A2(new_n473), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(G97), .B2(new_n712), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  INV_X1    g0557(.A(new_n713), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n756), .B1(new_n757), .B2(new_n758), .C1(new_n759), .C2(new_n696), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n754), .B(new_n760), .C1(G107), .C2(new_n724), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n712), .A2(G58), .B1(new_n727), .B2(G68), .ZN(new_n762));
  INV_X1    g0562(.A(G132), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n762), .B(new_n333), .C1(new_n763), .C2(new_n715), .ZN(new_n764));
  INV_X1    g0564(.A(new_n705), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n708), .A2(G143), .B1(new_n765), .B2(G159), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  INV_X1    g0567(.A(G150), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n766), .B1(new_n696), .B2(new_n767), .C1(new_n768), .C2(new_n758), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT34), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n764), .B(new_n771), .C1(G50), .C2(new_n724), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n761), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n417), .A2(new_n615), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n422), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n420), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n419), .A2(new_n616), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n750), .B1(new_n692), .B2(new_n774), .C1(new_n780), .C2(new_n734), .ZN(new_n781));
  INV_X1    g0581(.A(new_n607), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n779), .B1(new_n782), .B2(new_n615), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n616), .B(new_n780), .C1(new_n671), .C2(new_n672), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n667), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n686), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n785), .A2(new_n786), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n787), .B2(new_n788), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n781), .B1(new_n790), .B2(new_n792), .ZN(G384));
  AOI211_X1 g0593(.A(new_n503), .B(new_n219), .C1(new_n435), .C2(KEYINPUT35), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(KEYINPUT35), .B2(new_n435), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT36), .Z(new_n796));
  NAND3_X1  g0596(.A1(new_n640), .A2(G77), .A3(new_n320), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n697), .A2(G68), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n209), .B(G13), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n282), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n345), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n613), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT98), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n804), .A2(KEYINPUT98), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n376), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n804), .A2(new_n361), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n341), .A2(new_n345), .A3(new_n371), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT37), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n348), .A2(new_n349), .A3(new_n805), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT37), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n364), .A2(new_n816), .A3(new_n817), .A4(new_n813), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n811), .A2(KEYINPUT38), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT38), .B1(new_n811), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n784), .A2(new_n778), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n387), .A2(new_n615), .ZN(new_n824));
  AND3_X1   g0624(.A1(new_n402), .A2(new_n405), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n402), .B2(new_n405), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT97), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n827), .B1(new_n784), .B2(new_n778), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n586), .A2(new_n613), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n811), .A2(KEYINPUT38), .A3(new_n819), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT101), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n811), .A2(KEYINPUT101), .A3(KEYINPUT38), .A4(new_n819), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n816), .B1(new_n585), .B2(new_n373), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n816), .A2(new_n813), .A3(new_n584), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n818), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n842), .B1(new_n845), .B2(KEYINPUT100), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT100), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n844), .A2(new_n847), .A3(new_n818), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n836), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n820), .A2(new_n821), .A3(new_n836), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n402), .A2(new_n615), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT99), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n834), .B(new_n835), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n588), .B1(new_n678), .B2(new_n424), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n856), .B(new_n857), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n652), .A2(new_n860), .A3(KEYINPUT31), .A4(new_n615), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n665), .A2(new_n859), .A3(new_n861), .A4(new_n655), .ZN(new_n862));
  INV_X1    g0662(.A(new_n826), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n402), .A2(new_n405), .A3(new_n824), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n779), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT40), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n841), .B2(new_n849), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n811), .A2(new_n819), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n866), .B1(new_n872), .B2(new_n837), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(KEYINPUT40), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n424), .A2(new_n862), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(G330), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n858), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n209), .B2(new_n682), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n858), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n800), .B1(new_n880), .B2(new_n881), .ZN(G367));
  XOR2_X1   g0682(.A(new_n637), .B(KEYINPUT41), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n604), .A2(new_n615), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT104), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n663), .B1(new_n438), .B2(new_n616), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n626), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT44), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n626), .A2(new_n888), .ZN(new_n891));
  XOR2_X1   g0691(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n892));
  XNOR2_X1  g0692(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n633), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(KEYINPUT106), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(KEYINPUT106), .ZN(new_n896));
  INV_X1    g0696(.A(new_n681), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n622), .B(new_n623), .ZN(new_n898));
  MUX2_X1   g0698(.A(new_n631), .B(new_n897), .S(new_n898), .Z(new_n899));
  AND2_X1   g0699(.A1(new_n899), .A2(new_n679), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n890), .A2(new_n633), .A3(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n895), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n679), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n884), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n683), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n888), .A2(new_n624), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n888), .A2(new_n594), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n615), .B1(new_n909), .B2(new_n466), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT43), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n571), .A2(new_n616), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n568), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n602), .A2(new_n591), .A3(new_n912), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n908), .A2(new_n910), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n911), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n888), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n633), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n920), .B(new_n922), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n906), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n738), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n241), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n736), .B1(new_n213), .B2(new_n414), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n685), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n267), .B1(new_n699), .B2(new_n222), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT109), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n707), .A2(new_n768), .B1(new_n715), .B2(new_n767), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G50), .B2(new_n765), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n711), .A2(new_n202), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G58), .B2(new_n702), .ZN(new_n934));
  AOI22_X1  g0734(.A1(G143), .A2(new_n695), .B1(new_n713), .B2(G159), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n930), .A2(new_n932), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n712), .A2(G107), .B1(new_n765), .B2(G283), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(KEYINPUT107), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n696), .A2(new_n720), .B1(new_n699), .B2(new_n229), .ZN(new_n939));
  INV_X1    g0739(.A(G317), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n707), .A2(new_n759), .B1(new_n715), .B2(new_n940), .ZN(new_n941));
  NOR4_X1   g0741(.A1(new_n938), .A2(new_n939), .A3(new_n333), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n724), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n701), .A2(new_n503), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(KEYINPUT46), .B2(new_n944), .C1(new_n753), .C2(new_n758), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n942), .B1(KEYINPUT107), .B2(new_n937), .C1(KEYINPUT108), .C2(new_n945), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(KEYINPUT108), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n936), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT47), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n692), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n928), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n916), .B2(new_n745), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n924), .A2(new_n953), .ZN(G387));
  NOR2_X1   g0754(.A1(new_n899), .A2(new_n679), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n900), .A2(new_n955), .A3(G41), .A4(new_n636), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n899), .A2(new_n684), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT110), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n741), .A2(new_n638), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(G107), .B2(new_n213), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n238), .A2(new_n253), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n275), .A2(new_n697), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT50), .Z(new_n963));
  AOI211_X1 g0763(.A(G45), .B(new_n638), .C1(G68), .C2(G77), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n925), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n960), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n685), .B1(new_n966), .B2(new_n737), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n701), .A2(new_n222), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G97), .B2(new_n727), .ZN(new_n969));
  XNOR2_X1  g0769(.A(KEYINPUT111), .B(G150), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n969), .B(new_n333), .C1(new_n715), .C2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT112), .Z(new_n972));
  OAI22_X1  g0772(.A1(new_n707), .A2(new_n697), .B1(new_n705), .B2(new_n202), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(G159), .B2(new_n695), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n563), .A2(new_n712), .B1(new_n713), .B2(new_n275), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n333), .B1(new_n751), .B2(new_n726), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n708), .A2(G317), .B1(new_n765), .B2(G303), .ZN(new_n978));
  INV_X1    g0778(.A(G322), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n696), .B2(new_n979), .C1(new_n720), .C2(new_n758), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT48), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n712), .A2(G283), .B1(new_n702), .B2(G294), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT49), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n977), .B1(new_n503), .B2(new_n699), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n985), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n988), .A2(KEYINPUT49), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n976), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n967), .B1(new_n990), .B2(new_n691), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT113), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n622), .B2(new_n735), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n956), .A2(new_n958), .A3(new_n993), .ZN(G393));
  INV_X1    g0794(.A(new_n901), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n894), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n637), .B1(new_n996), .B2(new_n900), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n903), .A2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n736), .B1(new_n229), .B2(new_n213), .C1(new_n925), .C2(new_n245), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n686), .B1(new_n999), .B2(KEYINPUT114), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n758), .A2(new_n697), .B1(new_n701), .B2(new_n202), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n275), .A2(new_n765), .B1(new_n751), .B2(G143), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n333), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n711), .A2(new_n222), .ZN(new_n1004));
  NOR4_X1   g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n755), .A4(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n696), .A2(new_n768), .B1(new_n716), .B2(new_n707), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT51), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n696), .A2(new_n940), .B1(new_n720), .B2(new_n707), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT52), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n758), .A2(new_n759), .B1(new_n701), .B2(new_n757), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n262), .B1(new_n715), .B2(new_n979), .C1(new_n753), .C2(new_n705), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n711), .A2(new_n503), .B1(new_n699), .B2(new_n224), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1005), .A2(new_n1007), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1000), .B1(KEYINPUT114), .B2(new_n999), .C1(new_n1014), .C2(new_n692), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n921), .B2(new_n735), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n996), .B2(new_n684), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n998), .A2(new_n1017), .ZN(G390));
  NAND3_X1  g0818(.A1(new_n862), .A2(new_n865), .A3(G330), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT115), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT115), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n862), .A2(new_n865), .A3(new_n1021), .A4(G330), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n855), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n832), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n850), .B2(new_n852), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n841), .A2(new_n849), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n778), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n677), .B2(new_n777), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n855), .B1(new_n1029), .B2(new_n827), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1023), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n667), .A2(new_n780), .A3(new_n828), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n855), .B1(new_n1029), .B2(new_n827), .C1(new_n841), .C2(new_n849), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n844), .A2(new_n847), .A3(new_n818), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n847), .B1(new_n844), .B2(new_n818), .ZN(new_n1036));
  NOR3_X1   g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n842), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n839), .B(new_n840), .C1(new_n1037), .C2(KEYINPUT38), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n851), .B1(new_n1038), .B2(new_n836), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1033), .B(new_n1034), .C1(new_n1039), .C2(new_n1025), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1032), .A2(new_n684), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT117), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n424), .A2(G330), .A3(new_n862), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n857), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n828), .B1(new_n667), .B2(new_n780), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n823), .B1(new_n1046), .B2(new_n1023), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT116), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n862), .A2(new_n1048), .A3(G330), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n780), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1048), .B1(new_n862), .B2(G330), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n827), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n1033), .A3(new_n1029), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1045), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1043), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1032), .A2(new_n1040), .A3(new_n1054), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n637), .A3(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n707), .A2(new_n503), .B1(new_n705), .B2(new_n229), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n267), .B(new_n1059), .C1(G294), .C2(new_n751), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n724), .A2(G87), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1004), .B1(G68), .B2(new_n727), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G107), .A2(new_n713), .B1(new_n695), .B2(G283), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  INV_X1    g0865(.A(G125), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n705), .A2(new_n1065), .B1(new_n715), .B2(new_n1066), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n262), .B(new_n1067), .C1(G132), .C2(new_n708), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n701), .A2(new_n970), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT53), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n695), .A2(G128), .B1(new_n727), .B2(G50), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G159), .A2(new_n712), .B1(new_n713), .B2(G137), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n692), .B1(new_n1064), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n686), .B(new_n1074), .C1(new_n344), .C2(new_n749), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1039), .B2(new_n734), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1042), .A2(new_n1058), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(G378));
  INV_X1    g0878(.A(new_n856), .ZN(new_n1079));
  INV_X1    g0879(.A(G330), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n780), .B1(new_n825), .B2(new_n826), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n859), .A2(new_n861), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n661), .B1(new_n579), .B2(new_n616), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n820), .B2(new_n821), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1080), .B1(new_n1085), .B2(new_n867), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT120), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1086), .A2(new_n869), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1086), .B2(new_n869), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n290), .A2(new_n805), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT119), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n297), .B(new_n1091), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1088), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1095), .A2(new_n1086), .A3(new_n1087), .A4(new_n869), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1079), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1084), .A2(KEYINPUT40), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n839), .A2(new_n840), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n846), .A2(new_n848), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n871), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(G330), .B1(new_n873), .B2(KEYINPUT40), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT120), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1086), .A2(new_n869), .A3(new_n1087), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n1108), .A3(new_n1094), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n856), .A3(new_n1097), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1099), .A2(new_n1100), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1109), .A2(KEYINPUT121), .A3(new_n856), .A4(new_n1097), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1111), .A2(new_n684), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1095), .A2(new_n733), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1066), .A2(new_n696), .B1(new_n758), .B2(new_n763), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n708), .A2(G128), .B1(new_n765), .B2(G137), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n701), .B2(new_n1065), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(G150), .C2(new_n712), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n727), .A2(G159), .ZN(new_n1122));
  AOI211_X1 g0922(.A(G33), .B(G41), .C1(new_n751), .C2(G124), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n563), .A2(new_n765), .B1(new_n751), .B2(G283), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n224), .B2(new_n707), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1126), .A2(new_n933), .A3(new_n968), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n696), .A2(new_n503), .B1(new_n699), .B2(new_n201), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G97), .B2(new_n713), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n333), .A2(G41), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT58), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1134));
  AOI211_X1 g0934(.A(G50), .B(new_n1130), .C1(new_n250), .C2(new_n251), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT118), .Z(new_n1136));
  NAND4_X1  g0936(.A1(new_n1124), .A2(new_n1133), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1137), .A2(new_n691), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n686), .B(new_n1138), .C1(new_n697), .C2(new_n749), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1113), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1045), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1057), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1111), .A2(new_n1143), .A3(new_n1112), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1109), .A2(new_n856), .A3(new_n1097), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n856), .B1(new_n1109), .B2(new_n1097), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1143), .B(KEYINPUT57), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1149), .A2(new_n637), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1141), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G375));
  NAND2_X1  g0952(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n827), .A2(new_n733), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n763), .A2(new_n696), .B1(new_n758), .B2(new_n1065), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G50), .B2(new_n712), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n724), .A2(G159), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n707), .A2(new_n767), .B1(new_n715), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G150), .B2(new_n765), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n352), .B1(G58), .B2(new_n727), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n707), .A2(new_n757), .B1(new_n705), .B2(new_n224), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n267), .B(new_n1163), .C1(G303), .C2(new_n751), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n724), .A2(G97), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n712), .A2(new_n563), .B1(new_n727), .B2(G77), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(G116), .A2(new_n713), .B1(new_n695), .B2(G294), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n692), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n686), .B(new_n1169), .C1(new_n202), .C2(new_n749), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1153), .A2(new_n684), .B1(new_n1154), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1055), .A2(new_n884), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1153), .A2(new_n1142), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(G381));
  NOR4_X1   g0974(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1175), .A2(new_n924), .A3(new_n953), .ZN(new_n1176));
  OR4_X1    g0976(.A1(G378), .A2(G375), .A3(new_n1176), .A4(G381), .ZN(G407));
  NAND2_X1  g0977(.A1(new_n614), .A2(G213), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT122), .Z(new_n1179));
  NAND3_X1  g0979(.A1(new_n1151), .A2(new_n1077), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(G407), .A2(G213), .A3(new_n1180), .ZN(G409));
  OR2_X1    g0981(.A1(new_n1144), .A2(new_n883), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n684), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1183), .A2(new_n1140), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G378), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT123), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1151), .B2(G378), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1149), .A2(new_n637), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1145), .B2(new_n1144), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1190), .A2(KEYINPUT123), .A3(new_n1141), .A4(new_n1077), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1186), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1179), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT60), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1173), .B(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n637), .A3(new_n1055), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1171), .ZN(new_n1197));
  INV_X1    g0997(.A(G384), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(G384), .A3(new_n1171), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1192), .A2(KEYINPUT62), .A3(new_n1193), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1141), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(G378), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1151), .A2(new_n1187), .A3(G378), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1178), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1201), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1203), .B1(new_n1211), .B2(KEYINPUT62), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1199), .A2(new_n1200), .B1(G2897), .B2(new_n1179), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1210), .A2(G2897), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1202), .B2(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT127), .B1(new_n1216), .B2(KEYINPUT61), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1215), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1209), .B2(new_n1179), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT127), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1212), .A2(new_n1217), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT124), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G390), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n998), .A2(KEYINPUT124), .A3(new_n1017), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1225), .A2(new_n924), .A3(new_n953), .A4(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(G393), .B(new_n747), .ZN(new_n1228));
  INV_X1    g1028(.A(G387), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1228), .C1(new_n1229), .C2(new_n1225), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT125), .B1(new_n924), .B2(new_n953), .ZN(new_n1231));
  INV_X1    g1031(.A(G390), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1228), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1230), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1223), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1218), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1237), .A2(new_n1221), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT63), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1201), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1192), .A2(new_n1193), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1210), .B1(new_n1246), .B2(new_n1186), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT63), .B1(new_n1247), .B2(new_n1202), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT126), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1237), .A2(new_n1221), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1192), .A2(new_n1178), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1218), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1192), .A2(new_n1178), .A3(new_n1202), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1242), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .A4(new_n1244), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1249), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1239), .A2(new_n1257), .ZN(G405));
  OAI21_X1  g1058(.A(new_n1246), .B1(G378), .B2(new_n1151), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(new_n1202), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(new_n1238), .ZN(G402));
endmodule


