

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n571), .A2(n570), .ZN(n924) );
  INV_X1 U551 ( .A(n683), .ZN(n732) );
  NOR2_X1 U552 ( .A1(n610), .A2(n530), .ZN(n633) );
  NOR2_X2 U553 ( .A1(n569), .A2(n568), .ZN(n571) );
  NOR2_X4 U554 ( .A1(G2104), .A2(n520), .ZN(n901) );
  XOR2_X2 U555 ( .A(KEYINPUT1), .B(n527), .Z(n572) );
  NOR2_X1 U556 ( .A1(n693), .A2(n692), .ZN(n695) );
  INV_X1 U557 ( .A(KEYINPUT17), .ZN(n522) );
  NOR2_X2 U558 ( .A1(n674), .A2(n771), .ZN(n683) );
  XOR2_X1 U559 ( .A(n694), .B(KEYINPUT28), .Z(n515) );
  NOR2_X1 U560 ( .A1(n747), .A2(n765), .ZN(n516) );
  AND2_X1 U561 ( .A1(n896), .A2(G102), .ZN(n517) );
  NAND2_X1 U562 ( .A1(n711), .A2(G1348), .ZN(n696) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n765), .ZN(n726) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n772) );
  XNOR2_X1 U565 ( .A(n580), .B(n579), .ZN(n711) );
  XNOR2_X1 U566 ( .A(n522), .B(KEYINPUT64), .ZN(n523) );
  INV_X1 U567 ( .A(n711), .ZN(n932) );
  XNOR2_X1 U568 ( .A(n524), .B(n523), .ZN(n593) );
  AND2_X1 U569 ( .A1(n526), .A2(n525), .ZN(G164) );
  INV_X1 U570 ( .A(G2105), .ZN(n520) );
  NAND2_X1 U571 ( .A1(G126), .A2(n901), .ZN(n519) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n902) );
  NAND2_X1 U573 ( .A1(G114), .A2(n902), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n519), .A2(n518), .ZN(n521) );
  AND2_X2 U575 ( .A1(n520), .A2(G2104), .ZN(n896) );
  NOR2_X1 U576 ( .A1(n521), .A2(n517), .ZN(n526) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G138), .A2(n593), .ZN(n525) );
  AND2_X1 U579 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X1 U580 ( .A1(G543), .A2(G651), .ZN(n632) );
  NAND2_X1 U581 ( .A1(G91), .A2(n632), .ZN(n529) );
  INV_X1 U582 ( .A(G651), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G543), .A2(n530), .ZN(n527) );
  NAND2_X1 U584 ( .A1(G65), .A2(n572), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n610) );
  NAND2_X1 U587 ( .A1(G78), .A2(n633), .ZN(n532) );
  NOR2_X2 U588 ( .A1(n610), .A2(G651), .ZN(n636) );
  NAND2_X1 U589 ( .A1(G53), .A2(n636), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n925) );
  INV_X1 U592 ( .A(n925), .ZN(G299) );
  INV_X1 U593 ( .A(G108), .ZN(G238) );
  NAND2_X1 U594 ( .A1(G64), .A2(n572), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G52), .A2(n636), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G90), .A2(n632), .ZN(n538) );
  NAND2_X1 U598 ( .A1(G77), .A2(n633), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G101), .A2(n896), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(n542), .Z(n671) );
  NAND2_X1 U604 ( .A1(n593), .A2(G137), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT65), .B(n543), .Z(n673) );
  NAND2_X1 U606 ( .A1(n671), .A2(n673), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G125), .A2(n901), .ZN(n545) );
  NAND2_X1 U608 ( .A1(G113), .A2(n902), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n668) );
  NOR2_X1 U610 ( .A1(n546), .A2(n668), .ZN(G160) );
  NAND2_X1 U611 ( .A1(G63), .A2(n572), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G51), .A2(n636), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT6), .B(n549), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n632), .A2(G89), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G76), .A2(n633), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U619 ( .A(n553), .B(KEYINPUT5), .Z(n554) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT72), .B(n556), .Z(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  XOR2_X1 U623 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n559) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n558) );
  XOR2_X1 U627 ( .A(n559), .B(n558), .Z(n825) );
  NAND2_X1 U628 ( .A1(G567), .A2(n825), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G234) );
  NAND2_X1 U630 ( .A1(G56), .A2(n572), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n562), .Z(n569) );
  NAND2_X1 U632 ( .A1(G81), .A2(n632), .ZN(n563) );
  XOR2_X1 U633 ( .A(KEYINPUT69), .B(n563), .Z(n564) );
  XNOR2_X1 U634 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G68), .A2(n633), .ZN(n565) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NAND2_X1 U638 ( .A1(n636), .A2(G43), .ZN(n570) );
  INV_X1 U639 ( .A(G860), .ZN(n830) );
  OR2_X1 U640 ( .A1(n924), .A2(n830), .ZN(G153) );
  INV_X1 U641 ( .A(G868), .ZN(n650) );
  NOR2_X1 U642 ( .A1(G171), .A2(n650), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G92), .A2(n632), .ZN(n574) );
  NAND2_X1 U644 ( .A1(G66), .A2(n572), .ZN(n573) );
  NAND2_X1 U645 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G79), .A2(n633), .ZN(n576) );
  NAND2_X1 U647 ( .A1(G54), .A2(n636), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U650 ( .A(KEYINPUT70), .B(KEYINPUT15), .ZN(n579) );
  NOR2_X1 U651 ( .A1(G868), .A2(n932), .ZN(n581) );
  NOR2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U653 ( .A(KEYINPUT71), .B(n583), .ZN(G284) );
  XOR2_X1 U654 ( .A(KEYINPUT73), .B(n650), .Z(n584) );
  NOR2_X1 U655 ( .A1(G286), .A2(n584), .ZN(n586) );
  NOR2_X1 U656 ( .A1(G868), .A2(G299), .ZN(n585) );
  NOR2_X1 U657 ( .A1(n586), .A2(n585), .ZN(G297) );
  NAND2_X1 U658 ( .A1(n830), .A2(G559), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n587), .A2(n932), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U661 ( .A1(G868), .A2(n924), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n932), .A2(G868), .ZN(n589) );
  NOR2_X1 U663 ( .A1(G559), .A2(n589), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(G282) );
  NAND2_X1 U665 ( .A1(n901), .A2(G123), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT18), .ZN(n595) );
  BUF_X1 U667 ( .A(n593), .Z(n897) );
  NAND2_X1 U668 ( .A1(G135), .A2(n897), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U670 ( .A(KEYINPUT74), .B(n596), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G99), .A2(n896), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G111), .A2(n902), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n985) );
  XNOR2_X1 U675 ( .A(n985), .B(G2096), .ZN(n601) );
  INV_X1 U676 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U677 ( .A1(n601), .A2(n852), .ZN(G156) );
  NAND2_X1 U678 ( .A1(n633), .A2(G75), .ZN(n602) );
  XOR2_X1 U679 ( .A(KEYINPUT79), .B(n602), .Z(n604) );
  NAND2_X1 U680 ( .A1(n632), .A2(G88), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT80), .B(n605), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G62), .A2(n572), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G50), .A2(n636), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G166) );
  NAND2_X1 U687 ( .A1(G74), .A2(G651), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G87), .A2(n610), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n572), .A2(n613), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G49), .A2(n636), .ZN(n614) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(n614), .Z(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(G288) );
  XOR2_X1 U694 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n618) );
  NAND2_X1 U695 ( .A1(G73), .A2(n633), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n618), .B(n617), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G86), .A2(n632), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G61), .A2(n572), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n636), .A2(G48), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(G305) );
  NAND2_X1 U703 ( .A1(G85), .A2(n632), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G72), .A2(n633), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G47), .A2(n636), .ZN(n627) );
  XOR2_X1 U707 ( .A(KEYINPUT66), .B(n627), .Z(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n572), .A2(G60), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G67), .A2(n572), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G93), .A2(n632), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G80), .A2(n633), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G55), .A2(n636), .ZN(n637) );
  XNOR2_X1 U716 ( .A(KEYINPUT75), .B(n637), .ZN(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(KEYINPUT76), .ZN(n831) );
  XNOR2_X1 U720 ( .A(n831), .B(KEYINPUT19), .ZN(n644) );
  XOR2_X1 U721 ( .A(G305), .B(G299), .Z(n643) );
  XNOR2_X1 U722 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U723 ( .A(n645), .B(G290), .Z(n646) );
  XNOR2_X1 U724 ( .A(G288), .B(n646), .ZN(n647) );
  XNOR2_X1 U725 ( .A(G166), .B(n647), .ZN(n867) );
  NAND2_X1 U726 ( .A1(n932), .A2(G559), .ZN(n648) );
  XOR2_X1 U727 ( .A(n924), .B(n648), .Z(n829) );
  XOR2_X1 U728 ( .A(n867), .B(n829), .Z(n649) );
  NOR2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n652) );
  NOR2_X1 U730 ( .A1(n831), .A2(G868), .ZN(n651) );
  NOR2_X1 U731 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2084), .A2(G2078), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n653), .Z(n654) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n654), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT81), .B(KEYINPUT21), .Z(n655) );
  XNOR2_X1 U736 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G2072), .A2(n657), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U739 ( .A1(G120), .A2(G69), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT83), .B(n658), .Z(n659) );
  NOR2_X1 U741 ( .A1(G238), .A2(n659), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G57), .A2(n660), .ZN(n833) );
  NAND2_X1 U743 ( .A1(n833), .A2(G567), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G132), .A2(G82), .ZN(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(KEYINPUT22), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(KEYINPUT82), .ZN(n663) );
  NOR2_X1 U747 ( .A1(G218), .A2(n663), .ZN(n664) );
  NAND2_X1 U748 ( .A1(G96), .A2(n664), .ZN(n834) );
  NAND2_X1 U749 ( .A1(n834), .A2(G2106), .ZN(n665) );
  NAND2_X1 U750 ( .A1(n666), .A2(n665), .ZN(n845) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n667) );
  NOR2_X1 U752 ( .A1(n845), .A2(n667), .ZN(n828) );
  NAND2_X1 U753 ( .A1(n828), .A2(G36), .ZN(G176) );
  XOR2_X1 U754 ( .A(KEYINPUT84), .B(G166), .Z(G303) );
  INV_X1 U755 ( .A(G171), .ZN(G301) );
  INV_X1 U756 ( .A(n772), .ZN(n674) );
  INV_X1 U757 ( .A(G40), .ZN(n669) );
  NOR2_X1 U758 ( .A1(n669), .A2(n668), .ZN(n670) );
  AND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n771) );
  NAND2_X2 U761 ( .A1(G8), .A2(n732), .ZN(n765) );
  NOR2_X1 U762 ( .A1(G2084), .A2(n732), .ZN(n727) );
  NOR2_X1 U763 ( .A1(n726), .A2(n727), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n675), .A2(G8), .ZN(n678) );
  INV_X1 U765 ( .A(n678), .ZN(n677) );
  INV_X1 U766 ( .A(KEYINPUT30), .ZN(n676) );
  NAND2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n680) );
  NAND2_X1 U768 ( .A1(KEYINPUT30), .A2(n678), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U770 ( .A(KEYINPUT94), .B(n681), .ZN(n682) );
  NOR2_X1 U771 ( .A1(n682), .A2(G168), .ZN(n689) );
  NOR2_X1 U772 ( .A1(n683), .A2(G1961), .ZN(n684) );
  XNOR2_X1 U773 ( .A(n684), .B(KEYINPUT90), .ZN(n687) );
  XNOR2_X1 U774 ( .A(G2078), .B(KEYINPUT25), .ZN(n685) );
  XNOR2_X1 U775 ( .A(n685), .B(KEYINPUT91), .ZN(n1005) );
  NOR2_X1 U776 ( .A1(n732), .A2(n1005), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n687), .A2(n686), .ZN(n719) );
  AND2_X1 U778 ( .A1(G301), .A2(n719), .ZN(n688) );
  NOR2_X1 U779 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U780 ( .A(n690), .B(KEYINPUT31), .ZN(n723) );
  NAND2_X1 U781 ( .A1(n683), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  INV_X1 U783 ( .A(G1956), .ZN(n926) );
  NOR2_X1 U784 ( .A1(n926), .A2(n683), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n695), .A2(n925), .ZN(n694) );
  NAND2_X1 U786 ( .A1(n695), .A2(n925), .ZN(n715) );
  XNOR2_X1 U787 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n696), .A2(n705), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G1341), .A2(n697), .ZN(n698) );
  NOR2_X1 U790 ( .A1(n683), .A2(n698), .ZN(n699) );
  NOR2_X1 U791 ( .A1(n924), .A2(n699), .ZN(n704) );
  NAND2_X1 U792 ( .A1(n711), .A2(G2067), .ZN(n701) );
  NAND2_X1 U793 ( .A1(G1996), .A2(n705), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U795 ( .A1(n702), .A2(n683), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U797 ( .A1(G1996), .A2(n705), .ZN(n706) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n713) );
  NAND2_X1 U799 ( .A1(G1348), .A2(n732), .ZN(n709) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n683), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n515), .A2(n716), .ZN(n718) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(KEYINPUT93), .Z(n717) );
  XNOR2_X1 U807 ( .A(n718), .B(n717), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n719), .A2(G301), .ZN(n720) );
  NOR2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U811 ( .A(n724), .B(KEYINPUT95), .ZN(n731) );
  XOR2_X1 U812 ( .A(n731), .B(KEYINPUT96), .Z(n725) );
  NOR2_X1 U813 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U814 ( .A1(G8), .A2(n727), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n729), .A2(n728), .ZN(n743) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n740) );
  INV_X1 U818 ( .A(G8), .ZN(n738) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n765), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U822 ( .A(KEYINPUT97), .B(n735), .Z(n736) );
  NAND2_X1 U823 ( .A1(G303), .A2(n736), .ZN(n737) );
  OR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U826 ( .A(KEYINPUT32), .B(n741), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n751), .A2(n744), .ZN(n938) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n745) );
  AND2_X1 U832 ( .A1(n938), .A2(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n758), .A2(n746), .ZN(n749) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U835 ( .A(n927), .ZN(n747) );
  OR2_X1 U836 ( .A1(KEYINPUT33), .A2(n516), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U838 ( .A(n750), .B(KEYINPUT98), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n765), .A2(n752), .ZN(n753) );
  XOR2_X1 U841 ( .A(KEYINPUT99), .B(n753), .Z(n754) );
  NOR2_X2 U842 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n756), .B(KEYINPUT100), .ZN(n757) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U845 ( .A1(n757), .A2(n921), .ZN(n769) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n758), .A2(n760), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n765), .A2(n761), .ZN(n762) );
  XNOR2_X1 U850 ( .A(n762), .B(KEYINPUT101), .ZN(n767) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U852 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT102), .ZN(n806) );
  XNOR2_X1 U857 ( .A(G1986), .B(G290), .ZN(n930) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT85), .B(n773), .ZN(n802) );
  INV_X1 U860 ( .A(n802), .ZN(n820) );
  NAND2_X1 U861 ( .A1(n930), .A2(n820), .ZN(n804) );
  XOR2_X1 U862 ( .A(KEYINPUT37), .B(G2067), .Z(n817) );
  NAND2_X1 U863 ( .A1(n896), .A2(G104), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G140), .A2(n897), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U866 ( .A(KEYINPUT34), .B(n776), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G128), .A2(n901), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G116), .A2(n902), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT86), .B(n779), .Z(n780) );
  XNOR2_X1 U871 ( .A(KEYINPUT35), .B(n780), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U873 ( .A(n783), .B(KEYINPUT36), .Z(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT87), .B(n784), .Z(n912) );
  NAND2_X1 U875 ( .A1(n817), .A2(n912), .ZN(n992) );
  NOR2_X1 U876 ( .A1(n802), .A2(n992), .ZN(n785) );
  XNOR2_X1 U877 ( .A(KEYINPUT88), .B(n785), .ZN(n815) );
  NAND2_X1 U878 ( .A1(n896), .A2(G95), .ZN(n787) );
  NAND2_X1 U879 ( .A1(G131), .A2(n897), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G119), .A2(n901), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G107), .A2(n902), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n888) );
  INV_X1 U885 ( .A(G1991), .ZN(n862) );
  NOR2_X1 U886 ( .A1(n888), .A2(n862), .ZN(n801) );
  NAND2_X1 U887 ( .A1(G105), .A2(n896), .ZN(n792) );
  XNOR2_X1 U888 ( .A(n792), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n901), .A2(G129), .ZN(n794) );
  NAND2_X1 U890 ( .A1(G141), .A2(n897), .ZN(n793) );
  NAND2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G117), .A2(n902), .ZN(n795) );
  XNOR2_X1 U893 ( .A(KEYINPUT89), .B(n795), .ZN(n796) );
  NOR2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n889) );
  AND2_X1 U896 ( .A1(n889), .A2(G1996), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n987) );
  NOR2_X1 U898 ( .A1(n987), .A2(n802), .ZN(n811) );
  NOR2_X1 U899 ( .A1(n815), .A2(n811), .ZN(n803) );
  AND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n823) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n889), .ZN(n807) );
  XOR2_X1 U903 ( .A(KEYINPUT103), .B(n807), .Z(n982) );
  AND2_X1 U904 ( .A1(n862), .A2(n888), .ZN(n808) );
  XNOR2_X1 U905 ( .A(KEYINPUT104), .B(n808), .ZN(n989) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n989), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n982), .A2(n812), .ZN(n813) );
  XOR2_X1 U910 ( .A(KEYINPUT39), .B(n813), .Z(n814) );
  NOR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U912 ( .A(KEYINPUT105), .B(n816), .ZN(n819) );
  OR2_X1 U913 ( .A1(n912), .A2(n817), .ZN(n818) );
  XNOR2_X1 U914 ( .A(n818), .B(KEYINPUT106), .ZN(n993) );
  NAND2_X1 U915 ( .A1(n819), .A2(n993), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n825), .ZN(G217) );
  INV_X1 U920 ( .A(n825), .ZN(G223) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n826) );
  NAND2_X1 U922 ( .A1(G661), .A2(n826), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NAND2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(G145) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G82), .ZN(G220) );
  NOR2_X1 U932 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U934 ( .A(G1341), .B(G2454), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n835), .B(G2430), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n836), .B(G1348), .ZN(n842) );
  XOR2_X1 U937 ( .A(G2443), .B(G2427), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2438), .B(G2446), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n840) );
  XOR2_X1 U940 ( .A(G2451), .B(G2435), .Z(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U943 ( .A1(n843), .A2(G14), .ZN(n844) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(n844), .ZN(G401) );
  INV_X1 U945 ( .A(n845), .ZN(G319) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2678), .Z(n847) );
  XNOR2_X1 U947 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2090), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U952 ( .A(n851), .B(n850), .Z(n854) );
  XOR2_X1 U953 ( .A(G2096), .B(n852), .Z(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U955 ( .A(G2084), .B(G2078), .Z(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(G227) );
  XNOR2_X1 U957 ( .A(G1961), .B(n926), .ZN(n858) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1981), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n859), .B(G2474), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1976), .B(G1971), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT41), .B(G1966), .Z(n864) );
  XOR2_X1 U964 ( .A(G1996), .B(n862), .Z(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(G229) );
  XNOR2_X1 U967 ( .A(G286), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n932), .B(G171), .Z(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n870), .B(n924), .ZN(n871) );
  NOR2_X1 U971 ( .A1(G37), .A2(n871), .ZN(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT114), .B(n872), .ZN(G397) );
  NAND2_X1 U973 ( .A1(n901), .A2(G124), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G112), .A2(n902), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n896), .A2(G100), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G136), .A2(n897), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U981 ( .A1(n896), .A2(G103), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G139), .A2(n897), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G127), .A2(n901), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G115), .A2(n902), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(n884), .Z(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n975) );
  XOR2_X1 U990 ( .A(G162), .B(n975), .Z(n891) );
  XOR2_X1 U991 ( .A(n889), .B(n888), .Z(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U993 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  XNOR2_X1 U994 ( .A(G160), .B(KEYINPUT113), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n911) );
  NAND2_X1 U997 ( .A1(n896), .A2(G106), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G142), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(KEYINPUT45), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(G130), .A2(n901), .ZN(n904) );
  NAND2_X1 U1002 ( .A1(G118), .A2(n902), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT111), .B(n905), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(n985), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(G164), .B(n909), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G395) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n917), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G397), .A2(G395), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT115), .B(n918), .Z(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G96), .ZN(G221) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1021 ( .A(G1966), .B(G168), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1023 ( .A(KEYINPUT57), .B(n923), .Z(n946) );
  XOR2_X1 U1024 ( .A(n924), .B(G1341), .Z(n943) );
  XOR2_X1 U1025 ( .A(n926), .B(n925), .Z(n928) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n936) );
  XOR2_X1 U1028 ( .A(G301), .B(G1961), .Z(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT123), .ZN(n934) );
  XOR2_X1 U1030 ( .A(n932), .B(G1348), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(G1971), .A2(G303), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(KEYINPUT124), .B(n941), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT125), .B(n944), .Z(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n948) );
  XOR2_X1 U1040 ( .A(KEYINPUT56), .B(G16), .Z(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(n949), .B(KEYINPUT126), .ZN(n973) );
  XOR2_X1 U1043 ( .A(G1966), .B(G21), .Z(n959) );
  XOR2_X1 U1044 ( .A(G20), .B(G1956), .Z(n953) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1049 ( .A(KEYINPUT59), .B(G1348), .Z(n954) );
  XNOR2_X1 U1050 ( .A(G4), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(n957), .B(KEYINPUT60), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT127), .B(n960), .ZN(n969) );
  XNOR2_X1 U1055 ( .A(G1961), .B(G5), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT61), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n971), .A2(G16), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1004) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(n974), .ZN(n978) );
  XOR2_X1 U1069 ( .A(n975), .B(KEYINPUT117), .Z(n976) );
  XOR2_X1 U1070 ( .A(G2072), .B(n976), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT119), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n980), .B(KEYINPUT50), .ZN(n998) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n983), .Z(n991) );
  XOR2_X1 U1077 ( .A(G2084), .B(G160), .Z(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n995) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1084 ( .A(KEYINPUT116), .B(n996), .Z(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n999), .ZN(n1001) );
  INV_X1 U1087 ( .A(KEYINPUT55), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(G29), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1029) );
  XOR2_X1 U1091 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n1018) );
  XNOR2_X1 U1092 ( .A(n1005), .B(G27), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G2067), .B(G26), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G2072), .B(G33), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT121), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1016) );
  XOR2_X1 U1098 ( .A(G32), .B(G1996), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(G28), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G25), .B(G1991), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(KEYINPUT120), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(G35), .B(G2090), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(G2084), .B(G34), .Z(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT54), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT55), .B(n1024), .Z(n1026) );
  INV_X1 U1111 ( .A(G29), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(G11), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(n1030), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

