

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796;

  BUF_X1 U374 ( .A(n637), .Z(n609) );
  NOR2_X1 U375 ( .A1(n687), .A2(G902), .ZN(n586) );
  INV_X1 U376 ( .A(G902), .ZN(n573) );
  AND2_X1 U377 ( .A1(n511), .A2(n509), .ZN(n508) );
  XNOR2_X1 U378 ( .A(n548), .B(n547), .ZN(n736) );
  AND2_X1 U379 ( .A1(n437), .A2(n436), .ZN(n649) );
  NAND2_X1 U380 ( .A1(n665), .A2(n654), .ZN(n407) );
  XNOR2_X1 U381 ( .A(n435), .B(KEYINPUT39), .ZN(n665) );
  XNOR2_X1 U382 ( .A(n452), .B(KEYINPUT110), .ZN(n418) );
  NAND2_X2 U383 ( .A1(n422), .A2(n419), .ZN(n613) );
  NOR2_X2 U384 ( .A1(n635), .A2(n736), .ZN(n440) );
  XNOR2_X2 U385 ( .A(G143), .B(G128), .ZN(n557) );
  XNOR2_X2 U386 ( .A(n482), .B(n366), .ZN(n795) );
  XNOR2_X2 U387 ( .A(n440), .B(KEYINPUT68), .ZN(n733) );
  XNOR2_X2 U388 ( .A(n609), .B(KEYINPUT6), .ZN(n655) );
  XNOR2_X2 U389 ( .A(n425), .B(n363), .ZN(n596) );
  XNOR2_X2 U390 ( .A(n661), .B(KEYINPUT38), .ZN(n633) );
  XNOR2_X2 U391 ( .A(n586), .B(G472), .ZN(n637) );
  XNOR2_X1 U392 ( .A(G116), .B(G113), .ZN(n522) );
  XNOR2_X1 U393 ( .A(n395), .B(n426), .ZN(n514) );
  NAND2_X1 U394 ( .A1(n418), .A2(n417), .ZN(n601) );
  NAND2_X1 U395 ( .A1(n456), .A2(n454), .ZN(n482) );
  INV_X1 U396 ( .A(n759), .ZN(n455) );
  INV_X1 U397 ( .A(n644), .ZN(n501) );
  XNOR2_X1 U398 ( .A(G110), .B(KEYINPUT82), .ZN(n401) );
  AND2_X2 U399 ( .A1(n672), .A2(n403), .ZN(n766) );
  NAND2_X1 U400 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U401 ( .A1(n396), .A2(n376), .ZN(n395) );
  XNOR2_X1 U402 ( .A(n601), .B(KEYINPUT44), .ZN(n394) );
  AND2_X1 U403 ( .A1(n414), .A2(n485), .ZN(n376) );
  NAND2_X1 U404 ( .A1(n455), .A2(n459), .ZN(n454) );
  AND2_X1 U405 ( .A1(n460), .A2(n457), .ZN(n456) );
  XNOR2_X1 U406 ( .A(n406), .B(n365), .ZN(n411) );
  NOR2_X1 U407 ( .A1(n658), .A2(n661), .ZN(n413) );
  AND2_X1 U408 ( .A1(n470), .A2(n398), .ZN(n381) );
  AND2_X1 U409 ( .A1(n655), .A2(n493), .ZN(n492) );
  AND2_X1 U410 ( .A1(n399), .A2(n400), .ZN(n398) );
  OR2_X1 U411 ( .A1(n472), .A2(KEYINPUT41), .ZN(n400) );
  OR2_X1 U412 ( .A1(n633), .A2(KEYINPUT41), .ZN(n399) );
  XNOR2_X1 U413 ( .A(n441), .B(n595), .ZN(n635) );
  NOR2_X1 U414 ( .A1(n639), .A2(n357), .ZN(n515) );
  XNOR2_X1 U415 ( .A(n486), .B(n556), .ZN(n620) );
  XOR2_X1 U416 ( .A(KEYINPUT62), .B(n687), .Z(n688) );
  XNOR2_X1 U417 ( .A(n585), .B(n584), .ZN(n687) );
  XNOR2_X1 U418 ( .A(n451), .B(n579), .ZN(n585) );
  XNOR2_X1 U419 ( .A(n776), .B(n469), .ZN(n430) );
  XNOR2_X1 U420 ( .A(n370), .B(n587), .ZN(n783) );
  XNOR2_X1 U421 ( .A(n489), .B(KEYINPUT105), .ZN(n488) );
  XNOR2_X1 U422 ( .A(n784), .B(G146), .ZN(n451) );
  XNOR2_X1 U423 ( .A(n524), .B(n523), .ZN(n581) );
  XNOR2_X1 U424 ( .A(n568), .B(n567), .ZN(n784) );
  XNOR2_X1 U425 ( .A(n480), .B(KEYINPUT8), .ZN(n588) );
  XNOR2_X1 U426 ( .A(n438), .B(n549), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n530), .B(n573), .ZN(n668) );
  XNOR2_X1 U428 ( .A(n401), .B(KEYINPUT94), .ZN(n520) );
  XNOR2_X1 U429 ( .A(n557), .B(G134), .ZN(n568) );
  NOR2_X1 U430 ( .A1(n624), .A2(n562), .ZN(n480) );
  XNOR2_X1 U431 ( .A(n522), .B(n521), .ZN(n524) );
  XNOR2_X1 U432 ( .A(KEYINPUT69), .B(KEYINPUT10), .ZN(n439) );
  AND2_X1 U433 ( .A1(n672), .A2(n666), .ZN(n352) );
  XNOR2_X1 U434 ( .A(n581), .B(n505), .ZN(n775) );
  NAND2_X1 U435 ( .A1(n381), .A2(n501), .ZN(n406) );
  XNOR2_X2 U436 ( .A(n407), .B(KEYINPUT40), .ZN(n642) );
  INV_X1 U437 ( .A(KEYINPUT48), .ZN(n426) );
  XNOR2_X1 U438 ( .A(n465), .B(n533), .ZN(n632) );
  XNOR2_X1 U439 ( .A(n443), .B(KEYINPUT81), .ZN(n402) );
  NAND2_X1 U440 ( .A1(n421), .A2(n420), .ZN(n419) );
  AND2_X1 U441 ( .A1(n424), .A2(n423), .ZN(n422) );
  NOR2_X1 U442 ( .A1(n518), .A2(n361), .ZN(n420) );
  XNOR2_X1 U443 ( .A(n555), .B(n554), .ZN(n701) );
  NAND2_X1 U444 ( .A1(n394), .A2(n392), .ZN(n391) );
  XNOR2_X1 U445 ( .A(n367), .B(KEYINPUT89), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n477), .B(G146), .ZN(n549) );
  INV_X1 U447 ( .A(G125), .ZN(n477) );
  OR2_X1 U448 ( .A1(n728), .A2(n450), .ZN(n449) );
  NOR2_X1 U449 ( .A1(n448), .A2(n446), .ZN(n445) );
  NOR2_X1 U450 ( .A1(n716), .A2(n447), .ZN(n446) );
  INV_X1 U451 ( .A(n720), .ZN(n448) );
  INV_X1 U452 ( .A(n654), .ZN(n447) );
  AND2_X1 U453 ( .A1(n491), .A2(n490), .ZN(n576) );
  INV_X1 U454 ( .A(G237), .ZN(n490) );
  XNOR2_X1 U455 ( .A(n590), .B(n353), .ZN(n433) );
  XNOR2_X1 U456 ( .A(n462), .B(KEYINPUT19), .ZN(n643) );
  NOR2_X1 U457 ( .A1(n632), .A2(n746), .ZN(n462) );
  INV_X1 U458 ( .A(KEYINPUT1), .ZN(n429) );
  XNOR2_X1 U459 ( .A(n466), .B(n467), .ZN(n674) );
  XNOR2_X1 U460 ( .A(n468), .B(n528), .ZN(n467) );
  XNOR2_X1 U461 ( .A(n775), .B(n430), .ZN(n466) );
  NAND2_X1 U462 ( .A1(n507), .A2(KEYINPUT88), .ZN(n506) );
  BUF_X2 U463 ( .A(n632), .Z(n661) );
  AND2_X1 U464 ( .A1(n657), .A2(n494), .ZN(n493) );
  NOR2_X1 U465 ( .A1(n357), .A2(n746), .ZN(n494) );
  INV_X1 U466 ( .A(n606), .ZN(n459) );
  NAND2_X1 U467 ( .A1(n613), .A2(n354), .ZN(n425) );
  NAND2_X1 U468 ( .A1(n701), .A2(n573), .ZN(n486) );
  BUF_X1 U469 ( .A(n643), .Z(n484) );
  INV_X1 U470 ( .A(KEYINPUT115), .ZN(n478) );
  NOR2_X1 U471 ( .A1(n766), .A2(n371), .ZN(n410) );
  INV_X1 U472 ( .A(G472), .ZN(n371) );
  NOR2_X1 U473 ( .A1(n766), .A2(n373), .ZN(n409) );
  INV_X1 U474 ( .A(G475), .ZN(n373) );
  INV_X1 U475 ( .A(n766), .ZN(n374) );
  NOR2_X1 U476 ( .A1(n766), .A2(n372), .ZN(n408) );
  INV_X1 U477 ( .A(G210), .ZN(n372) );
  AND2_X1 U478 ( .A1(n500), .A2(n647), .ZN(n498) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT100), .Z(n543) );
  INV_X1 U480 ( .A(KEYINPUT46), .ZN(n427) );
  NOR2_X1 U481 ( .A1(n431), .A2(n739), .ZN(n740) );
  OR2_X1 U482 ( .A1(G237), .A2(G902), .ZN(n534) );
  XOR2_X1 U483 ( .A(G122), .B(G104), .Z(n552) );
  XNOR2_X1 U484 ( .A(G143), .B(G113), .ZN(n551) );
  XNOR2_X1 U485 ( .A(n488), .B(n487), .ZN(n550) );
  XNOR2_X1 U486 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n487) );
  NAND2_X1 U487 ( .A1(n576), .A2(G214), .ZN(n489) );
  XNOR2_X1 U488 ( .A(n439), .B(n481), .ZN(n438) );
  INV_X1 U489 ( .A(G140), .ZN(n481) );
  XNOR2_X1 U490 ( .A(KEYINPUT71), .B(G137), .ZN(n587) );
  XNOR2_X1 U491 ( .A(n504), .B(n527), .ZN(n468) );
  XNOR2_X1 U492 ( .A(n549), .B(n529), .ZN(n504) );
  NOR2_X1 U493 ( .A1(n513), .A2(KEYINPUT88), .ZN(n512) );
  NOR2_X1 U494 ( .A1(n510), .A2(n684), .ZN(n509) );
  NOR2_X1 U495 ( .A1(n663), .A2(n664), .ZN(n510) );
  AND2_X1 U496 ( .A1(n444), .A2(n685), .ZN(n368) );
  NAND2_X1 U497 ( .A1(n795), .A2(KEYINPUT44), .ZN(n369) );
  AND2_X1 U498 ( .A1(n449), .A2(n445), .ZN(n444) );
  NAND2_X1 U499 ( .A1(G234), .A2(G237), .ZN(n535) );
  OR2_X1 U500 ( .A1(n746), .A2(n473), .ZN(n471) );
  NOR2_X1 U501 ( .A1(n474), .A2(n746), .ZN(n472) );
  XNOR2_X1 U502 ( .A(n464), .B(n463), .ZN(n746) );
  INV_X1 U503 ( .A(KEYINPUT96), .ZN(n463) );
  NAND2_X1 U504 ( .A1(n534), .A2(G214), .ZN(n464) );
  XOR2_X1 U505 ( .A(KEYINPUT4), .B(G101), .Z(n580) );
  XOR2_X1 U506 ( .A(KEYINPUT103), .B(KEYINPUT5), .Z(n578) );
  XNOR2_X1 U507 ( .A(G107), .B(G104), .ZN(n519) );
  XNOR2_X1 U508 ( .A(n525), .B(G122), .ZN(n505) );
  XOR2_X1 U509 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n525) );
  XNOR2_X1 U510 ( .A(G122), .B(KEYINPUT106), .ZN(n559) );
  XNOR2_X1 U511 ( .A(G116), .B(G107), .ZN(n558) );
  AND2_X1 U512 ( .A1(n458), .A2(n652), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n615), .A2(n459), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n614), .B(KEYINPUT104), .ZN(n442) );
  INV_X1 U515 ( .A(KEYINPUT109), .ZN(n387) );
  NOR2_X1 U516 ( .A1(n734), .A2(KEYINPUT109), .ZN(n384) );
  XNOR2_X1 U517 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U518 ( .A(n674), .B(n676), .ZN(n677) );
  XOR2_X1 U519 ( .A(KEYINPUT92), .B(n679), .Z(n704) );
  INV_X1 U520 ( .A(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U521 ( .A(n413), .B(KEYINPUT36), .ZN(n412) );
  NAND2_X1 U522 ( .A1(n653), .A2(n652), .ZN(n683) );
  NOR2_X1 U523 ( .A1(n644), .A2(n484), .ZN(n726) );
  INV_X1 U524 ( .A(G953), .ZN(n491) );
  XOR2_X1 U525 ( .A(KEYINPUT24), .B(G128), .Z(n353) );
  NOR2_X1 U526 ( .A1(n736), .A2(n474), .ZN(n354) );
  XOR2_X1 U527 ( .A(n560), .B(n559), .Z(n355) );
  XNOR2_X1 U528 ( .A(n574), .B(G469), .ZN(n356) );
  AND2_X1 U529 ( .A1(n627), .A2(n626), .ZN(n357) );
  AND2_X1 U530 ( .A1(n613), .A2(n606), .ZN(n358) );
  NOR2_X1 U531 ( .A1(n474), .A2(n471), .ZN(n359) );
  OR2_X1 U532 ( .A1(n597), .A2(n387), .ZN(n360) );
  XNOR2_X1 U533 ( .A(KEYINPUT0), .B(KEYINPUT67), .ZN(n361) );
  AND2_X1 U534 ( .A1(n645), .A2(KEYINPUT80), .ZN(n362) );
  XOR2_X1 U535 ( .A(n566), .B(KEYINPUT22), .Z(n363) );
  AND2_X1 U536 ( .A1(n633), .A2(n475), .ZN(n364) );
  XNOR2_X1 U537 ( .A(KEYINPUT116), .B(KEYINPUT42), .ZN(n365) );
  INV_X1 U538 ( .A(n746), .ZN(n475) );
  XOR2_X1 U539 ( .A(KEYINPUT87), .B(KEYINPUT35), .Z(n366) );
  XNOR2_X1 U540 ( .A(n550), .B(n370), .ZN(n555) );
  AND2_X2 U541 ( .A1(n382), .A2(n374), .ZN(n708) );
  NAND2_X1 U542 ( .A1(n608), .A2(n656), .ZN(n685) );
  NAND2_X1 U543 ( .A1(n503), .A2(n362), .ZN(n502) );
  NAND2_X1 U544 ( .A1(n412), .A2(n734), .ZN(n375) );
  NAND2_X1 U545 ( .A1(n412), .A2(n734), .ZN(n485) );
  INV_X1 U546 ( .A(n609), .ZN(n431) );
  NAND2_X1 U547 ( .A1(n783), .A2(n432), .ZN(n379) );
  NAND2_X1 U548 ( .A1(n377), .A2(n378), .ZN(n380) );
  NAND2_X1 U549 ( .A1(n379), .A2(n380), .ZN(n591) );
  INV_X1 U550 ( .A(n783), .ZN(n377) );
  INV_X1 U551 ( .A(n432), .ZN(n378) );
  XNOR2_X1 U552 ( .A(n434), .B(n433), .ZN(n432) );
  AND2_X1 U553 ( .A1(n749), .A2(n495), .ZN(n500) );
  XNOR2_X1 U554 ( .A(n415), .B(KEYINPUT79), .ZN(n414) );
  NAND2_X1 U555 ( .A1(n591), .A2(n573), .ZN(n441) );
  XNOR2_X1 U556 ( .A(n397), .B(n427), .ZN(n396) );
  NOR2_X1 U557 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U558 ( .A1(n382), .A2(n410), .ZN(n689) );
  NAND2_X1 U559 ( .A1(n382), .A2(n408), .ZN(n678) );
  NAND2_X1 U560 ( .A1(n382), .A2(n409), .ZN(n703) );
  NAND2_X2 U561 ( .A1(n453), .A2(n671), .ZN(n382) );
  NAND2_X1 U562 ( .A1(n385), .A2(n597), .ZN(n607) );
  NAND2_X1 U563 ( .A1(n386), .A2(n383), .ZN(n389) );
  NAND2_X1 U564 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U565 ( .A(n596), .ZN(n385) );
  AND2_X1 U566 ( .A1(n388), .A2(n360), .ZN(n386) );
  NAND2_X1 U567 ( .A1(n596), .A2(KEYINPUT109), .ZN(n388) );
  NAND2_X1 U568 ( .A1(n389), .A2(n517), .ZN(n452) );
  NAND2_X1 U569 ( .A1(n391), .A2(n390), .ZN(n405) );
  NAND2_X1 U570 ( .A1(n393), .A2(n795), .ZN(n392) );
  INV_X1 U571 ( .A(n601), .ZN(n393) );
  NAND2_X1 U572 ( .A1(n642), .A2(n411), .ZN(n397) );
  NAND2_X1 U573 ( .A1(n402), .A2(n431), .ZN(n614) );
  XNOR2_X1 U574 ( .A(n402), .B(n603), .ZN(n604) );
  NOR2_X1 U575 ( .A1(n673), .A2(n404), .ZN(n403) );
  XNOR2_X2 U576 ( .A(n405), .B(KEYINPUT45), .ZN(n672) );
  OR2_X1 U577 ( .A1(n633), .A2(n475), .ZN(n748) );
  NAND2_X1 U578 ( .A1(n359), .A2(n633), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n411), .B(G137), .ZN(G39) );
  NAND2_X1 U580 ( .A1(n416), .A2(n683), .ZN(n415) );
  NAND2_X1 U581 ( .A1(n499), .A2(n497), .ZN(n416) );
  INV_X1 U582 ( .A(n796), .ZN(n417) );
  XNOR2_X1 U583 ( .A(n418), .B(G110), .ZN(G12) );
  NAND2_X1 U584 ( .A1(n643), .A2(n361), .ZN(n424) );
  INV_X1 U585 ( .A(n643), .ZN(n421) );
  NAND2_X1 U586 ( .A1(n518), .A2(n361), .ZN(n423) );
  NAND2_X1 U587 ( .A1(n421), .A2(n749), .ZN(n503) );
  XNOR2_X1 U588 ( .A(n428), .B(n355), .ZN(n564) );
  XNOR2_X1 U589 ( .A(n568), .B(n561), .ZN(n428) );
  XNOR2_X1 U590 ( .A(n639), .B(n429), .ZN(n602) );
  XNOR2_X2 U591 ( .A(n575), .B(n356), .ZN(n639) );
  XNOR2_X1 U592 ( .A(n430), .B(n572), .ZN(n461) );
  XNOR2_X1 U593 ( .A(n663), .B(G140), .ZN(G42) );
  NAND2_X1 U594 ( .A1(n662), .A2(n661), .ZN(n663) );
  INV_X1 U595 ( .A(n591), .ZN(n692) );
  NAND2_X1 U596 ( .A1(n588), .A2(G221), .ZN(n434) );
  NAND2_X1 U597 ( .A1(n649), .A2(n633), .ZN(n435) );
  XNOR2_X1 U598 ( .A(n631), .B(n630), .ZN(n436) );
  XNOR2_X1 U599 ( .A(n629), .B(n628), .ZN(n437) );
  NOR2_X1 U600 ( .A1(n442), .A2(n615), .ZN(n616) );
  NAND2_X1 U601 ( .A1(n742), .A2(n442), .ZN(n743) );
  NAND2_X1 U602 ( .A1(n602), .A2(n733), .ZN(n443) );
  OR2_X1 U603 ( .A1(n728), .A2(n611), .ZN(n731) );
  NOR2_X1 U604 ( .A1(n722), .A2(n654), .ZN(n450) );
  XNOR2_X1 U605 ( .A(n451), .B(n461), .ZN(n711) );
  NAND2_X1 U606 ( .A1(n352), .A2(n667), .ZN(n453) );
  NOR2_X1 U607 ( .A1(n484), .A2(n362), .ZN(n495) );
  NAND2_X1 U608 ( .A1(n759), .A2(n358), .ZN(n460) );
  XNOR2_X2 U609 ( .A(n605), .B(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U610 ( .A1(n674), .A2(n668), .ZN(n465) );
  XNOR2_X1 U611 ( .A(n580), .B(KEYINPUT74), .ZN(n469) );
  INV_X1 U612 ( .A(KEYINPUT41), .ZN(n473) );
  INV_X1 U613 ( .A(n747), .ZN(n474) );
  XNOR2_X2 U614 ( .A(n622), .B(n621), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n476), .A2(n475), .ZN(n631) );
  INV_X1 U616 ( .A(n637), .ZN(n476) );
  NAND2_X1 U617 ( .A1(n725), .A2(n492), .ZN(n658) );
  XNOR2_X2 U618 ( .A(n479), .B(n478), .ZN(n644) );
  NAND2_X1 U619 ( .A1(n641), .A2(n640), .ZN(n479) );
  NAND2_X1 U620 ( .A1(n498), .A2(n501), .ZN(n497) );
  NAND2_X2 U621 ( .A1(n508), .A2(n506), .ZN(n673) );
  NAND2_X1 U622 ( .A1(n483), .A2(n647), .ZN(n499) );
  NAND2_X1 U623 ( .A1(n496), .A2(n502), .ZN(n483) );
  XNOR2_X1 U624 ( .A(n375), .B(n732), .ZN(G27) );
  NAND2_X1 U625 ( .A1(n619), .A2(n620), .ZN(n622) );
  NAND2_X1 U626 ( .A1(n644), .A2(n362), .ZN(n496) );
  INV_X1 U627 ( .A(n514), .ZN(n507) );
  NAND2_X1 U628 ( .A1(n514), .A2(n512), .ZN(n511) );
  INV_X1 U629 ( .A(n663), .ZN(n513) );
  INV_X1 U630 ( .A(n642), .ZN(n686) );
  NAND2_X1 U631 ( .A1(n515), .A2(n733), .ZN(n629) );
  AND2_X1 U632 ( .A1(n733), .A2(n640), .ZN(n516) );
  NAND2_X1 U633 ( .A1(n516), .A2(n722), .ZN(n612) );
  NAND2_X1 U634 ( .A1(n618), .A2(n516), .ZN(n716) );
  INV_X1 U635 ( .A(n557), .ZN(n526) );
  AND2_X1 U636 ( .A1(n609), .A2(n737), .ZN(n517) );
  XNOR2_X1 U637 ( .A(KEYINPUT99), .B(n542), .ZN(n518) );
  INV_X1 U638 ( .A(n668), .ZN(n666) );
  INV_X1 U639 ( .A(KEYINPUT111), .ZN(n603) );
  INV_X1 U640 ( .A(KEYINPUT88), .ZN(n664) );
  INV_X1 U641 ( .A(n656), .ZN(n737) );
  INV_X1 U642 ( .A(KEYINPUT56), .ZN(n681) );
  XNOR2_X2 U643 ( .A(n520), .B(n519), .ZN(n776) );
  INV_X1 U644 ( .A(KEYINPUT3), .ZN(n521) );
  XOR2_X1 U645 ( .A(KEYINPUT73), .B(G119), .Z(n523) );
  XOR2_X1 U646 ( .A(n526), .B(KEYINPUT18), .Z(n528) );
  XNOR2_X2 U647 ( .A(KEYINPUT64), .B(G953), .ZN(n624) );
  INV_X1 U648 ( .A(n624), .ZN(n790) );
  NAND2_X1 U649 ( .A1(n790), .A2(G224), .ZN(n527) );
  XNOR2_X1 U650 ( .A(KEYINPUT17), .B(KEYINPUT91), .ZN(n529) );
  XNOR2_X1 U651 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n530) );
  NAND2_X1 U652 ( .A1(G210), .A2(n534), .ZN(n532) );
  INV_X1 U653 ( .A(KEYINPUT95), .ZN(n531) );
  XNOR2_X1 U654 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U655 ( .A(n535), .B(KEYINPUT14), .ZN(n539) );
  NAND2_X1 U656 ( .A1(G952), .A2(n539), .ZN(n536) );
  XOR2_X1 U657 ( .A(KEYINPUT97), .B(n536), .Z(n758) );
  NOR2_X1 U658 ( .A1(G953), .A2(n758), .ZN(n538) );
  INV_X1 U659 ( .A(KEYINPUT98), .ZN(n537) );
  XNOR2_X1 U660 ( .A(n538), .B(n537), .ZN(n627) );
  NAND2_X1 U661 ( .A1(G902), .A2(n539), .ZN(n623) );
  INV_X1 U662 ( .A(n623), .ZN(n540) );
  NOR2_X1 U663 ( .A1(G898), .A2(n491), .ZN(n780) );
  NAND2_X1 U664 ( .A1(n540), .A2(n780), .ZN(n541) );
  NAND2_X1 U665 ( .A1(n627), .A2(n541), .ZN(n542) );
  NAND2_X1 U666 ( .A1(n668), .A2(G234), .ZN(n544) );
  XNOR2_X1 U667 ( .A(n544), .B(n543), .ZN(n592) );
  INV_X1 U668 ( .A(G221), .ZN(n545) );
  OR2_X1 U669 ( .A1(n592), .A2(n545), .ZN(n548) );
  INV_X1 U670 ( .A(KEYINPUT101), .ZN(n546) );
  XNOR2_X1 U671 ( .A(n546), .B(KEYINPUT21), .ZN(n547) );
  XOR2_X1 U672 ( .A(KEYINPUT70), .B(G131), .Z(n567) );
  XNOR2_X1 U673 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U674 ( .A(n567), .B(n553), .ZN(n554) );
  XOR2_X1 U675 ( .A(KEYINPUT13), .B(G475), .Z(n556) );
  XNOR2_X1 U676 ( .A(n558), .B(KEYINPUT9), .ZN(n561) );
  XOR2_X1 U677 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n560) );
  INV_X1 U678 ( .A(G234), .ZN(n562) );
  NAND2_X1 U679 ( .A1(n588), .A2(G217), .ZN(n563) );
  XNOR2_X1 U680 ( .A(n564), .B(n563), .ZN(n696) );
  NAND2_X1 U681 ( .A1(n696), .A2(n573), .ZN(n565) );
  XNOR2_X1 U682 ( .A(n565), .B(G478), .ZN(n610) );
  NOR2_X1 U683 ( .A1(n620), .A2(n610), .ZN(n747) );
  XNOR2_X1 U684 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n566) );
  XNOR2_X1 U685 ( .A(n587), .B(G140), .ZN(n571) );
  INV_X1 U686 ( .A(G227), .ZN(n569) );
  NOR2_X1 U687 ( .A1(n624), .A2(n569), .ZN(n570) );
  XNOR2_X1 U688 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U689 ( .A1(n711), .A2(n573), .ZN(n575) );
  INV_X1 U690 ( .A(KEYINPUT72), .ZN(n574) );
  INV_X1 U691 ( .A(n602), .ZN(n597) );
  INV_X1 U692 ( .A(n597), .ZN(n734) );
  NAND2_X1 U693 ( .A1(n576), .A2(G210), .ZN(n577) );
  XNOR2_X1 U694 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U695 ( .A(KEYINPUT102), .B(n580), .Z(n583) );
  XNOR2_X1 U696 ( .A(n581), .B(G137), .ZN(n582) );
  XNOR2_X1 U697 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U698 ( .A(G119), .B(G110), .ZN(n589) );
  XNOR2_X1 U699 ( .A(n589), .B(KEYINPUT23), .ZN(n590) );
  INV_X1 U700 ( .A(n592), .ZN(n593) );
  NAND2_X1 U701 ( .A1(n593), .A2(G217), .ZN(n594) );
  XNOR2_X1 U702 ( .A(n594), .B(KEYINPUT25), .ZN(n595) );
  INV_X1 U703 ( .A(n635), .ZN(n656) );
  NOR2_X1 U704 ( .A1(n655), .A2(n596), .ZN(n599) );
  NOR2_X1 U705 ( .A1(n597), .A2(n656), .ZN(n598) );
  NAND2_X1 U706 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U707 ( .A(KEYINPUT32), .B(n600), .Z(n796) );
  AND2_X1 U708 ( .A1(n610), .A2(n620), .ZN(n652) );
  NAND2_X1 U709 ( .A1(n604), .A2(n655), .ZN(n605) );
  XNOR2_X1 U710 ( .A(KEYINPUT34), .B(KEYINPUT75), .ZN(n606) );
  NOR2_X1 U711 ( .A1(n607), .A2(n655), .ZN(n608) );
  NAND2_X1 U712 ( .A1(n609), .A2(n613), .ZN(n617) );
  INV_X1 U713 ( .A(n610), .ZN(n619) );
  OR2_X1 U714 ( .A1(n620), .A2(n619), .ZN(n611) );
  INV_X1 U715 ( .A(n611), .ZN(n722) );
  OR2_X1 U716 ( .A1(n617), .A2(n612), .ZN(n720) );
  INV_X1 U717 ( .A(n613), .ZN(n615) );
  XNOR2_X1 U718 ( .A(KEYINPUT31), .B(n616), .ZN(n728) );
  INV_X1 U719 ( .A(n617), .ZN(n618) );
  INV_X1 U720 ( .A(KEYINPUT108), .ZN(n621) );
  INV_X1 U721 ( .A(n672), .ZN(n764) );
  NOR2_X1 U722 ( .A1(G900), .A2(n623), .ZN(n625) );
  NAND2_X1 U723 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U724 ( .A(KEYINPUT84), .ZN(n628) );
  XNOR2_X1 U725 ( .A(KEYINPUT113), .B(KEYINPUT30), .ZN(n630) );
  NOR2_X1 U726 ( .A1(n357), .A2(n736), .ZN(n634) );
  NAND2_X1 U727 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U728 ( .A(n638), .B(KEYINPUT28), .ZN(n641) );
  INV_X1 U729 ( .A(n639), .ZN(n640) );
  OR2_X1 U730 ( .A1(n654), .A2(n722), .ZN(n749) );
  INV_X1 U731 ( .A(KEYINPUT47), .ZN(n645) );
  INV_X1 U732 ( .A(KEYINPUT80), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n646), .A2(KEYINPUT47), .ZN(n647) );
  INV_X1 U734 ( .A(n661), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U736 ( .A(KEYINPUT114), .ZN(n650) );
  XNOR2_X1 U737 ( .A(n651), .B(n650), .ZN(n653) );
  XNOR2_X1 U738 ( .A(n654), .B(KEYINPUT112), .ZN(n725) );
  NOR2_X1 U739 ( .A1(n656), .A2(n736), .ZN(n657) );
  NOR2_X1 U740 ( .A1(n658), .A2(n734), .ZN(n660) );
  INV_X1 U741 ( .A(KEYINPUT43), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n660), .B(n659), .ZN(n662) );
  AND2_X1 U743 ( .A1(n665), .A2(n722), .ZN(n684) );
  XNOR2_X2 U744 ( .A(n673), .B(KEYINPUT86), .ZN(n763) );
  XNOR2_X1 U745 ( .A(n763), .B(KEYINPUT83), .ZN(n667) );
  XNOR2_X1 U746 ( .A(n668), .B(KEYINPUT85), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n669), .A2(KEYINPUT2), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT66), .ZN(n671) );
  XOR2_X1 U749 ( .A(KEYINPUT90), .B(KEYINPUT54), .Z(n675) );
  XNOR2_X1 U750 ( .A(n675), .B(KEYINPUT55), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n678), .B(n677), .ZN(n680) );
  NOR2_X1 U752 ( .A1(n790), .A2(G952), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n680), .A2(n704), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(n681), .ZN(G51) );
  XNOR2_X1 U755 ( .A(n683), .B(G143), .ZN(G45) );
  XOR2_X1 U756 ( .A(G134), .B(n684), .Z(G36) );
  XNOR2_X1 U757 ( .A(n685), .B(G101), .ZN(G3) );
  XOR2_X1 U758 ( .A(G131), .B(n686), .Z(G33) );
  XNOR2_X1 U759 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n690), .A2(n704), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n691), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U762 ( .A1(n708), .A2(G217), .ZN(n694) );
  XOR2_X1 U763 ( .A(KEYINPUT123), .B(n692), .Z(n693) );
  XNOR2_X1 U764 ( .A(n694), .B(n693), .ZN(n695) );
  INV_X1 U765 ( .A(n704), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n695), .A2(n714), .ZN(G66) );
  NAND2_X1 U767 ( .A1(n708), .A2(G478), .ZN(n698) );
  XOR2_X1 U768 ( .A(n696), .B(KEYINPUT122), .Z(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U770 ( .A1(n699), .A2(n714), .ZN(G63) );
  XNOR2_X1 U771 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n707) );
  XNOR2_X1 U774 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n707), .B(n706), .ZN(G60) );
  NAND2_X1 U776 ( .A1(n708), .A2(G469), .ZN(n713) );
  XNOR2_X1 U777 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n709) );
  XNOR2_X1 U778 ( .A(n709), .B(KEYINPUT58), .ZN(n710) );
  XNOR2_X1 U779 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U780 ( .A(n713), .B(n712), .ZN(n715) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(G54) );
  INV_X1 U782 ( .A(n725), .ZN(n729) );
  NOR2_X1 U783 ( .A1(n716), .A2(n729), .ZN(n718) );
  XNOR2_X1 U784 ( .A(G104), .B(KEYINPUT117), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n718), .B(n717), .ZN(G6) );
  XOR2_X1 U786 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n719) );
  XNOR2_X1 U787 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U788 ( .A(G107), .B(n721), .ZN(G9) );
  XOR2_X1 U789 ( .A(G128), .B(KEYINPUT29), .Z(n724) );
  NAND2_X1 U790 ( .A1(n726), .A2(n722), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n724), .B(n723), .ZN(G30) );
  NAND2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U793 ( .A(n727), .B(G146), .ZN(G48) );
  NOR2_X1 U794 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U795 ( .A(G113), .B(n730), .Z(G15) );
  XNOR2_X1 U796 ( .A(G116), .B(n731), .ZN(G18) );
  XOR2_X1 U797 ( .A(G125), .B(KEYINPUT37), .Z(n732) );
  NOR2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U799 ( .A(KEYINPUT50), .B(n735), .Z(n741) );
  NAND2_X1 U800 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U801 ( .A(n738), .B(KEYINPUT49), .ZN(n739) );
  NAND2_X1 U802 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U803 ( .A(KEYINPUT118), .B(n743), .Z(n744) );
  XNOR2_X1 U804 ( .A(KEYINPUT51), .B(n744), .ZN(n745) );
  NAND2_X1 U805 ( .A1(n381), .A2(n745), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n748), .A2(n747), .ZN(n752) );
  NAND2_X1 U807 ( .A1(n364), .A2(n749), .ZN(n750) );
  XOR2_X1 U808 ( .A(KEYINPUT119), .B(n750), .Z(n751) );
  NAND2_X1 U809 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U810 ( .A1(n759), .A2(n753), .ZN(n754) );
  NAND2_X1 U811 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U812 ( .A(KEYINPUT52), .B(n756), .Z(n757) );
  NOR2_X1 U813 ( .A1(n758), .A2(n757), .ZN(n761) );
  AND2_X1 U814 ( .A1(n759), .A2(n381), .ZN(n760) );
  NOR2_X1 U815 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U816 ( .A1(n762), .A2(n491), .ZN(n769) );
  NOR2_X1 U817 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U818 ( .A1(n765), .A2(KEYINPUT2), .ZN(n767) );
  NOR2_X1 U819 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U820 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n770), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U822 ( .A1(n491), .A2(n672), .ZN(n774) );
  NAND2_X1 U823 ( .A1(G953), .A2(G224), .ZN(n771) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n771), .ZN(n772) );
  NAND2_X1 U825 ( .A1(n772), .A2(G898), .ZN(n773) );
  NAND2_X1 U826 ( .A1(n774), .A2(n773), .ZN(n782) );
  XNOR2_X1 U827 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U828 ( .A(n777), .B(KEYINPUT124), .ZN(n778) );
  XNOR2_X1 U829 ( .A(n778), .B(G101), .ZN(n779) );
  NOR2_X1 U830 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U831 ( .A(n782), .B(n781), .ZN(G69) );
  XNOR2_X1 U832 ( .A(n783), .B(KEYINPUT125), .ZN(n786) );
  XNOR2_X1 U833 ( .A(n784), .B(KEYINPUT4), .ZN(n785) );
  XNOR2_X1 U834 ( .A(n786), .B(n785), .ZN(n789) );
  XOR2_X1 U835 ( .A(G227), .B(n789), .Z(n787) );
  NAND2_X1 U836 ( .A1(n787), .A2(G900), .ZN(n788) );
  NAND2_X1 U837 ( .A1(n788), .A2(G953), .ZN(n794) );
  XOR2_X1 U838 ( .A(n763), .B(n789), .Z(n791) );
  NAND2_X1 U839 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U840 ( .A(n792), .B(KEYINPUT126), .ZN(n793) );
  NAND2_X1 U841 ( .A1(n794), .A2(n793), .ZN(G72) );
  XOR2_X1 U842 ( .A(n795), .B(G122), .Z(G24) );
  XOR2_X1 U843 ( .A(G119), .B(n796), .Z(G21) );
endmodule

