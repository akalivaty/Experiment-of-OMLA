//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G97), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n225), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  AND3_X1   g0046(.A1(new_n205), .A2(KEYINPUT66), .A3(G20), .ZN(new_n247));
  AOI21_X1  g0047(.A(KEYINPUT66), .B1(new_n205), .B2(G20), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n206), .A3(G1), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n214), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n251), .A2(new_n256), .B1(new_n253), .B2(new_n250), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT73), .ZN(new_n258));
  AND3_X1   g0058(.A1(KEYINPUT71), .A2(G58), .A3(G68), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT71), .B1(G58), .B2(G68), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G58), .A2(G68), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G159), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n206), .A2(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n262), .A2(new_n206), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT70), .B(KEYINPUT3), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n264), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n266), .B1(new_n276), .B2(G68), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n258), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n264), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n275), .B1(new_n282), .B2(new_n271), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n271), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT7), .B1(new_n285), .B2(new_n206), .ZN(new_n286));
  OAI21_X1  g0086(.A(G68), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n265), .A2(new_n263), .ZN(new_n288));
  OR3_X1    g0088(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n278), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(KEYINPUT73), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n279), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n255), .ZN(new_n295));
  INV_X1    g0095(.A(G68), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n280), .A2(new_n281), .A3(new_n264), .ZN(new_n297));
  INV_X1    g0097(.A(new_n284), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n206), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n296), .B1(new_n299), .B2(KEYINPUT7), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n270), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(G33), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(G20), .B1(new_n304), .B2(new_n284), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n267), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n266), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n295), .B1(new_n307), .B2(KEYINPUT16), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n294), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT74), .B1(new_n294), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n257), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G41), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(G1), .A3(G13), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n280), .A2(new_n281), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n298), .B1(new_n314), .B2(G33), .ZN(new_n315));
  MUX2_X1   g0115(.A(G223), .B(G226), .S(G1698), .Z(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G87), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G274), .ZN(new_n320));
  AND2_X1   g0120(.A1(G1), .A2(G13), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n312), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n323), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n225), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G179), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT75), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n319), .B2(new_n327), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n311), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT18), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n328), .A2(G200), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n319), .A2(KEYINPUT76), .A3(G190), .A4(new_n327), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n328), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT76), .B1(new_n340), .B2(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n257), .B(new_n342), .C1(new_n309), .C2(new_n310), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n257), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT74), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT73), .B1(new_n291), .B2(new_n292), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n258), .B(new_n278), .C1(new_n287), .C2(new_n290), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n306), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n305), .B2(new_n267), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n290), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n255), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n347), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n294), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n346), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT17), .A3(new_n342), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n311), .A2(new_n360), .A3(new_n334), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n336), .A2(new_n345), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n268), .A2(G222), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n268), .A2(G1698), .ZN(new_n366));
  INV_X1    g0166(.A(G223), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n365), .B1(new_n218), .B2(new_n268), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n313), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n325), .ZN(new_n371));
  INV_X1    g0171(.A(new_n326), .ZN(new_n372));
  XNOR2_X1  g0172(.A(KEYINPUT65), .B(G226), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G169), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n253), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n295), .ZN(new_n379));
  INV_X1    g0179(.A(G50), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n249), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n380), .B2(new_n253), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n206), .A2(G33), .ZN(new_n383));
  INV_X1    g0183(.A(G150), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n250), .A2(new_n383), .B1(new_n384), .B2(new_n265), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G50), .A2(G58), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n206), .B1(new_n386), .B2(new_n296), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n255), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n377), .B(new_n389), .C1(G179), .C2(new_n375), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n389), .B(KEYINPUT9), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n375), .A2(G200), .ZN(new_n393));
  INV_X1    g0193(.A(new_n375), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT10), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT10), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n392), .A2(new_n398), .A3(new_n393), .A4(new_n395), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n253), .A2(new_n296), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT12), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n296), .A2(G20), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n403), .B1(new_n383), .B2(new_n218), .C1(new_n380), .C2(new_n265), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n404), .A2(new_n255), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n402), .B1(KEYINPUT11), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(KEYINPUT11), .B2(new_n405), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n379), .A2(new_n249), .A3(new_n296), .ZN(new_n408));
  XOR2_X1   g0208(.A(new_n408), .B(KEYINPUT69), .Z(new_n409));
  OR2_X1    g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n225), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n268), .B(new_n411), .C1(G226), .C2(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n313), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G238), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n325), .B1(new_n415), .B2(new_n326), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n414), .A2(KEYINPUT13), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT13), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(G169), .ZN(new_n421));
  INV_X1    g0221(.A(G179), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(new_n419), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n419), .B2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n410), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n407), .A2(new_n409), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n419), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(G190), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n427), .C1(new_n428), .C2(new_n419), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n431), .A2(new_n383), .B1(new_n206), .B2(new_n218), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n250), .A2(new_n265), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n255), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G77), .B1(new_n247), .B2(new_n248), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n434), .B1(G77), .B2(new_n378), .C1(new_n379), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT67), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G107), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n366), .A2(new_n415), .B1(new_n440), .B2(new_n268), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n285), .A2(new_n225), .A3(G1698), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n369), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n371), .B1(G244), .B2(new_n372), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT68), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n436), .B1(new_n446), .B2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT68), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n445), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G190), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n376), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n422), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n436), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n400), .A2(new_n430), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n363), .A2(KEYINPUT77), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n362), .B2(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n256), .B1(G1), .B2(new_n264), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT25), .B1(new_n253), .B2(new_n220), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n463), .A2(new_n220), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n437), .A2(new_n439), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT23), .B1(new_n467), .B2(new_n206), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n206), .A2(G87), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n285), .B2(new_n470), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT24), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n304), .A2(KEYINPUT22), .A3(G87), .A4(new_n284), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT83), .B(G116), .Z(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G33), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n473), .B(new_n474), .C1(new_n478), .C2(G20), .ZN(new_n479));
  AOI21_X1  g0279(.A(G20), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT24), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n466), .B1(new_n483), .B2(new_n255), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT80), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT80), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n489));
  AOI21_X1  g0289(.A(G41), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G41), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n205), .B(G45), .C1(new_n491), .C2(KEYINPUT5), .ZN(new_n492));
  OAI211_X1 g0292(.A(G264), .B(new_n313), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G250), .A2(G1698), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n227), .B2(G1698), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n304), .A3(new_n284), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n313), .B1(new_n499), .B2(KEYINPUT84), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n494), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n487), .A2(new_n489), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n491), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT79), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n492), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n486), .A2(G41), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(KEYINPUT79), .A3(new_n205), .A4(G45), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n505), .A2(new_n507), .A3(new_n322), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n422), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n510), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n376), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n485), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n500), .A2(new_n502), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n428), .A2(new_n515), .A3(new_n510), .A4(new_n493), .ZN(new_n516));
  AOI21_X1  g0316(.A(G200), .B1(new_n503), .B2(new_n510), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n484), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n514), .A2(new_n521), .A3(new_n518), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(new_n313), .C1(new_n490), .C2(new_n492), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT81), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n219), .A2(G1698), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n315), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT78), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n219), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(new_n364), .A3(new_n284), .A4(new_n271), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n284), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n369), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n510), .A2(new_n524), .A3(KEYINPUT81), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n527), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT82), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n527), .A2(new_n537), .A3(new_n541), .A4(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(G200), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(G33), .B1(new_n302), .B2(new_n303), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT7), .B(new_n206), .C1(new_n544), .C2(new_n272), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n440), .B1(new_n545), .B2(new_n269), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n547), .A2(new_n226), .A3(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n550), .A2(new_n206), .B1(new_n218), .B2(new_n265), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n255), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n378), .A2(G97), .ZN(new_n553));
  INV_X1    g0353(.A(new_n463), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n536), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n304), .A2(new_n284), .ZN(new_n558));
  INV_X1    g0358(.A(new_n528), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n532), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n313), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(new_n525), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n556), .B1(G190), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n543), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n525), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n537), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n376), .A2(new_n566), .B1(new_n552), .B2(new_n555), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n527), .A2(new_n537), .A3(new_n422), .A4(new_n538), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G87), .A2(G97), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n437), .A2(new_n439), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n413), .A2(new_n206), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n383), .A2(KEYINPUT19), .A3(new_n226), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n206), .A2(G68), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n558), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n255), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n463), .A2(new_n431), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n431), .A2(new_n253), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(G238), .A2(G1698), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n219), .B2(G1698), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(new_n304), .A3(new_n284), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n313), .B1(new_n585), .B2(new_n477), .ZN(new_n586));
  INV_X1    g0386(.A(G250), .ZN(new_n587));
  INV_X1    g0387(.A(G45), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G1), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n205), .A2(new_n320), .A3(G45), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n313), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n586), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n422), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n582), .B(new_n594), .C1(G169), .C2(new_n593), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n578), .A2(new_n255), .B1(new_n253), .B2(new_n431), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n315), .A2(new_n584), .B1(G33), .B2(new_n476), .ZN(new_n597));
  OAI211_X1 g0397(.A(G190), .B(new_n591), .C1(new_n597), .C2(new_n313), .ZN(new_n598));
  OAI21_X1  g0398(.A(G200), .B1(new_n586), .B2(new_n592), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n554), .A2(G87), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(G257), .A2(G1698), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n221), .B2(G1698), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n315), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n285), .A2(G303), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n313), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n313), .B1(new_n490), .B2(new_n492), .ZN(new_n608));
  INV_X1    g0408(.A(G270), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n510), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G190), .ZN(new_n612));
  INV_X1    g0412(.A(G116), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n463), .A2(new_n613), .B1(new_n378), .B2(new_n476), .ZN(new_n614));
  XNOR2_X1  g0414(.A(KEYINPUT83), .B(G116), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n295), .B1(G20), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G20), .B1(new_n264), .B2(G97), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n531), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n618), .A3(KEYINPUT20), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G200), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n612), .B(new_n623), .C1(new_n624), .C2(new_n611), .ZN(new_n625));
  OAI21_X1  g0425(.A(G169), .B1(new_n607), .B2(new_n610), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n622), .ZN(new_n628));
  INV_X1    g0428(.A(new_n614), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n630), .A3(KEYINPUT21), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n623), .B2(new_n626), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(G179), .A3(new_n611), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n625), .A2(new_n631), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n570), .A2(new_n602), .A3(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n462), .A2(new_n523), .A3(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n591), .A2(KEYINPUT86), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT86), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n313), .A2(new_n589), .A3(new_n590), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(G200), .B1(new_n586), .B2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n596), .A2(new_n598), .A3(new_n600), .A4(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n376), .B1(new_n586), .B2(new_n641), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT87), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(KEYINPUT87), .B(new_n376), .C1(new_n586), .C2(new_n641), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n596), .A2(new_n580), .B1(new_n422), .B2(new_n593), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n643), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n564), .A2(new_n518), .A3(new_n650), .A4(new_n569), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n376), .B1(new_n561), .B2(new_n525), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n556), .A2(new_n568), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n543), .B2(new_n563), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n656), .A2(KEYINPUT88), .A3(new_n518), .A4(new_n650), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n514), .A2(new_n633), .A3(new_n634), .A4(new_n631), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n646), .A2(new_n582), .A3(new_n594), .A4(new_n647), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT89), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n648), .A2(new_n662), .A3(new_n649), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n596), .A2(new_n598), .A3(new_n600), .A4(new_n642), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n660), .A2(new_n567), .A3(new_n568), .A4(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n661), .B(new_n663), .C1(new_n665), .C2(KEYINPUT26), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n595), .A2(new_n601), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n655), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT90), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n650), .A2(new_n667), .A3(new_n655), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n663), .A2(new_n661), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT26), .B1(new_n602), .B2(new_n569), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT90), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n671), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n462), .B1(new_n659), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n329), .A2(new_n331), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT18), .B1(new_n358), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n311), .A2(new_n360), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n345), .A2(new_n359), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n452), .A2(new_n453), .A3(new_n436), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n429), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n425), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n682), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT91), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n688), .A2(KEYINPUT91), .B1(new_n397), .B2(new_n399), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n391), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n677), .A2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(G213), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n523), .B1(new_n484), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT92), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n485), .A2(new_n511), .A3(new_n513), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n698), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n631), .A2(new_n634), .A3(new_n633), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n623), .A2(new_n699), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n635), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n708), .A2(new_n699), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n701), .A2(new_n702), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n704), .A2(new_n699), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OR2_X1    g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n209), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G1), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n440), .A2(new_n613), .A3(new_n572), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n723), .B1(new_n212), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n636), .A2(new_n520), .A3(new_n522), .A4(new_n699), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n562), .A2(new_n611), .A3(G179), .A4(new_n593), .ZN(new_n728));
  INV_X1    g0528(.A(new_n503), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n586), .A2(new_n641), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n611), .A2(G179), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n512), .A3(new_n539), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n728), .A2(new_n727), .A3(new_n729), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n698), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n726), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n668), .A2(new_n667), .A3(new_n655), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n672), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n704), .A2(new_n708), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT93), .B1(new_n746), .B2(new_n651), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT93), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n518), .A2(new_n650), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n658), .A2(new_n748), .A3(new_n749), .A4(new_n656), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n745), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n698), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT29), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n699), .B1(new_n659), .B2(new_n676), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT29), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n742), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n725), .B1(new_n757), .B2(G1), .ZN(G364));
  NOR2_X1   g0558(.A1(new_n252), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n205), .B1(new_n759), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n720), .A2(new_n761), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n206), .A2(new_n428), .A3(new_n624), .A4(G179), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G87), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n206), .A2(G190), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(new_n422), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n285), .B(new_n766), .C1(G107), .C2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT95), .Z(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n263), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT32), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n767), .A2(G179), .A3(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n206), .A2(new_n422), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n428), .A3(new_n624), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n776), .B1(new_n296), .B2(new_n777), .C1(new_n218), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n624), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n224), .B1(new_n785), .B2(new_n380), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n206), .B1(new_n772), .B2(G190), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n774), .A2(new_n775), .B1(new_n226), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n780), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n268), .B1(new_n763), .B2(G303), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  INV_X1    g0592(.A(G326), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n783), .A2(new_n792), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n777), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  INV_X1    g0596(.A(new_n773), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n799), .B2(new_n768), .C1(new_n800), .C2(new_n779), .ZN(new_n801));
  INV_X1    g0601(.A(new_n787), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n794), .B(new_n801), .C1(G294), .C2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n771), .A2(new_n789), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n214), .B1(G20), .B2(new_n376), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n762), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n805), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n242), .A2(G45), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n719), .A2(new_n315), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n588), .B2(new_n213), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n719), .A2(new_n285), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G355), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n209), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n812), .A2(new_n815), .B1(new_n818), .B2(KEYINPUT94), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(KEYINPUT94), .B2(new_n818), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n807), .B1(new_n811), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n810), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n711), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n762), .B1(new_n711), .B2(G330), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(G330), .B2(new_n711), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n685), .A2(new_n699), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n447), .A2(new_n450), .B1(new_n436), .B2(new_n698), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n685), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n754), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n829), .A2(new_n685), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n454), .A2(new_n698), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n699), .B(new_n834), .C1(new_n659), .C2(new_n676), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n762), .B1(new_n836), .B2(new_n741), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n742), .A2(new_n831), .A3(new_n835), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n805), .A2(new_n808), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n762), .B1(G77), .B2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT97), .Z(new_n843));
  OAI22_X1  g0643(.A1(new_n768), .A2(new_n765), .B1(new_n773), .B2(new_n800), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n285), .B1(new_n764), .B2(new_n220), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(G303), .C2(new_n784), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n782), .A2(G294), .B1(G97), .B2(new_n802), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n779), .A2(new_n615), .B1(new_n777), .B2(new_n799), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT98), .Z(new_n850));
  AND3_X1   g0650(.A1(new_n846), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n779), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G159), .A2(new_n852), .B1(new_n795), .B2(G150), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G143), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n785), .C1(new_n855), .C2(new_n783), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT34), .ZN(new_n857));
  INV_X1    g0657(.A(G132), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n764), .A2(new_n380), .B1(new_n773), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n315), .B1(new_n224), .B2(new_n787), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n768), .A2(new_n296), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n851), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n843), .B1(new_n806), .B2(new_n863), .C1(new_n834), .C2(new_n809), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT100), .Z(new_n865));
  NOR2_X1   g0665(.A1(new_n839), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  INV_X1    g0667(.A(new_n550), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n868), .A2(KEYINPUT35), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(KEYINPUT35), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n869), .A2(G116), .A3(new_n215), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT36), .Z(new_n872));
  OR4_X1    g0672(.A1(new_n218), .A2(new_n259), .A3(new_n260), .A4(new_n212), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n380), .A2(G68), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n205), .B(G13), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n308), .B1(new_n307), .B2(new_n278), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n696), .B1(new_n877), .B2(new_n257), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n362), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n343), .B1(new_n358), .B2(new_n696), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n332), .A2(new_n333), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n881), .B1(new_n358), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n877), .A2(new_n257), .B1(new_n678), .B2(new_n696), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n358), .B2(new_n342), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n880), .A2(new_n883), .B1(new_n885), .B2(new_n881), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT104), .ZN(new_n888));
  INV_X1    g0688(.A(new_n696), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n311), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n335), .A2(new_n890), .A3(new_n881), .A4(new_n343), .ZN(new_n891));
  INV_X1    g0691(.A(new_n343), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n892), .B2(new_n884), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n888), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n879), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT38), .B(new_n879), .C1(new_n887), .C2(new_n894), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n358), .A2(new_n678), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n880), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n891), .ZN(new_n902));
  INV_X1    g0702(.A(new_n890), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n682), .B2(new_n683), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n896), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n425), .A2(new_n698), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n833), .B(KEYINPUT101), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n835), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT102), .B1(new_n835), .B2(new_n914), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n423), .A2(new_n424), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n410), .A2(new_n698), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n425), .A2(new_n429), .A3(new_n919), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(KEYINPUT103), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n425), .A2(new_n923), .A3(new_n429), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n898), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n891), .A2(new_n893), .A3(new_n888), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n929), .B2(new_n879), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n917), .B(new_n925), .C1(new_n926), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n682), .A2(new_n696), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n912), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n462), .A2(new_n753), .A3(new_n756), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n691), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT105), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n933), .B(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT106), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n902), .B2(new_n904), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n927), .A2(new_n928), .B1(new_n362), .B2(new_n878), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n939), .B1(new_n940), .B2(KEYINPUT38), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n830), .B1(new_n922), .B2(new_n924), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n740), .A3(KEYINPUT40), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n938), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n907), .A2(KEYINPUT106), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n740), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n897), .B2(new_n898), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(KEYINPUT40), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n462), .A2(new_n740), .ZN(new_n951));
  OAI21_X1  g0751(.A(G330), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n937), .A2(new_n953), .B1(new_n205), .B2(new_n759), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n937), .A2(new_n953), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n876), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT107), .ZN(G367));
  NAND2_X1  g0757(.A1(new_n596), .A2(new_n600), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n698), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n650), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n672), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n704), .A2(new_n564), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n698), .B1(new_n963), .B2(new_n569), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n556), .A2(new_n698), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n656), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n655), .A2(new_n698), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n715), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n964), .B1(new_n972), .B2(KEYINPUT42), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT42), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT109), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n972), .A2(new_n976), .A3(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n973), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n713), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n969), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n981), .B1(new_n978), .B2(new_n982), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n962), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n985), .ZN(new_n987));
  INV_X1    g0787(.A(new_n962), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n988), .A3(new_n983), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n720), .B(KEYINPUT41), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n717), .A2(new_n969), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT44), .Z(new_n993));
  NOR2_X1   g0793(.A1(new_n717), .A2(new_n969), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT45), .ZN(new_n995));
  AND3_X1   g0795(.A1(new_n993), .A2(new_n979), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n979), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n715), .B1(new_n706), .B2(new_n714), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(new_n712), .Z(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n757), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n996), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n991), .B1(new_n1001), .B2(new_n757), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n760), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n990), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g0805(.A1(new_n763), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G97), .B2(new_n769), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n795), .A2(G294), .B1(new_n797), .B2(G317), .ZN(new_n1008));
  AOI21_X1  g0808(.A(KEYINPUT46), .B1(new_n763), .B2(new_n476), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(G311), .B2(new_n784), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n315), .B1(G303), .B2(new_n782), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n852), .A2(G283), .B1(new_n802), .B2(new_n467), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT111), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n779), .A2(new_n380), .B1(new_n777), .B2(new_n263), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT112), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n285), .B1(new_n763), .B2(G58), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n769), .A2(G77), .B1(new_n797), .B2(G137), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n787), .A2(new_n296), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n782), .B2(G150), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n855), .B2(new_n785), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1012), .A2(new_n1014), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT47), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n806), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n811), .B1(new_n209), .B2(new_n431), .C1(new_n814), .C2(new_n238), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n762), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT110), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n961), .B2(new_n822), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1005), .A2(new_n1032), .ZN(G387));
  INV_X1    g0833(.A(new_n1000), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n721), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n757), .B2(new_n999), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n999), .A2(new_n761), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n783), .A2(new_n380), .B1(new_n785), .B2(new_n263), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n787), .A2(new_n431), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n764), .A2(new_n218), .B1(new_n773), .B2(new_n384), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G68), .B2(new_n852), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n250), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n795), .A2(new_n1043), .B1(new_n769), .B2(G97), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n315), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(G294), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n764), .A2(new_n1046), .B1(new_n787), .B2(new_n799), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G303), .A2(new_n852), .B1(new_n795), .B2(G311), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n782), .A2(G317), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n792), .C2(new_n785), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n768), .A2(new_n615), .B1(new_n773), .B2(new_n793), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n315), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1045), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n805), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n762), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n235), .A2(new_n588), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1062), .A2(new_n813), .B1(new_n723), .B2(new_n816), .ZN(new_n1063));
  AOI211_X1 g0863(.A(G45), .B(new_n723), .C1(G68), .C2(G77), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1043), .A2(new_n380), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT113), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT50), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1063), .A2(new_n1069), .B1(G107), .B2(new_n209), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1061), .B1(new_n1070), .B2(new_n811), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1060), .B(new_n1071), .C1(new_n706), .C2(new_n822), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1036), .A2(new_n1037), .A3(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n1001), .A2(new_n720), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT114), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n996), .B2(new_n997), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n997), .A2(new_n1075), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1034), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1074), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n761), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n811), .B1(new_n226), .B2(new_n209), .C1(new_n814), .C2(new_n245), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1081), .A2(new_n762), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n285), .B1(new_n787), .B2(new_n615), .C1(new_n220), .C2(new_n768), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(G294), .A2(new_n852), .B1(new_n795), .B2(G303), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n799), .B2(new_n764), .C1(new_n792), .C2(new_n773), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G311), .A2(new_n782), .B1(new_n784), .B2(G317), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1083), .B(new_n1085), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n852), .A2(new_n1043), .B1(new_n797), .B2(G143), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n380), .B2(new_n777), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n764), .A2(new_n296), .B1(new_n765), .B2(new_n768), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n787), .A2(new_n218), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1091), .A2(new_n558), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G150), .A2(new_n784), .B1(new_n782), .B2(G159), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1088), .A2(new_n1089), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1082), .B1(new_n806), .B2(new_n1098), .C1(new_n968), .C2(new_n822), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1080), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1079), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n742), .A2(new_n834), .A3(new_n925), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(KEYINPUT117), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n925), .B1(new_n915), .B2(new_n916), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n909), .A2(new_n899), .B1(new_n1108), .B2(new_n911), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n907), .A2(new_n911), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n913), .B1(new_n752), .B2(new_n834), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n925), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1106), .B(new_n1107), .C1(new_n1109), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1108), .A2(new_n911), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n910), .A2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1117), .A2(new_n1105), .A3(new_n1104), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1112), .B1(new_n741), .B2(new_n830), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1103), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n917), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1103), .A2(new_n1111), .A3(new_n1121), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n462), .A2(new_n742), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n934), .A2(new_n691), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n934), .A2(new_n691), .A3(new_n1126), .A4(KEYINPUT118), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n721), .B1(new_n1120), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1115), .A2(new_n1119), .A3(new_n1131), .A4(KEYINPUT119), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1115), .A2(new_n1119), .A3(new_n1131), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT120), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1133), .A2(new_n1137), .A3(KEYINPUT120), .A4(new_n1134), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n779), .A2(new_n1143), .B1(new_n773), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n763), .A2(G150), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(G137), .C2(new_n795), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n268), .B1(new_n768), .B2(new_n380), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n783), .A2(new_n858), .B1(new_n787), .B2(new_n263), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G128), .C2(new_n784), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n779), .A2(new_n226), .B1(new_n773), .B2(new_n1046), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n861), .B(new_n1153), .C1(new_n467), .C2(new_n795), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n783), .A2(new_n613), .B1(new_n785), .B2(new_n799), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1155), .A2(new_n766), .A3(new_n268), .A4(new_n1093), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1149), .A2(new_n1152), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n762), .B1(new_n1043), .B2(new_n841), .C1(new_n1157), .C2(new_n806), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n910), .B2(new_n808), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1120), .B2(new_n761), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1142), .A2(new_n1160), .ZN(G378));
  NAND2_X1  g0961(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1120), .B2(new_n1132), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT57), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT106), .B1(new_n907), .B2(new_n945), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n938), .B(new_n943), .C1(new_n898), .C2(new_n906), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(G330), .B1(new_n949), .B2(KEYINPUT40), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT122), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G330), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n948), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n926), .B2(new_n930), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT40), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT122), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n947), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n389), .A2(new_n889), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n400), .B(new_n1178), .Z(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1170), .A2(new_n1177), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1175), .A2(new_n947), .A3(new_n1181), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1184), .A2(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1175), .A2(new_n947), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1181), .B1(new_n1187), .B2(KEYINPUT122), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT123), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n1177), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1186), .A2(new_n933), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n933), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1165), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n933), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1184), .A2(KEYINPUT123), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1188), .B2(new_n1177), .ZN(new_n1196));
  AND4_X1   g0996(.A1(new_n1189), .A2(new_n1170), .A3(new_n1177), .A4(new_n1182), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1186), .A2(new_n933), .A3(new_n1190), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1163), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1193), .B(new_n720), .C1(new_n1200), .C2(KEYINPUT57), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1182), .A2(new_n808), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n762), .B1(G50), .B2(new_n841), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n782), .A2(G128), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n785), .B2(new_n1144), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1143), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n795), .A2(G132), .B1(new_n763), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n854), .B2(new_n779), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(G150), .C2(new_n802), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n769), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n768), .A2(new_n224), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G97), .B2(new_n795), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n315), .A2(G41), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n799), .C2(new_n773), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n783), .A2(new_n220), .B1(new_n785), .B2(new_n613), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n764), .A2(new_n218), .B1(new_n431), .B2(new_n779), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1021), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1219), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n380), .C1(G33), .C2(G41), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1223), .A2(KEYINPUT58), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1216), .A2(new_n1224), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1204), .B1(new_n1228), .B2(new_n805), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1202), .A2(new_n761), .B1(new_n1203), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1201), .A2(new_n1230), .ZN(G375));
  NAND3_X1  g1031(.A1(new_n1162), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n991), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1131), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1112), .A2(new_n808), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n783), .A2(new_n854), .B1(new_n787), .B2(new_n380), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G132), .B2(new_n784), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n852), .A2(G150), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n795), .A2(new_n1207), .B1(new_n797), .B2(G128), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n558), .B(new_n1217), .C1(G159), .C2(new_n763), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n268), .B(new_n1039), .C1(G77), .C2(new_n769), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n467), .A2(new_n852), .B1(new_n795), .B2(new_n476), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G303), .A2(new_n797), .B1(new_n763), .B2(G97), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G283), .A2(new_n782), .B1(new_n784), .B2(G294), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n806), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1061), .B(new_n1247), .C1(new_n296), .C2(new_n840), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1125), .A2(new_n761), .B1(new_n1235), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1234), .A2(new_n1249), .ZN(G381));
  NAND3_X1  g1050(.A1(new_n1005), .A2(new_n1032), .A3(new_n1101), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1138), .A2(new_n1160), .ZN(new_n1252));
  OR4_X1    g1052(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1253));
  OR4_X1    g1053(.A1(G375), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(G407));
  INV_X1    g1054(.A(new_n1252), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n697), .A2(G213), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G407), .B(G213), .C1(G375), .C2(new_n1258), .ZN(G409));
  AOI22_X1  g1059(.A1(new_n986), .A2(new_n989), .B1(new_n1003), .B2(new_n760), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1032), .ZN(new_n1261));
  OAI21_X1  g1061(.A(G390), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(new_n826), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1251), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1251), .B2(new_n1262), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n1232), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n720), .B1(new_n1270), .B2(new_n1232), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1249), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(new_n866), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n866), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(G2897), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1276), .B(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1200), .A2(new_n1233), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1252), .B1(new_n1230), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1201), .A2(G378), .A3(new_n1230), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1201), .A2(G378), .A3(KEYINPUT125), .A4(new_n1230), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1280), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1278), .B1(new_n1285), .B2(new_n1257), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1285), .A2(new_n1257), .A3(new_n1276), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1269), .B(new_n1286), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1280), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1257), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1276), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1268), .B1(new_n1289), .B2(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1286), .A2(new_n1269), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1295), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1298), .A2(new_n1267), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1302), .ZN(G405));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1251), .A2(new_n1262), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1263), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1251), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(KEYINPUT127), .A3(new_n1308), .ZN(new_n1309));
  XOR2_X1   g1109(.A(new_n1276), .B(KEYINPUT126), .Z(new_n1310));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1255), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1290), .B2(new_n1311), .ZN(new_n1312));
  OR2_X1    g1112(.A1(new_n1276), .A2(KEYINPUT126), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1290), .A2(new_n1311), .A3(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1305), .B(new_n1309), .C1(new_n1312), .C2(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1312), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1267), .A2(KEYINPUT127), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(G402));
endmodule


