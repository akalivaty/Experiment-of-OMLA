

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742;

  NOR2_X2 U371 ( .A1(n619), .A2(n714), .ZN(n622) );
  NOR2_X2 U372 ( .A1(n695), .A2(n714), .ZN(n697) );
  XNOR2_X1 U373 ( .A(n370), .B(n369), .ZN(n609) );
  NOR2_X1 U374 ( .A1(n373), .A2(n359), .ZN(n372) );
  NOR2_X1 U375 ( .A1(n742), .A2(n739), .ZN(n580) );
  NOR2_X1 U376 ( .A1(n664), .A2(n513), .ZN(n629) );
  NAND2_X1 U377 ( .A1(n396), .A2(n656), .ZN(n524) );
  NAND2_X1 U378 ( .A1(n522), .A2(n523), .ZN(n579) );
  NOR2_X2 U379 ( .A1(G902), .A2(n698), .ZN(n452) );
  INV_X1 U380 ( .A(KEYINPUT48), .ZN(n369) );
  INV_X4 U381 ( .A(G953), .ZN(n729) );
  AND2_X2 U382 ( .A1(n614), .A2(n649), .ZN(n710) );
  AND2_X1 U383 ( .A1(n647), .A2(n603), .ZN(n602) );
  NAND2_X1 U384 ( .A1(n372), .A2(n371), .ZN(n370) );
  XNOR2_X1 U385 ( .A(n580), .B(KEYINPUT46), .ZN(n371) );
  NOR2_X1 U386 ( .A1(n415), .A2(n629), .ZN(n519) );
  XNOR2_X1 U387 ( .A(n506), .B(KEYINPUT35), .ZN(n415) );
  NOR2_X1 U388 ( .A1(n712), .A2(G902), .ZN(n472) );
  XNOR2_X1 U389 ( .A(n365), .B(n364), .ZN(n712) );
  XNOR2_X1 U390 ( .A(n368), .B(n483), .ZN(n365) );
  XNOR2_X1 U391 ( .A(n366), .B(n466), .ZN(n364) );
  XNOR2_X1 U392 ( .A(n727), .B(n400), .ZN(n483) );
  XNOR2_X1 U393 ( .A(n402), .B(n401), .ZN(n727) );
  XNOR2_X1 U394 ( .A(n403), .B(KEYINPUT10), .ZN(n402) );
  XNOR2_X1 U395 ( .A(n363), .B(G110), .ZN(n446) );
  XNOR2_X1 U396 ( .A(n388), .B(G146), .ZN(n444) );
  NOR2_X2 U397 ( .A1(n553), .A2(n515), .ZN(n520) );
  OR2_X1 U398 ( .A1(G237), .A2(G902), .ZN(n433) );
  XNOR2_X1 U399 ( .A(n445), .B(n479), .ZN(n424) );
  XNOR2_X1 U400 ( .A(n444), .B(n387), .ZN(n445) );
  INV_X1 U401 ( .A(G137), .ZN(n387) );
  AND2_X1 U402 ( .A1(n417), .A2(n592), .ZN(n528) );
  INV_X1 U403 ( .A(n524), .ZN(n417) );
  XNOR2_X1 U404 ( .A(n664), .B(n418), .ZN(n553) );
  INV_X1 U405 ( .A(KEYINPUT6), .ZN(n418) );
  XNOR2_X1 U406 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U407 ( .A(n592), .ZN(n658) );
  NOR2_X1 U408 ( .A1(n409), .A2(n641), .ZN(n532) );
  XNOR2_X1 U409 ( .A(n591), .B(n360), .ZN(n359) );
  NOR2_X1 U410 ( .A1(n568), .A2(n567), .ZN(n581) );
  XNOR2_X1 U411 ( .A(n475), .B(KEYINPUT72), .ZN(n422) );
  XNOR2_X1 U412 ( .A(G125), .B(KEYINPUT68), .ZN(n401) );
  INV_X1 U413 ( .A(G140), .ZN(n403) );
  XNOR2_X1 U414 ( .A(n392), .B(KEYINPUT75), .ZN(n443) );
  XNOR2_X1 U415 ( .A(G143), .B(G128), .ZN(n392) );
  INV_X1 U416 ( .A(KEYINPUT4), .ZN(n388) );
  AND2_X1 U417 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U418 ( .A1(n578), .A2(n356), .ZN(n385) );
  NAND2_X1 U419 ( .A1(n586), .A2(n356), .ZN(n386) );
  NAND2_X1 U420 ( .A1(n383), .A2(n350), .ZN(n382) );
  OR2_X1 U421 ( .A1(n691), .A2(n603), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n428), .B(n427), .ZN(n473) );
  INV_X1 U423 ( .A(G119), .ZN(n427) );
  INV_X1 U424 ( .A(G107), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n460), .B(n459), .ZN(n500) );
  XOR2_X1 U426 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n459) );
  XNOR2_X1 U427 ( .A(n458), .B(n457), .ZN(n460) );
  INV_X1 U428 ( .A(KEYINPUT78), .ZN(n457) );
  XNOR2_X1 U429 ( .A(n498), .B(n351), .ZN(n391) );
  XOR2_X1 U430 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n498) );
  XNOR2_X1 U431 ( .A(n497), .B(n496), .ZN(n390) );
  INV_X1 U432 ( .A(KEYINPUT9), .ZN(n496) );
  XNOR2_X1 U433 ( .A(G116), .B(KEYINPUT7), .ZN(n497) );
  XNOR2_X1 U434 ( .A(n443), .B(n423), .ZN(n499) );
  INV_X1 U435 ( .A(G134), .ZN(n423) );
  NOR2_X1 U436 ( .A1(n539), .A2(n538), .ZN(n541) );
  AND2_X1 U437 ( .A1(n637), .A2(n551), .ZN(n552) );
  XNOR2_X1 U438 ( .A(n503), .B(n393), .ZN(n523) );
  XNOR2_X1 U439 ( .A(n504), .B(n394), .ZN(n393) );
  NOR2_X1 U440 ( .A1(G902), .A2(n708), .ZN(n503) );
  INV_X1 U441 ( .A(G472), .ZN(n419) );
  INV_X1 U442 ( .A(KEYINPUT101), .ZN(n395) );
  INV_X1 U443 ( .A(KEYINPUT1), .ZN(n416) );
  XNOR2_X1 U444 ( .A(n408), .B(n705), .ZN(n407) );
  XNOR2_X1 U445 ( .A(n704), .B(n357), .ZN(n705) );
  INV_X1 U446 ( .A(KEYINPUT76), .ZN(n360) );
  XOR2_X1 U447 ( .A(KEYINPUT69), .B(G131), .Z(n479) );
  NAND2_X1 U448 ( .A1(G953), .A2(G902), .ZN(n542) );
  INV_X1 U449 ( .A(G143), .ZN(n480) );
  INV_X1 U450 ( .A(n579), .ZN(n381) );
  INV_X1 U451 ( .A(G478), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n726), .B(n420), .ZN(n615) );
  XOR2_X1 U453 ( .A(G122), .B(G104), .Z(n486) );
  XNOR2_X1 U454 ( .A(G119), .B(G128), .ZN(n464) );
  XNOR2_X1 U455 ( .A(n463), .B(n367), .ZN(n366) );
  INV_X1 U456 ( .A(KEYINPUT24), .ZN(n367) );
  XNOR2_X1 U457 ( .A(G137), .B(G110), .ZN(n461) );
  INV_X1 U458 ( .A(G146), .ZN(n400) );
  XOR2_X1 U459 ( .A(G101), .B(G104), .Z(n449) );
  XNOR2_X1 U460 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n444), .B(n352), .ZN(n411) );
  XNOR2_X1 U462 ( .A(n443), .B(n432), .ZN(n412) );
  XNOR2_X1 U463 ( .A(n611), .B(n610), .ZN(n613) );
  INV_X1 U464 ( .A(KEYINPUT80), .ZN(n610) );
  NAND2_X1 U465 ( .A1(n384), .A2(n382), .ZN(n598) );
  OR2_X1 U466 ( .A1(n381), .A2(KEYINPUT40), .ZN(n380) );
  AND2_X1 U467 ( .A1(n381), .A2(KEYINPUT40), .ZN(n377) );
  XNOR2_X1 U468 ( .A(n477), .B(n355), .ZN(n684) );
  AND2_X1 U469 ( .A1(n553), .A2(n528), .ZN(n477) );
  NAND2_X1 U470 ( .A1(n577), .A2(n397), .ZN(n586) );
  XNOR2_X1 U471 ( .A(n398), .B(KEYINPUT73), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n435), .B(n434), .ZN(n564) );
  XNOR2_X1 U473 ( .A(n495), .B(n494), .ZN(n522) );
  XNOR2_X1 U474 ( .A(KEYINPUT13), .B(G475), .ZN(n494) );
  XNOR2_X1 U475 ( .A(n413), .B(n473), .ZN(n715) );
  XNOR2_X1 U476 ( .A(n429), .B(n486), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n446), .B(n362), .ZN(n429) );
  INV_X1 U478 ( .A(KEYINPUT16), .ZN(n362) );
  XNOR2_X1 U479 ( .A(n499), .B(n389), .ZN(n502) );
  XNOR2_X1 U480 ( .A(n391), .B(n390), .ZN(n389) );
  NAND2_X1 U481 ( .A1(n379), .A2(n376), .ZN(n739) );
  NAND2_X1 U482 ( .A1(n375), .A2(n374), .ZN(n379) );
  NAND2_X1 U483 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U484 ( .A1(n380), .A2(KEYINPUT40), .ZN(n374) );
  NOR2_X1 U485 ( .A1(n596), .A2(n593), .ZN(n554) );
  XNOR2_X1 U486 ( .A(n518), .B(n517), .ZN(n737) );
  NOR2_X1 U487 ( .A1(n564), .A2(n573), .ZN(n635) );
  XNOR2_X1 U488 ( .A(n527), .B(KEYINPUT93), .ZN(n409) );
  XNOR2_X1 U489 ( .A(n414), .B(KEYINPUT91), .ZN(n526) );
  INV_X1 U490 ( .A(KEYINPUT60), .ZN(n404) );
  NAND2_X1 U491 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U492 ( .A(n714), .ZN(n406) );
  NOR2_X1 U493 ( .A1(n578), .A2(n356), .ZN(n350) );
  NOR2_X1 U494 ( .A1(n556), .A2(n524), .ZN(n525) );
  XOR2_X1 U495 ( .A(G122), .B(G107), .Z(n351) );
  AND2_X1 U496 ( .A1(G224), .A2(n729), .ZN(n352) );
  AND2_X1 U497 ( .A1(G210), .A2(n433), .ZN(n353) );
  AND2_X1 U498 ( .A1(n382), .A2(n380), .ZN(n354) );
  XOR2_X1 U499 ( .A(KEYINPUT83), .B(KEYINPUT33), .Z(n355) );
  XOR2_X1 U500 ( .A(KEYINPUT39), .B(KEYINPUT70), .Z(n356) );
  XNOR2_X1 U501 ( .A(n424), .B(n499), .ZN(n726) );
  XNOR2_X1 U502 ( .A(n715), .B(n410), .ZN(n691) );
  XNOR2_X1 U503 ( .A(n726), .B(n451), .ZN(n698) );
  XNOR2_X1 U504 ( .A(G902), .B(KEYINPUT15), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n357) );
  NAND2_X1 U506 ( .A1(n358), .A2(n584), .ZN(n590) );
  NAND2_X1 U507 ( .A1(n583), .A2(KEYINPUT47), .ZN(n358) );
  INV_X1 U508 ( .A(n664), .ZN(n559) );
  BUF_X1 U509 ( .A(n612), .Z(n718) );
  XNOR2_X2 U510 ( .A(n361), .B(n353), .ZN(n569) );
  NAND2_X1 U511 ( .A1(n500), .A2(G221), .ZN(n368) );
  INV_X1 U512 ( .A(n581), .ZN(n373) );
  NAND2_X1 U513 ( .A1(n354), .A2(n384), .ZN(n375) );
  INV_X1 U514 ( .A(n598), .ZN(n378) );
  INV_X1 U515 ( .A(n586), .ZN(n383) );
  XNOR2_X2 U516 ( .A(n556), .B(n416), .ZN(n592) );
  XNOR2_X2 U517 ( .A(n452), .B(G469), .ZN(n556) );
  XNOR2_X2 U518 ( .A(n579), .B(KEYINPUT103), .ZN(n637) );
  NOR2_X1 U519 ( .A1(n396), .A2(n576), .ZN(n549) );
  XNOR2_X1 U520 ( .A(n396), .B(n395), .ZN(n655) );
  NOR2_X1 U521 ( .A1(n515), .A2(n396), .ZN(n512) );
  XNOR2_X2 U522 ( .A(n472), .B(n471), .ZN(n396) );
  NAND2_X1 U523 ( .A1(n525), .A2(n399), .ZN(n398) );
  INV_X1 U524 ( .A(n576), .ZN(n399) );
  XNOR2_X1 U525 ( .A(n405), .B(n404), .ZN(G60) );
  NAND2_X1 U526 ( .A1(n710), .A2(G475), .ZN(n408) );
  NOR2_X2 U527 ( .A1(n564), .A2(n440), .ZN(n441) );
  NAND2_X1 U528 ( .A1(n409), .A2(n640), .ZN(n625) );
  NAND2_X1 U529 ( .A1(n409), .A2(n637), .ZN(n624) );
  INV_X1 U530 ( .A(n530), .ZN(n507) );
  NAND2_X1 U531 ( .A1(n530), .A2(n525), .ZN(n414) );
  XNOR2_X2 U532 ( .A(n441), .B(n442), .ZN(n530) );
  XNOR2_X1 U533 ( .A(n415), .B(G122), .ZN(n736) );
  XNOR2_X2 U534 ( .A(n476), .B(n419), .ZN(n664) );
  XNOR2_X1 U535 ( .A(n473), .B(n421), .ZN(n420) );
  XNOR2_X1 U536 ( .A(n422), .B(n474), .ZN(n421) );
  AND2_X2 U537 ( .A1(n609), .A2(n607), .ZN(n647) );
  NOR2_X1 U538 ( .A1(n615), .A2(G902), .ZN(n476) );
  INV_X1 U539 ( .A(n669), .ZN(n550) );
  XNOR2_X1 U540 ( .A(n470), .B(KEYINPUT74), .ZN(n471) );
  XNOR2_X1 U541 ( .A(n541), .B(n540), .ZN(n612) );
  INV_X1 U542 ( .A(KEYINPUT100), .ZN(n504) );
  INV_X1 U543 ( .A(KEYINPUT19), .ZN(n434) );
  XNOR2_X1 U544 ( .A(n616), .B(KEYINPUT62), .ZN(n617) );
  XNOR2_X1 U545 ( .A(n691), .B(n692), .ZN(n693) );
  XNOR2_X1 U546 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U547 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U548 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n517) );
  XNOR2_X1 U549 ( .A(n620), .B(KEYINPUT63), .ZN(n621) );
  NOR2_X1 U550 ( .A1(G952), .A2(n729), .ZN(n714) );
  XNOR2_X1 U551 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n442) );
  NAND2_X1 U552 ( .A1(G214), .A2(n433), .ZN(n669) );
  INV_X1 U553 ( .A(n453), .ZN(n603) );
  XOR2_X1 U554 ( .A(KEYINPUT3), .B(G116), .Z(n426) );
  XNOR2_X1 U555 ( .A(G113), .B(G101), .ZN(n425) );
  XNOR2_X1 U556 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n431) );
  XNOR2_X1 U558 ( .A(G125), .B(KEYINPUT18), .ZN(n430) );
  XNOR2_X1 U559 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U560 ( .A1(n669), .A2(n569), .ZN(n435) );
  NAND2_X1 U561 ( .A1(G952), .A2(n729), .ZN(n546) );
  INV_X1 U562 ( .A(n546), .ZN(n437) );
  NOR2_X1 U563 ( .A1(G898), .A2(n542), .ZN(n436) );
  NOR2_X1 U564 ( .A1(n437), .A2(n436), .ZN(n439) );
  NAND2_X1 U565 ( .A1(G234), .A2(G237), .ZN(n438) );
  XNOR2_X1 U566 ( .A(KEYINPUT14), .B(n438), .ZN(n654) );
  INV_X1 U567 ( .A(n654), .ZN(n545) );
  OR2_X1 U568 ( .A1(n439), .A2(n545), .ZN(n440) );
  XOR2_X1 U569 ( .A(G140), .B(n446), .Z(n448) );
  NAND2_X1 U570 ( .A1(G227), .A2(n729), .ZN(n447) );
  XNOR2_X1 U571 ( .A(n448), .B(n447), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U573 ( .A1(G234), .A2(n453), .ZN(n454) );
  XNOR2_X1 U574 ( .A(KEYINPUT20), .B(n454), .ZN(n467) );
  NAND2_X1 U575 ( .A1(n467), .A2(G221), .ZN(n455) );
  XNOR2_X1 U576 ( .A(n455), .B(KEYINPUT21), .ZN(n456) );
  XOR2_X1 U577 ( .A(KEYINPUT90), .B(n456), .Z(n656) );
  NAND2_X1 U578 ( .A1(G234), .A2(n729), .ZN(n458) );
  XOR2_X1 U579 ( .A(KEYINPUT87), .B(KEYINPUT23), .Z(n462) );
  XNOR2_X1 U580 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U581 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n465) );
  XNOR2_X1 U582 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U583 ( .A(KEYINPUT25), .B(KEYINPUT89), .Z(n469) );
  NAND2_X1 U584 ( .A1(n467), .A2(G217), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U586 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n474) );
  NOR2_X1 U587 ( .A1(G953), .A2(G237), .ZN(n487) );
  AND2_X1 U588 ( .A1(n487), .A2(G210), .ZN(n475) );
  NOR2_X1 U589 ( .A1(n507), .A2(n684), .ZN(n478) );
  XNOR2_X1 U590 ( .A(n478), .B(KEYINPUT34), .ZN(n505) );
  XNOR2_X1 U591 ( .A(G113), .B(n479), .ZN(n481) );
  XNOR2_X1 U592 ( .A(n483), .B(n482), .ZN(n493) );
  XOR2_X1 U593 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n485) );
  XNOR2_X1 U594 ( .A(KEYINPUT95), .B(KEYINPUT97), .ZN(n484) );
  XNOR2_X1 U595 ( .A(n485), .B(n484), .ZN(n491) );
  XOR2_X1 U596 ( .A(KEYINPUT12), .B(n486), .Z(n489) );
  NAND2_X1 U597 ( .A1(G214), .A2(n487), .ZN(n488) );
  XNOR2_X1 U598 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U599 ( .A(n491), .B(n490), .Z(n492) );
  XNOR2_X1 U600 ( .A(n493), .B(n492), .ZN(n704) );
  NOR2_X1 U601 ( .A1(G902), .A2(n704), .ZN(n495) );
  INV_X1 U602 ( .A(n522), .ZN(n508) );
  NAND2_X1 U603 ( .A1(G217), .A2(n500), .ZN(n501) );
  XNOR2_X1 U604 ( .A(n502), .B(n501), .ZN(n708) );
  NOR2_X1 U605 ( .A1(n508), .A2(n523), .ZN(n585) );
  NAND2_X1 U606 ( .A1(n505), .A2(n585), .ZN(n506) );
  INV_X1 U607 ( .A(n656), .ZN(n509) );
  NAND2_X1 U608 ( .A1(n523), .A2(n508), .ZN(n672) );
  NOR2_X1 U609 ( .A1(n509), .A2(n672), .ZN(n510) );
  NAND2_X1 U610 ( .A1(n530), .A2(n510), .ZN(n511) );
  XNOR2_X1 U611 ( .A(KEYINPUT22), .B(n511), .ZN(n515) );
  NAND2_X1 U612 ( .A1(n658), .A2(n512), .ZN(n513) );
  NOR2_X1 U613 ( .A1(n658), .A2(n655), .ZN(n514) );
  XNOR2_X1 U614 ( .A(KEYINPUT102), .B(n514), .ZN(n516) );
  NAND2_X1 U615 ( .A1(n516), .A2(n520), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n519), .A2(n737), .ZN(n537) );
  NAND2_X1 U617 ( .A1(n537), .A2(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U618 ( .A1(n520), .A2(n655), .ZN(n521) );
  NOR2_X1 U619 ( .A1(n592), .A2(n521), .ZN(n623) );
  NOR2_X1 U620 ( .A1(n522), .A2(n523), .ZN(n640) );
  INV_X1 U621 ( .A(n640), .ZN(n599) );
  NAND2_X1 U622 ( .A1(n599), .A2(n579), .ZN(n565) );
  INV_X1 U623 ( .A(n565), .ZN(n675) );
  NAND2_X1 U624 ( .A1(n526), .A2(n559), .ZN(n527) );
  NAND2_X1 U625 ( .A1(n528), .A2(n664), .ZN(n529) );
  XOR2_X1 U626 ( .A(KEYINPUT94), .B(n529), .Z(n666) );
  NAND2_X1 U627 ( .A1(n666), .A2(n530), .ZN(n531) );
  XNOR2_X1 U628 ( .A(n531), .B(KEYINPUT31), .ZN(n641) );
  NOR2_X1 U629 ( .A1(n675), .A2(n532), .ZN(n533) );
  NOR2_X1 U630 ( .A1(n623), .A2(n533), .ZN(n534) );
  NAND2_X1 U631 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT82), .ZN(n539) );
  NOR2_X1 U633 ( .A1(n537), .A2(KEYINPUT44), .ZN(n538) );
  INV_X1 U634 ( .A(KEYINPUT45), .ZN(n540) );
  INV_X1 U635 ( .A(n569), .ZN(n596) );
  NOR2_X1 U636 ( .A1(n545), .A2(n542), .ZN(n543) );
  XOR2_X1 U637 ( .A(KEYINPUT104), .B(n543), .Z(n544) );
  NOR2_X1 U638 ( .A1(G900), .A2(n544), .ZN(n548) );
  NOR2_X1 U639 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U640 ( .A1(n548), .A2(n547), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n656), .A2(n549), .ZN(n558) );
  NOR2_X1 U642 ( .A1(n558), .A2(n550), .ZN(n551) );
  NAND2_X1 U643 ( .A1(n553), .A2(n552), .ZN(n593) );
  XNOR2_X1 U644 ( .A(n554), .B(KEYINPUT36), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n555), .A2(n592), .ZN(n645) );
  XNOR2_X1 U646 ( .A(n645), .B(KEYINPUT81), .ZN(n568) );
  INV_X1 U647 ( .A(n556), .ZN(n557) );
  XOR2_X1 U648 ( .A(KEYINPUT107), .B(n557), .Z(n563) );
  NOR2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U650 ( .A(KEYINPUT28), .B(KEYINPUT108), .ZN(n560) );
  XNOR2_X1 U651 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n573) );
  NAND2_X1 U653 ( .A1(n635), .A2(n565), .ZN(n566) );
  NOR2_X1 U654 ( .A1(n566), .A2(KEYINPUT47), .ZN(n567) );
  XNOR2_X1 U655 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n570) );
  XOR2_X1 U656 ( .A(n570), .B(n569), .Z(n578) );
  INV_X1 U657 ( .A(n578), .ZN(n670) );
  NAND2_X1 U658 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U659 ( .A1(n672), .A2(n674), .ZN(n572) );
  XOR2_X1 U660 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n571) );
  XNOR2_X1 U661 ( .A(n572), .B(n571), .ZN(n685) );
  NOR2_X1 U662 ( .A1(n685), .A2(n573), .ZN(n574) );
  XNOR2_X1 U663 ( .A(n574), .B(KEYINPUT42), .ZN(n742) );
  NAND2_X1 U664 ( .A1(n664), .A2(n669), .ZN(n575) );
  XOR2_X1 U665 ( .A(KEYINPUT30), .B(n575), .Z(n577) );
  NAND2_X1 U666 ( .A1(n675), .A2(KEYINPUT47), .ZN(n582) );
  XOR2_X1 U667 ( .A(n582), .B(KEYINPUT77), .Z(n584) );
  INV_X1 U668 ( .A(n635), .ZN(n583) );
  INV_X1 U669 ( .A(n585), .ZN(n589) );
  NOR2_X1 U670 ( .A1(n596), .A2(n586), .ZN(n587) );
  XOR2_X1 U671 ( .A(KEYINPUT106), .B(n587), .Z(n588) );
  NOR2_X1 U672 ( .A1(n589), .A2(n588), .ZN(n633) );
  NOR2_X1 U673 ( .A1(n590), .A2(n633), .ZN(n591) );
  XOR2_X1 U674 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n595) );
  OR2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U676 ( .A(n595), .B(n594), .ZN(n597) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(n646) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT110), .ZN(n741) );
  INV_X1 U680 ( .A(n741), .ZN(n601) );
  AND2_X1 U681 ( .A1(n646), .A2(n601), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n612), .A2(n602), .ZN(n606) );
  INV_X1 U683 ( .A(KEYINPUT2), .ZN(n604) );
  OR2_X1 U684 ( .A1(n453), .A2(n604), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n614) );
  AND2_X1 U686 ( .A1(n607), .A2(KEYINPUT2), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n649) );
  NAND2_X1 U689 ( .A1(n710), .A2(G472), .ZN(n618) );
  XOR2_X1 U690 ( .A(n615), .B(KEYINPUT111), .Z(n616) );
  XOR2_X1 U691 ( .A(KEYINPUT84), .B(KEYINPUT112), .Z(n620) );
  XNOR2_X1 U692 ( .A(n622), .B(n621), .ZN(G57) );
  XOR2_X1 U693 ( .A(G101), .B(n623), .Z(G3) );
  XNOR2_X1 U694 ( .A(n624), .B(G104), .ZN(G6) );
  XOR2_X1 U695 ( .A(G107), .B(KEYINPUT27), .Z(n626) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(n628) );
  XOR2_X1 U697 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(G9) );
  XOR2_X1 U699 ( .A(G110), .B(n629), .Z(G12) );
  XOR2_X1 U700 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n631) );
  NAND2_X1 U701 ( .A1(n635), .A2(n640), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(G128), .B(n632), .ZN(G30) );
  XNOR2_X1 U704 ( .A(G143), .B(n633), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT115), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n635), .A2(n637), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n637), .A2(n641), .ZN(n638) );
  XNOR2_X1 U709 ( .A(n638), .B(KEYINPUT116), .ZN(n639) );
  XNOR2_X1 U710 ( .A(G113), .B(n639), .ZN(G15) );
  XOR2_X1 U711 ( .A(G116), .B(KEYINPUT117), .Z(n643) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G18) );
  XOR2_X1 U714 ( .A(G125), .B(KEYINPUT37), .Z(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G140), .B(n646), .ZN(G42) );
  NOR2_X1 U717 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n648), .B(KEYINPUT79), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n652) );
  NOR2_X1 U720 ( .A1(n718), .A2(KEYINPUT2), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U722 ( .A1(G953), .A2(n653), .ZN(n689) );
  NAND2_X1 U723 ( .A1(G952), .A2(n654), .ZN(n683) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT49), .B(n657), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n524), .A2(n658), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n659), .B(KEYINPUT50), .ZN(n660) );
  XNOR2_X1 U728 ( .A(KEYINPUT118), .B(n660), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n667), .Z(n668) );
  NOR2_X1 U733 ( .A1(n685), .A2(n668), .ZN(n680) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U736 ( .A(KEYINPUT119), .B(n673), .Z(n677) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n684), .A2(n678), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U741 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  NOR2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n687) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U746 ( .A(KEYINPUT53), .B(n690), .Z(G75) );
  NAND2_X1 U747 ( .A1(n710), .A2(G210), .ZN(n694) );
  XOR2_X1 U748 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n692) );
  XNOR2_X1 U749 ( .A(KEYINPUT56), .B(KEYINPUT120), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(G51) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n700) );
  XNOR2_X1 U752 ( .A(n698), .B(KEYINPUT121), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n710), .A2(G469), .ZN(n701) );
  XOR2_X1 U755 ( .A(n702), .B(n701), .Z(n703) );
  NOR2_X1 U756 ( .A1(n714), .A2(n703), .ZN(G54) );
  NAND2_X1 U757 ( .A1(n710), .A2(G478), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n706), .B(KEYINPUT122), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U760 ( .A1(n714), .A2(n709), .ZN(G63) );
  NAND2_X1 U761 ( .A1(G217), .A2(n710), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U763 ( .A1(n714), .A2(n713), .ZN(G66) );
  OR2_X1 U764 ( .A1(G898), .A2(n729), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n717), .B(KEYINPUT124), .ZN(n725) );
  NAND2_X1 U767 ( .A1(n718), .A2(n729), .ZN(n723) );
  NAND2_X1 U768 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U770 ( .A1(n720), .A2(G898), .ZN(n721) );
  XOR2_X1 U771 ( .A(KEYINPUT123), .B(n721), .Z(n722) );
  NAND2_X1 U772 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U773 ( .A(n725), .B(n724), .Z(G69) );
  XOR2_X1 U774 ( .A(n726), .B(n727), .Z(n731) );
  INV_X1 U775 ( .A(n731), .ZN(n728) );
  XOR2_X1 U776 ( .A(n728), .B(n647), .Z(n730) );
  NAND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n735) );
  XOR2_X1 U778 ( .A(G227), .B(n731), .Z(n732) );
  NAND2_X1 U779 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U780 ( .A1(n733), .A2(G953), .ZN(n734) );
  NAND2_X1 U781 ( .A1(n735), .A2(n734), .ZN(G72) );
  XNOR2_X1 U782 ( .A(n736), .B(KEYINPUT125), .ZN(G24) );
  XNOR2_X1 U783 ( .A(G119), .B(KEYINPUT126), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n738), .B(n737), .ZN(G21) );
  XNOR2_X1 U785 ( .A(G131), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(G33) );
  XOR2_X1 U787 ( .A(G134), .B(n741), .Z(G36) );
  XOR2_X1 U788 ( .A(G137), .B(n742), .Z(G39) );
endmodule

