//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n205), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G107), .A2(G264), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n211), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n227), .A2(G20), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n214), .A2(new_n223), .A3(new_n224), .A4(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT66), .Z(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT76), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(G232), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT74), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT74), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G232), .A4(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1698), .B1(new_n257), .B2(new_n258), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n263), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n250), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(new_n250), .A3(G274), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n228), .B2(new_n249), .ZN(new_n273));
  AOI21_X1  g0073(.A(KEYINPUT68), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  INV_X1    g0074(.A(G238), .ZN(new_n275));
  INV_X1    g0075(.A(new_n268), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n250), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n271), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT13), .B1(new_n265), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n270), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n282));
  INV_X1    g0082(.A(new_n250), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n268), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n281), .A2(new_n282), .B1(new_n284), .B2(G238), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  OAI211_X1 g0086(.A(G226), .B(new_n286), .C1(new_n251), .C2(new_n252), .ZN(new_n287));
  INV_X1    g0087(.A(G97), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n256), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n261), .B2(new_n254), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n280), .B(new_n285), .C1(new_n290), .C2(new_n250), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n279), .A2(new_n291), .A3(G190), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G1), .A2(G13), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n209), .A2(G33), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n296), .A2(new_n205), .B1(new_n209), .B2(G68), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n297), .A2(new_n298), .B1(new_n202), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT11), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  OAI211_X1 g0110(.A(KEYINPUT11), .B(new_n295), .C1(new_n301), .C2(new_n302), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT73), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n307), .B2(new_n295), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n294), .A4(new_n293), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n208), .A2(G20), .ZN(new_n315));
  AND3_X1   g0115(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G68), .ZN(new_n317));
  AND4_X1   g0117(.A1(new_n305), .A2(new_n310), .A3(new_n311), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n292), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n279), .B2(new_n291), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n248), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n321), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n323), .A2(KEYINPUT76), .A3(new_n292), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n318), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n279), .A2(new_n291), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G169), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n279), .A2(new_n291), .A3(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n328), .B1(new_n327), .B2(G169), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n208), .B2(G20), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n307), .A2(new_n295), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(new_n307), .B2(new_n336), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n257), .A2(new_n209), .A3(new_n258), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n308), .B1(new_n340), .B2(KEYINPUT7), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n251), .A2(new_n252), .A3(G20), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G58), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n308), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n347), .B2(new_n201), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n299), .A2(G159), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(new_n351), .A3(KEYINPUT16), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n295), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n258), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n342), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n350), .B1(new_n356), .B2(G68), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT16), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n339), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G232), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n271), .A2(new_n274), .B1(new_n360), .B2(new_n277), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n286), .B1(new_n257), .B2(new_n258), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n263), .A2(G223), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n250), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(G226), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G87), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n283), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n281), .A2(new_n282), .B1(new_n284), .B2(G232), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n359), .A2(new_n373), .A3(KEYINPUT18), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT18), .B1(new_n359), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n339), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n350), .B1(new_n344), .B2(new_n341), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(KEYINPUT16), .B1(new_n294), .B2(new_n293), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n356), .A2(G68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n351), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT78), .B(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n370), .A2(new_n371), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G200), .B1(new_n361), .B2(new_n365), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n384), .A2(KEYINPUT17), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n352), .B(new_n295), .C1(KEYINPUT16), .C2(new_n357), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n389), .A2(new_n339), .A3(new_n387), .A4(new_n386), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n376), .A2(new_n393), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n271), .A2(new_n274), .B1(new_n215), .B2(new_n277), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n263), .A2(G232), .ZN(new_n397));
  INV_X1    g0197(.A(G107), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(new_n398), .B2(new_n259), .ZN(new_n399));
  XOR2_X1   g0199(.A(new_n362), .B(KEYINPUT69), .Z(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(G238), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n396), .B1(new_n401), .B2(new_n250), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n316), .A2(G77), .ZN(new_n406));
  INV_X1    g0206(.A(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT15), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n296), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n336), .A2(new_n300), .B1(new_n209), .B2(new_n205), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n295), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n406), .B(new_n415), .C1(G77), .C2(new_n306), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G169), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n402), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n405), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n403), .A2(new_n320), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n417), .B1(new_n402), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n394), .B(new_n420), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n271), .A2(new_n274), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(G226), .B2(new_n284), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n263), .A2(G222), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n205), .B2(new_n259), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n400), .B2(G223), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(new_n250), .ZN(new_n430));
  INV_X1    g0230(.A(G150), .ZN(new_n431));
  OAI22_X1  g0231(.A1(new_n336), .A2(new_n296), .B1(new_n431), .B2(new_n300), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n204), .A2(new_n209), .B1(new_n432), .B2(KEYINPUT70), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(KEYINPUT70), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n295), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n338), .A2(new_n436), .B1(new_n202), .B2(new_n307), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT9), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n430), .A2(G200), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n430), .A2(new_n422), .B1(new_n438), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT10), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n442), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT10), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n440), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n430), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n438), .B1(new_n448), .B2(G169), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT71), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT72), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n430), .B2(G179), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT71), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n438), .C1(new_n448), .C2(G169), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(KEYINPUT72), .A3(new_n404), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n450), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n335), .A2(new_n424), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n411), .A2(new_n306), .ZN(new_n460));
  NAND3_X1  g0260(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n209), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n407), .A2(new_n288), .A3(new_n398), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n209), .B(G68), .C1(new_n251), .C2(new_n252), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n296), .B2(new_n288), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n460), .B1(new_n468), .B2(new_n295), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT85), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n275), .A2(new_n286), .ZN(new_n472));
  INV_X1    g0272(.A(G244), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n472), .B(new_n474), .C1(new_n251), .C2(new_n252), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n256), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT84), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(KEYINPUT84), .A3(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n283), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n208), .A2(G45), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n250), .A2(G250), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  AND2_X1   g0286(.A1(G33), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(G274), .B1(new_n487), .B2(new_n294), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n484), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n267), .A2(G1), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n273), .A2(KEYINPUT83), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G200), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n338), .B1(G1), .B2(new_n256), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n483), .A2(G190), .A3(new_n492), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n471), .A2(new_n494), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n468), .A2(new_n295), .ZN(new_n500));
  INV_X1    g0300(.A(new_n460), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n470), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g0302(.A(KEYINPUT85), .B(new_n460), .C1(new_n468), .C2(new_n295), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n502), .A2(new_n503), .B1(new_n495), .B2(new_n412), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n493), .A2(new_n418), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n483), .A2(new_n404), .A3(new_n492), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n356), .A2(KEYINPUT80), .A3(G107), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT79), .B(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n288), .A2(KEYINPUT6), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n288), .A2(new_n398), .A3(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n513), .A3(new_n512), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(G20), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n299), .A2(G77), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT80), .B1(new_n356), .B2(G107), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n295), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n306), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n496), .B2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(new_n286), .C1(new_n251), .C2(new_n252), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT4), .B1(new_n263), .B2(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n283), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(KEYINPUT5), .A2(G41), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT5), .A2(G41), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n490), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT81), .B1(new_n535), .B2(new_n488), .ZN(new_n536));
  OR2_X1    g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n484), .B1(new_n537), .B2(new_n532), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n539), .A3(new_n273), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT5), .B(G41), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n490), .B1(new_n228), .B2(new_n249), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n536), .A2(new_n540), .B1(new_n542), .B2(G257), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT82), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n531), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n536), .A2(new_n540), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(G257), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n546), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n418), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n535), .A2(new_n488), .A3(KEYINPUT81), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n539), .B1(new_n538), .B2(new_n273), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n543), .A2(new_n544), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n404), .A4(new_n531), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n524), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n422), .A4(new_n531), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n545), .A2(new_n548), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n557), .B1(new_n558), .B2(G200), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n521), .A2(new_n523), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n508), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n398), .A3(G20), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n565), .C1(new_n476), .C2(new_n296), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n256), .A2(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G116), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n570), .A2(KEYINPUT87), .A3(new_n565), .A4(new_n563), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n209), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n259), .A2(new_n576), .A3(new_n209), .A4(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n572), .A2(new_n573), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n572), .B2(new_n578), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n295), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT25), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n306), .B2(G107), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n306), .A2(new_n582), .A3(G107), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n496), .A2(G107), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G257), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G1698), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G250), .B2(G1698), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n251), .A2(new_n252), .ZN(new_n591));
  INV_X1    g0391(.A(G294), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n590), .A2(new_n591), .B1(new_n256), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n283), .B1(new_n542), .B2(G264), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(KEYINPUT88), .A3(G179), .A4(new_n546), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n283), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n542), .A2(G264), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n546), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(G169), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n404), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n550), .A2(new_n551), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n286), .A2(G264), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G257), .A2(G1698), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(new_n251), .B2(new_n252), .ZN(new_n607));
  INV_X1    g0407(.A(G303), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n257), .A2(new_n608), .A3(new_n258), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n283), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n535), .A2(G270), .A3(new_n250), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n604), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n307), .A2(new_n476), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n293), .A2(new_n294), .B1(G20), .B2(new_n476), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n526), .B(new_n209), .C1(G33), .C2(new_n288), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n615), .A2(KEYINPUT20), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT20), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n476), .B1(new_n208), .B2(G33), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n313), .A2(new_n314), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n250), .B1(new_n591), .B2(new_n608), .ZN(new_n624));
  AOI22_X1  g0424(.A1(G270), .A2(new_n542), .B1(new_n624), .B2(new_n607), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n546), .A3(new_n385), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n613), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT86), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n613), .A2(new_n623), .A3(new_n626), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n621), .B(new_n614), .C1(new_n618), .C2(new_n617), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n611), .B(new_n610), .C1(new_n550), .C2(new_n551), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT21), .A4(G169), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n632), .A2(G179), .A3(new_n546), .A4(new_n625), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n418), .B1(new_n625), .B2(new_n546), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT21), .B1(new_n637), .B2(new_n632), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n599), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n599), .A2(G190), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n581), .B(new_n586), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n603), .A2(new_n631), .A3(new_n639), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n459), .A2(new_n562), .A3(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n456), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n388), .A2(new_n392), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n420), .B1(new_n322), .B2(new_n324), .ZN(new_n648));
  INV_X1    g0448(.A(new_n333), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT92), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n374), .B2(new_n375), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n359), .A2(new_n373), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n389), .A2(new_n339), .B1(new_n366), .B2(new_n372), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT18), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n657), .A3(KEYINPUT92), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n650), .A2(new_n652), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n646), .B1(new_n659), .B2(new_n447), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n524), .A2(new_n549), .A3(new_n555), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n508), .A2(new_n661), .A3(KEYINPUT26), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n499), .A2(new_n507), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n556), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n507), .A2(KEYINPUT90), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n504), .A2(new_n505), .A3(new_n668), .A4(new_n506), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT91), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n670), .B1(new_n662), .B2(new_n665), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n603), .B(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n636), .A2(new_n638), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n404), .A2(new_n558), .B1(new_n521), .B2(new_n523), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(new_n549), .B1(new_n559), .B2(new_n560), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n682), .A2(new_n508), .A3(new_n643), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n673), .A2(new_n676), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n660), .B1(new_n459), .B2(new_n684), .ZN(G369));
  NAND3_X1  g0485(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n632), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT93), .Z(new_n693));
  AND2_X1   g0493(.A1(new_n631), .A2(new_n639), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT94), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n639), .ZN(new_n698));
  OAI21_X1  g0498(.A(G330), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n587), .A2(new_n691), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n603), .A2(new_n700), .A3(new_n643), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n587), .A2(new_n602), .A3(new_n691), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n691), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n679), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n603), .A2(new_n643), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n691), .B(KEYINPUT95), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n678), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n706), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n212), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n463), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n226), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n712), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n553), .A2(new_n554), .A3(new_n531), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n483), .A2(new_n492), .A3(new_n594), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n625), .A2(G179), .A3(new_n546), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n725), .A2(new_n726), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(new_n558), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n724), .A2(new_n599), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT97), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G238), .A2(G1698), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n473), .B2(G1698), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n477), .B1(new_n735), .B2(new_n259), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n283), .B1(new_n736), .B2(KEYINPUT84), .ZN(new_n737));
  INV_X1    g0537(.A(new_n482), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT96), .B(new_n492), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n625), .B2(new_n546), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT96), .B1(new_n483), .B2(new_n492), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n733), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n493), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(KEYINPUT97), .A3(new_n739), .A4(new_n740), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n732), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n723), .B1(new_n731), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n743), .A2(new_n746), .ZN(new_n749));
  INV_X1    g0549(.A(new_n732), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n483), .A2(new_n492), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n633), .A2(new_n404), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n594), .ZN(new_n754));
  OAI21_X1  g0554(.A(KEYINPUT30), .B1(new_n754), .B2(new_n724), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n558), .A2(new_n729), .A3(new_n728), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n707), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n748), .B1(new_n758), .B2(KEYINPUT31), .ZN(new_n759));
  INV_X1    g0559(.A(new_n712), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n562), .A2(new_n644), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(G330), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT98), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND4_X1   g0564(.A1(new_n603), .A2(new_n631), .A3(new_n639), .A4(new_n643), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(new_n682), .A3(new_n508), .A4(new_n712), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n749), .A2(new_n750), .B1(new_n755), .B2(new_n756), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n722), .B1(new_n767), .B2(new_n707), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n768), .A3(new_n748), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT98), .A3(G330), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT99), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n684), .B2(new_n760), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT29), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n683), .B1(new_n679), .B2(new_n678), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n675), .B1(new_n666), .B2(new_n671), .ZN(new_n776));
  AOI211_X1 g0576(.A(KEYINPUT91), .B(new_n670), .C1(new_n662), .C2(new_n665), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(KEYINPUT99), .A3(new_n712), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n773), .A2(new_n774), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n603), .A2(new_n639), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n683), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n691), .B1(new_n782), .B2(new_n674), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT29), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n771), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n721), .B1(new_n785), .B2(G1), .ZN(G364));
  AOI21_X1  g0586(.A(new_n294), .B1(G20), .B2(new_n418), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n422), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n209), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n209), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n789), .A2(new_n592), .B1(new_n791), .B2(new_n608), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n790), .A2(new_n422), .A3(new_n320), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n259), .B1(new_n794), .B2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n790), .A2(new_n422), .A3(G200), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(G20), .A2(G179), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(G200), .A3(new_n385), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n792), .B(new_n798), .C1(G326), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(new_n422), .A3(new_n320), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n800), .A2(new_n422), .A3(G200), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT33), .B(G317), .Z(new_n807));
  OAI221_X1 g0607(.A(new_n803), .B1(new_n804), .B2(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n800), .A2(new_n320), .A3(new_n385), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT101), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n809), .A2(KEYINPUT101), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n808), .B1(G322), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n794), .A2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(new_n789), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(KEYINPUT32), .B1(G97), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(KEYINPUT32), .B2(new_n816), .C1(new_n398), .C2(new_n797), .ZN(new_n819));
  INV_X1    g0619(.A(new_n805), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(G77), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n791), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G87), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n259), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(KEYINPUT102), .ZN(new_n825));
  INV_X1    g0625(.A(new_n806), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G68), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n802), .A2(G50), .B1(new_n824), .B2(KEYINPUT102), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n821), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G58), .B2(new_n814), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n787), .B1(new_n815), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n209), .A2(G13), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n208), .B1(new_n832), .B2(G45), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n716), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n715), .A2(new_n259), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n267), .B2(new_n227), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n267), .B2(new_n243), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n715), .A2(new_n591), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n841), .A2(G355), .B1(new_n476), .B2(new_n715), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(G13), .A2(G33), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(G20), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n787), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n836), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n831), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n697), .A2(new_n698), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n699), .A2(new_n836), .ZN(new_n852));
  INV_X1    g0652(.A(G330), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G396));
  OAI22_X1  g0656(.A1(new_n421), .A2(new_n423), .B1(new_n417), .B2(new_n707), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n420), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n405), .A2(new_n419), .A3(new_n707), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n773), .A2(new_n779), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n778), .A2(new_n712), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n771), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT106), .Z(new_n867));
  NAND2_X1  g0667(.A1(new_n864), .A2(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n836), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G137), .A2(new_n802), .B1(new_n820), .B2(G159), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n431), .B2(new_n806), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G143), .B2(new_n814), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT34), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(KEYINPUT34), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n817), .A2(G58), .B1(new_n822), .B2(G50), .ZN(new_n875));
  INV_X1    g0675(.A(new_n797), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(G68), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n591), .B1(new_n794), .B2(G132), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n873), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n591), .B1(new_n791), .B2(new_n398), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT104), .Z(new_n882));
  OAI22_X1  g0682(.A1(new_n476), .A2(new_n805), .B1(new_n806), .B2(new_n796), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n797), .A2(new_n407), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n789), .A2(new_n288), .B1(new_n793), .B2(new_n804), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n802), .C2(G303), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n884), .B(new_n887), .C1(new_n592), .C2(new_n813), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  INV_X1    g0693(.A(new_n787), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n787), .A2(new_n844), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n835), .B1(G77), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n898), .B(KEYINPUT103), .Z(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n862), .B2(new_n845), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n867), .A2(new_n869), .B1(new_n895), .B2(new_n900), .ZN(G384));
  NOR3_X1   g0701(.A1(new_n294), .A2(new_n209), .A3(new_n476), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n515), .A2(new_n516), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT35), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n226), .A2(new_n205), .A3(new_n347), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n202), .A2(G68), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n208), .B(G13), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n751), .A2(new_n757), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n766), .A2(new_n914), .A3(new_n768), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n862), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n326), .A2(new_n691), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n331), .A2(new_n332), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n917), .B1(new_n325), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n325), .A2(new_n333), .A3(new_n917), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n325), .A2(new_n333), .A3(KEYINPUT108), .A4(new_n917), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n916), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n689), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n359), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n653), .A2(new_n927), .A3(new_n390), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT37), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n390), .A2(KEYINPUT37), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n339), .B1(new_n353), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n373), .B2(new_n926), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n926), .B(new_n933), .C1(new_n376), .C2(new_n393), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n933), .A2(new_n926), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n655), .A2(new_n657), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n940), .B1(new_n647), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n930), .A2(new_n935), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n942), .A2(new_n943), .A3(new_n939), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n652), .A2(new_n658), .A3(new_n647), .ZN(new_n948));
  INV_X1    g0748(.A(new_n927), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n927), .A2(new_n390), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n927), .A2(new_n651), .A3(new_n390), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(new_n653), .B1(new_n953), .B2(KEYINPUT37), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n951), .A2(new_n651), .A3(new_n929), .A4(new_n656), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n947), .B1(new_n957), .B2(new_n939), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n958), .A2(new_n916), .A3(new_n924), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT40), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n946), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT109), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n458), .A2(new_n915), .ZN(new_n963));
  OAI21_X1  g0763(.A(G330), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n780), .A2(new_n458), .A3(new_n784), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n660), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n652), .A2(new_n658), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n689), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n938), .A2(new_n944), .A3(KEYINPUT39), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n958), .B2(KEYINPUT39), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n649), .A2(new_n707), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n938), .A2(new_n944), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n859), .B(KEYINPUT107), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n924), .B1(new_n863), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n973), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n967), .B(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n965), .A2(new_n979), .B1(new_n208), .B2(new_n832), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n965), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n912), .B1(new_n980), .B2(new_n981), .ZN(G367));
  OAI21_X1  g0782(.A(new_n847), .B1(new_n212), .B2(new_n412), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n837), .B2(new_n239), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT111), .Z(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n591), .B1(new_n793), .B2(new_n986), .C1(new_n288), .C2(new_n797), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n791), .A2(new_n476), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT46), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G107), .C2(new_n817), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n796), .A2(new_n805), .B1(new_n806), .B2(new_n592), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G311), .B2(new_n802), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(new_n608), .C2(new_n813), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n789), .A2(new_n308), .B1(new_n797), .B2(new_n205), .ZN(new_n994));
  INV_X1    g0794(.A(G137), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n259), .B1(new_n793), .B2(new_n995), .C1(new_n346), .C2(new_n791), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(G143), .C2(new_n802), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G50), .A2(new_n820), .B1(new_n826), .B2(G159), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(new_n431), .C2(new_n813), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n836), .B(new_n985), .C1(new_n1001), .C2(new_n787), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n846), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n471), .A2(new_n497), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n691), .ZN(new_n1005));
  MUX2_X1   g0805(.A(new_n671), .B(new_n664), .S(new_n1005), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1002), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT112), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n682), .B1(new_n560), .B2(new_n712), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n556), .B2(new_n712), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1014), .A2(KEYINPUT110), .A3(new_n711), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT110), .B1(new_n1014), .B2(new_n711), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1015), .A2(new_n1016), .A3(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n556), .B1(new_n1013), .B2(new_n603), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n712), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT42), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1012), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n705), .A2(new_n1014), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n713), .A2(new_n1014), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT45), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT44), .ZN(new_n1032));
  OR3_X1    g0832(.A1(new_n713), .A2(new_n1032), .A3(new_n1014), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n713), .B2(new_n1014), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n705), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1031), .A2(new_n706), .A3(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n704), .A2(new_n708), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n710), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n699), .B(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n785), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n716), .B(KEYINPUT41), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n834), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1010), .B1(new_n1028), .B2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n718), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n841), .A2(new_n1048), .B1(new_n398), .B2(new_n715), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n236), .A2(new_n267), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n336), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n202), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n718), .B(new_n267), .C1(new_n308), .C2(new_n205), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n837), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1049), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n836), .B1(new_n1056), .B2(new_n847), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n703), .B2(new_n1003), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n806), .A2(new_n336), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n259), .B1(new_n793), .B2(new_n431), .C1(new_n288), .C2(new_n797), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n789), .A2(new_n412), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n791), .A2(new_n205), .ZN(new_n1062));
  NOR4_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G68), .A2(new_n820), .B1(new_n802), .B2(G159), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n202), .C2(new_n813), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n259), .B1(new_n794), .B2(G326), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n789), .A2(new_n796), .B1(new_n791), .B2(new_n592), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n608), .A2(new_n805), .B1(new_n806), .B2(new_n804), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G322), .B2(new_n802), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n813), .B2(new_n986), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT49), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1066), .B1(new_n476), .B2(new_n797), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1065), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1058), .B1(new_n1077), .B2(new_n787), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT113), .Z(new_n1079));
  INV_X1    g0879(.A(new_n1042), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n834), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n717), .B1(new_n785), .B2(new_n1080), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT114), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1082), .A2(new_n1083), .B1(new_n785), .B2(new_n1080), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(G393));
  NAND3_X1  g0886(.A1(new_n1037), .A2(new_n834), .A3(new_n1038), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n847), .B1(new_n288), .B2(new_n212), .C1(new_n838), .C2(new_n246), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n835), .ZN(new_n1089));
  INV_X1    g0889(.A(G159), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n813), .A2(new_n1090), .B1(new_n431), .B2(new_n801), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  AOI211_X1 g0892(.A(new_n591), .B(new_n885), .C1(G143), .C2(new_n794), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n817), .A2(G77), .B1(new_n822), .B2(G68), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n202), .B2(new_n806), .C1(new_n336), .C2(new_n805), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n813), .A2(new_n804), .B1(new_n986), .B2(new_n801), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  NOR2_X1   g0898(.A1(new_n797), .A2(new_n398), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n259), .B(new_n1099), .C1(G322), .C2(new_n794), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n817), .A2(G116), .B1(new_n822), .B2(G283), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n592), .B2(new_n805), .C1(new_n608), .C2(new_n806), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1092), .A2(new_n1096), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n1104), .B2(new_n787), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1014), .B2(new_n1003), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1087), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT115), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1087), .A2(new_n1109), .A3(new_n1106), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n785), .A2(new_n1080), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1039), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n716), .B1(new_n1039), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(G390));
  NAND2_X1  g0915(.A1(new_n863), .A2(new_n976), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n691), .B1(new_n731), .B2(new_n747), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(new_n722), .B1(new_n913), .B2(new_n723), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n763), .B(new_n853), .C1(new_n1118), .C2(new_n766), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT98), .B1(new_n769), .B2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n862), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(KEYINPUT116), .A3(new_n924), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n916), .A2(new_n853), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n922), .A2(new_n923), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n919), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT116), .B1(new_n1121), .B2(new_n924), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1116), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n975), .B1(new_n783), .B2(new_n862), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n860), .B1(new_n764), .B2(new_n770), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1132), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n458), .A2(G330), .A3(new_n915), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n966), .A2(new_n660), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n972), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n971), .B1(new_n977), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1133), .A2(new_n1126), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n957), .A2(new_n939), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n938), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n972), .B(new_n1144), .C1(new_n1131), .C2(new_n924), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1127), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1136), .A2(new_n1139), .A3(new_n1146), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT116), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1134), .B1(new_n1153), .B2(new_n1116), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1127), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1154), .A2(new_n1138), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1150), .A2(new_n716), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT119), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1155), .A2(new_n1156), .A3(new_n833), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G107), .A2(new_n826), .B1(new_n802), .B2(G283), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n288), .B2(new_n805), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT117), .Z(new_n1163));
  AOI21_X1  g0963(.A(new_n259), .B1(new_n794), .B2(G294), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n817), .A2(G77), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n1165), .A3(new_n823), .A4(new_n877), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n814), .B2(G116), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n814), .A2(G132), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n591), .B1(new_n794), .B2(G125), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n202), .B2(new_n797), .C1(new_n1090), .C2(new_n789), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n802), .A2(G128), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n791), .A2(new_n431), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n995), .C2(new_n806), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT54), .B(G143), .Z(new_n1175));
  AOI211_X1 g0975(.A(new_n1170), .B(new_n1174), .C1(new_n820), .C2(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1163), .A2(new_n1167), .B1(new_n1168), .B2(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n835), .B1(new_n1051), .B2(new_n897), .C1(new_n1177), .C2(new_n894), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n971), .B2(new_n844), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT118), .Z(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1159), .B1(new_n1160), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1149), .A2(new_n1146), .ZN(new_n1183));
  OAI211_X1 g0983(.A(KEYINPUT119), .B(new_n1180), .C1(new_n1183), .C2(new_n833), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1158), .A2(new_n1182), .A3(new_n1184), .ZN(G378));
  NOR2_X1   g0985(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1138), .B1(new_n1186), .B2(new_n1136), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n977), .A2(new_n974), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n969), .C1(new_n972), .C2(new_n971), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n438), .A2(new_n926), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT55), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n457), .A2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1194));
  NAND3_X1  g0994(.A1(new_n447), .A2(new_n456), .A3(new_n1191), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n915), .A2(new_n862), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1126), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT40), .B1(new_n1200), .B2(new_n958), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n853), .B(new_n1198), .C1(new_n1201), .C2(new_n946), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n961), .B2(G330), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1189), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1144), .A2(new_n1126), .A3(new_n1199), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n1206), .A2(KEYINPUT40), .B1(new_n925), .B2(new_n945), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1198), .B1(new_n1207), .B2(new_n853), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n961), .A2(G330), .A3(new_n1203), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n978), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(KEYINPUT57), .A3(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n716), .B1(new_n1187), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1139), .B1(new_n1183), .B2(new_n1154), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1210), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n978), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(KEYINPUT57), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1205), .A2(new_n834), .A3(new_n1210), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n814), .A2(G107), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n802), .A2(G116), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n266), .B(new_n591), .C1(new_n793), .C2(new_n796), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n789), .A2(new_n308), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n797), .A2(new_n346), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1062), .A4(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G97), .A2(new_n826), .B1(new_n820), .B2(new_n411), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1220), .A2(new_n1221), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n591), .A2(new_n266), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G50), .B1(new_n256), .B2(new_n266), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1227), .A2(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G132), .A2(new_n826), .B1(new_n820), .B2(G137), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n802), .A2(G125), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n817), .A2(G150), .B1(new_n822), .B2(new_n1175), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G128), .B2(new_n814), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n876), .A2(G159), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1237), .A2(KEYINPUT59), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1231), .B1(new_n1228), .B2(new_n1227), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n787), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n836), .B1(new_n202), .B2(new_n896), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(new_n1198), .C2(new_n845), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1219), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1218), .A2(new_n1248), .ZN(G375));
  NAND2_X1  g1049(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1154), .A2(new_n1138), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1045), .A3(new_n1251), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n789), .A2(new_n412), .B1(new_n791), .B2(new_n288), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n591), .B1(new_n793), .B2(new_n608), .C1(new_n205), .C2(new_n797), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(G107), .C2(new_n820), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G116), .A2(new_n826), .B1(new_n802), .B2(G294), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(new_n796), .C2(new_n813), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n591), .B(new_n1224), .C1(G128), .C2(new_n794), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n817), .A2(G50), .B1(new_n822), .B2(G159), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1258), .B(new_n1259), .C1(new_n431), .C2(new_n805), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT121), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G132), .A2(new_n802), .B1(new_n826), .B2(new_n1175), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n813), .B2(new_n995), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1257), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n787), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n836), .B1(new_n308), .B2(new_n896), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1265), .B(new_n1266), .C1(new_n1126), .C2(new_n845), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1136), .B2(new_n834), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1252), .A2(new_n1269), .ZN(G381));
  OAI211_X1 g1070(.A(new_n855), .B(new_n1081), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G384), .A2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT122), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1160), .A2(new_n1181), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1158), .A2(new_n1274), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G387), .A2(G390), .A3(new_n1275), .A4(G381), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1273), .A2(new_n1276), .A3(G375), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT123), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1279), .A2(new_n1280), .ZN(G407));
  OAI21_X1  g1081(.A(new_n1180), .B1(new_n1183), .B2(new_n833), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n717), .B1(new_n1250), .B2(new_n1183), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1150), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n690), .ZN(new_n1285));
  OAI221_X1 g1085(.A(G213), .B1(G375), .B2(new_n1285), .C1(new_n1279), .C2(new_n1280), .ZN(G409));
  NAND2_X1  g1086(.A1(G393), .A2(G396), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1271), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(G387), .A2(G390), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G390), .A2(new_n1290), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1111), .B(KEYINPUT125), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1289), .B(new_n1291), .C1(new_n1294), .C2(G387), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G390), .ZN(new_n1298));
  INV_X1    g1098(.A(G390), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1299), .A2(new_n1296), .A3(G387), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1300), .A3(new_n1288), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1248), .C1(new_n1217), .C2(new_n1212), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1205), .A2(new_n1045), .A3(new_n1210), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1247), .B1(new_n1213), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1305), .B1(new_n1308), .B2(new_n1275), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1219), .B(new_n1246), .C1(new_n1187), .C2(new_n1306), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1284), .A2(new_n1310), .A3(KEYINPUT124), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1304), .A2(new_n1309), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1154), .A2(new_n1138), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1251), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1154), .A2(KEYINPUT60), .A3(new_n1138), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1315), .A2(new_n716), .A3(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1317), .A2(G384), .A3(new_n1269), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1317), .B2(new_n1269), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n690), .A2(G213), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1312), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1312), .A2(new_n1325), .A3(new_n1321), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1312), .B2(new_n1321), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NOR3_X1   g1128(.A1(new_n1318), .A2(new_n1319), .A3(new_n1323), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1324), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(G2897), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1321), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1320), .A2(new_n1332), .ZN(new_n1333));
  OAI22_X1  g1133(.A1(new_n1318), .A2(new_n1319), .B1(new_n1331), .B2(new_n1321), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1335), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1303), .B1(new_n1330), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1302), .A2(new_n1337), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1312), .A2(new_n1321), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1341), .B2(new_n1335), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1320), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1322), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1342), .A2(new_n1343), .A3(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1339), .A2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1284), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1304), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1303), .A2(new_n1349), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1302), .A2(new_n1304), .A3(new_n1348), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1320), .ZN(G402));
endmodule


