

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U566 ( .A1(n536), .A2(G2105), .ZN(n894) );
  NOR2_X1 U567 ( .A1(n808), .A2(n790), .ZN(n791) );
  NOR2_X2 U568 ( .A1(G2105), .A2(n536), .ZN(n887) );
  NOR2_X2 U569 ( .A1(n545), .A2(n544), .ZN(G160) );
  NOR2_X1 U570 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U571 ( .A1(n732), .A2(n731), .ZN(n733) );
  OR2_X1 U572 ( .A1(n996), .A2(n734), .ZN(n741) );
  INV_X1 U573 ( .A(KEYINPUT97), .ZN(n742) );
  XNOR2_X1 U574 ( .A(n743), .B(n742), .ZN(n749) );
  NOR2_X1 U575 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U576 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U577 ( .A1(G651), .A2(n646), .ZN(n659) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n553), .Z(n658) );
  INV_X1 U579 ( .A(G2104), .ZN(n536) );
  NAND2_X1 U580 ( .A1(G125), .A2(n894), .ZN(n535) );
  XNOR2_X1 U581 ( .A(n535), .B(KEYINPUT64), .ZN(n539) );
  NAND2_X1 U582 ( .A1(G101), .A2(n887), .ZN(n537) );
  XOR2_X1 U583 ( .A(n537), .B(KEYINPUT23), .Z(n538) );
  NAND2_X1 U584 ( .A1(n539), .A2(n538), .ZN(n545) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U586 ( .A1(G113), .A2(n891), .ZN(n543) );
  XNOR2_X1 U587 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n541) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  XNOR2_X2 U589 ( .A(n541), .B(n540), .ZN(n886) );
  NAND2_X1 U590 ( .A1(G137), .A2(n886), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U592 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U593 ( .A1(G89), .A2(n653), .ZN(n546) );
  XNOR2_X1 U594 ( .A(n546), .B(KEYINPUT4), .ZN(n547) );
  XNOR2_X1 U595 ( .A(KEYINPUT76), .B(n547), .ZN(n550) );
  XOR2_X1 U596 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  INV_X1 U597 ( .A(G651), .ZN(n552) );
  NOR2_X2 U598 ( .A1(n646), .A2(n552), .ZN(n654) );
  NAND2_X1 U599 ( .A1(n654), .A2(G76), .ZN(n548) );
  XOR2_X1 U600 ( .A(KEYINPUT77), .B(n548), .Z(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U602 ( .A(n551), .B(KEYINPUT5), .ZN(n558) );
  NOR2_X1 U603 ( .A1(G543), .A2(n552), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G63), .A2(n658), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G51), .A2(n659), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U608 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U609 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G64), .A2(n658), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G52), .A2(n659), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U614 ( .A1(G90), .A2(n653), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G77), .A2(n654), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U617 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U618 ( .A1(n566), .A2(n565), .ZN(G171) );
  NAND2_X1 U619 ( .A1(G88), .A2(n653), .ZN(n568) );
  NAND2_X1 U620 ( .A1(G62), .A2(n658), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U622 ( .A1(G75), .A2(n654), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G50), .A2(n659), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U626 ( .A(KEYINPUT85), .B(n573), .Z(G166) );
  INV_X1 U627 ( .A(G166), .ZN(G303) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U629 ( .A(G57), .ZN(G237) );
  INV_X1 U630 ( .A(G132), .ZN(G219) );
  INV_X1 U631 ( .A(G82), .ZN(G220) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U633 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U634 ( .A(G223), .ZN(n836) );
  NAND2_X1 U635 ( .A1(n836), .A2(G567), .ZN(n575) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n658), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n576), .Z(n584) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(KEYINPUT12), .Z(n578) );
  NAND2_X1 U640 ( .A1(G81), .A2(n653), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n578), .B(n577), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n654), .A2(G68), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT13), .ZN(n583) );
  NOR2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U646 ( .A1(n659), .A2(G43), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n586), .A2(n585), .ZN(n983) );
  INV_X1 U648 ( .A(G860), .ZN(n611) );
  OR2_X1 U649 ( .A1(n983), .A2(n611), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U652 ( .A1(n659), .A2(G54), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT74), .ZN(n589) );
  NAND2_X1 U654 ( .A1(G79), .A2(n654), .ZN(n588) );
  NAND2_X1 U655 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U657 ( .A1(G92), .A2(n653), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT73), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G66), .A2(n658), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U661 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X2 U663 ( .A(n597), .B(KEYINPUT15), .ZN(n996) );
  OR2_X1 U664 ( .A1(n996), .A2(G868), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G65), .A2(n658), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G53), .A2(n659), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(KEYINPUT69), .B(n602), .ZN(n608) );
  NAND2_X1 U670 ( .A1(G91), .A2(n653), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT67), .ZN(n606) );
  NAND2_X1 U672 ( .A1(G78), .A2(n654), .ZN(n604) );
  XOR2_X1 U673 ( .A(KEYINPUT68), .B(n604), .Z(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n608), .A2(n607), .ZN(G299) );
  INV_X1 U676 ( .A(G868), .ZN(n672) );
  NOR2_X1 U677 ( .A1(G286), .A2(n672), .ZN(n610) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n611), .A2(G559), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n612), .A2(n996), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n996), .A2(G868), .ZN(n614) );
  NOR2_X1 U684 ( .A1(G559), .A2(n614), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT78), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n983), .A2(G868), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n894), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  XNOR2_X1 U690 ( .A(n619), .B(KEYINPUT79), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G111), .A2(n891), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G135), .A2(n886), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G99), .A2(n887), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n935) );
  XOR2_X1 U697 ( .A(n935), .B(G2096), .Z(n627) );
  XNOR2_X1 U698 ( .A(G2100), .B(KEYINPUT80), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT81), .B(n628), .ZN(G156) );
  NAND2_X1 U701 ( .A1(n996), .A2(G559), .ZN(n670) );
  XNOR2_X1 U702 ( .A(n983), .B(n670), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n629), .A2(G860), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G67), .A2(n658), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G55), .A2(n659), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G93), .A2(n653), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G80), .A2(n654), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n673) );
  XOR2_X1 U711 ( .A(n636), .B(n673), .Z(G145) );
  NAND2_X1 U712 ( .A1(n659), .A2(G48), .ZN(n637) );
  XNOR2_X1 U713 ( .A(KEYINPUT84), .B(n637), .ZN(n645) );
  NAND2_X1 U714 ( .A1(G86), .A2(n653), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G61), .A2(n658), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n654), .A2(G73), .ZN(n640) );
  XOR2_X1 U718 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT83), .B(n643), .Z(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U723 ( .A1(G49), .A2(n659), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G87), .A2(n646), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n658), .A2(n649), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U729 ( .A1(G85), .A2(n653), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G72), .A2(n654), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U732 ( .A(KEYINPUT66), .B(n657), .Z(n663) );
  NAND2_X1 U733 ( .A1(G60), .A2(n658), .ZN(n661) );
  NAND2_X1 U734 ( .A1(G47), .A2(n659), .ZN(n660) );
  AND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(G290) );
  INV_X1 U737 ( .A(G299), .ZN(n986) );
  XNOR2_X1 U738 ( .A(n986), .B(KEYINPUT19), .ZN(n664) );
  XOR2_X1 U739 ( .A(n664), .B(n673), .Z(n667) );
  XNOR2_X1 U740 ( .A(G288), .B(G290), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(G303), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U743 ( .A(n668), .B(n983), .ZN(n669) );
  XNOR2_X1 U744 ( .A(G305), .B(n669), .ZN(n908) );
  XOR2_X1 U745 ( .A(n908), .B(n670), .Z(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(n675) );
  NOR2_X1 U747 ( .A1(G868), .A2(n673), .ZN(n674) );
  NOR2_X1 U748 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U758 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U759 ( .A1(G96), .A2(n683), .ZN(n841) );
  NAND2_X1 U760 ( .A1(n841), .A2(G2106), .ZN(n687) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U762 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G108), .A2(n685), .ZN(n842) );
  NAND2_X1 U764 ( .A1(n842), .A2(G567), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n687), .A2(n686), .ZN(n843) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U767 ( .A1(n843), .A2(n688), .ZN(n840) );
  NAND2_X1 U768 ( .A1(n840), .A2(G36), .ZN(n689) );
  XOR2_X1 U769 ( .A(KEYINPUT87), .B(n689), .Z(G176) );
  NAND2_X1 U770 ( .A1(G126), .A2(n894), .ZN(n691) );
  NAND2_X1 U771 ( .A1(G114), .A2(n891), .ZN(n690) );
  NAND2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U773 ( .A(KEYINPUT88), .B(n692), .ZN(n696) );
  NAND2_X1 U774 ( .A1(G138), .A2(n886), .ZN(n694) );
  NAND2_X1 U775 ( .A1(G102), .A2(n887), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U777 ( .A1(n696), .A2(n695), .ZN(G164) );
  XNOR2_X1 U778 ( .A(G1986), .B(G290), .ZN(n985) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n830) );
  NAND2_X1 U782 ( .A1(n985), .A2(n830), .ZN(n818) );
  NAND2_X1 U783 ( .A1(G140), .A2(n886), .ZN(n698) );
  NAND2_X1 U784 ( .A1(G104), .A2(n887), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n699), .ZN(n704) );
  NAND2_X1 U787 ( .A1(G128), .A2(n894), .ZN(n701) );
  NAND2_X1 U788 ( .A1(G116), .A2(n891), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U790 ( .A(n702), .B(KEYINPUT35), .Z(n703) );
  NOR2_X1 U791 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U792 ( .A(KEYINPUT36), .B(n705), .Z(n706) );
  XNOR2_X1 U793 ( .A(KEYINPUT89), .B(n706), .ZN(n904) );
  XNOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U795 ( .A1(n904), .A2(n819), .ZN(n934) );
  NAND2_X1 U796 ( .A1(n830), .A2(n934), .ZN(n827) );
  NAND2_X1 U797 ( .A1(G119), .A2(n894), .ZN(n708) );
  NAND2_X1 U798 ( .A1(G107), .A2(n891), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n713) );
  NAND2_X1 U800 ( .A1(G131), .A2(n886), .ZN(n710) );
  NAND2_X1 U801 ( .A1(G95), .A2(n887), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U803 ( .A(KEYINPUT90), .B(n711), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U805 ( .A(n714), .B(KEYINPUT91), .Z(n899) );
  INV_X1 U806 ( .A(G1991), .ZN(n960) );
  NOR2_X1 U807 ( .A1(n899), .A2(n960), .ZN(n723) );
  NAND2_X1 U808 ( .A1(G129), .A2(n894), .ZN(n716) );
  NAND2_X1 U809 ( .A1(G141), .A2(n886), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n887), .A2(G105), .ZN(n717) );
  XOR2_X1 U812 ( .A(KEYINPUT38), .B(n717), .Z(n718) );
  NOR2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n891), .A2(G117), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n871) );
  AND2_X1 U816 ( .A1(n871), .A2(G1996), .ZN(n722) );
  NOR2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n932) );
  INV_X1 U818 ( .A(n830), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n932), .A2(n724), .ZN(n823) );
  INV_X1 U820 ( .A(n823), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n827), .A2(n725), .ZN(n726) );
  XNOR2_X1 U822 ( .A(n726), .B(KEYINPUT92), .ZN(n816) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n998) );
  INV_X1 U824 ( .A(n727), .ZN(n729) );
  NAND2_X2 U825 ( .A1(n729), .A2(n728), .ZN(n771) );
  NAND2_X1 U826 ( .A1(G8), .A2(n771), .ZN(n808) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n988) );
  INV_X1 U828 ( .A(G1996), .ZN(n954) );
  NOR2_X1 U829 ( .A1(n771), .A2(n954), .ZN(n730) );
  XNOR2_X1 U830 ( .A(n730), .B(KEYINPUT26), .ZN(n732) );
  AND2_X1 U831 ( .A1(n771), .A2(G1341), .ZN(n731) );
  NOR2_X1 U832 ( .A1(n983), .A2(n733), .ZN(n734) );
  NAND2_X1 U833 ( .A1(n996), .A2(n734), .ZN(n739) );
  INV_X1 U834 ( .A(G2067), .ZN(n961) );
  NOR2_X1 U835 ( .A1(n771), .A2(n961), .ZN(n735) );
  XOR2_X1 U836 ( .A(n735), .B(KEYINPUT96), .Z(n737) );
  NAND2_X1 U837 ( .A1(n771), .A2(G1348), .ZN(n736) );
  NAND2_X1 U838 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U839 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U840 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n771), .A2(G1956), .ZN(n746) );
  INV_X1 U842 ( .A(n771), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n757), .A2(G2072), .ZN(n744) );
  XOR2_X1 U844 ( .A(KEYINPUT27), .B(n744), .Z(n745) );
  NAND2_X1 U845 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U846 ( .A(n747), .B(KEYINPUT95), .ZN(n750) );
  NAND2_X1 U847 ( .A1(n750), .A2(n986), .ZN(n748) );
  NAND2_X1 U848 ( .A1(n749), .A2(n748), .ZN(n753) );
  NOR2_X1 U849 ( .A1(n750), .A2(n986), .ZN(n751) );
  XOR2_X1 U850 ( .A(n751), .B(KEYINPUT28), .Z(n752) );
  NAND2_X1 U851 ( .A1(n753), .A2(n752), .ZN(n755) );
  XOR2_X1 U852 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n754) );
  XNOR2_X1 U853 ( .A(n755), .B(n754), .ZN(n761) );
  INV_X1 U854 ( .A(G1961), .ZN(n1030) );
  NAND2_X1 U855 ( .A1(n771), .A2(n1030), .ZN(n759) );
  XNOR2_X1 U856 ( .A(G2078), .B(KEYINPUT25), .ZN(n756) );
  XNOR2_X1 U857 ( .A(n756), .B(KEYINPUT94), .ZN(n955) );
  NAND2_X1 U858 ( .A1(n757), .A2(n955), .ZN(n758) );
  NAND2_X1 U859 ( .A1(n759), .A2(n758), .ZN(n765) );
  NAND2_X1 U860 ( .A1(n765), .A2(G171), .ZN(n760) );
  NAND2_X1 U861 ( .A1(n761), .A2(n760), .ZN(n770) );
  NOR2_X1 U862 ( .A1(G1966), .A2(n808), .ZN(n783) );
  NOR2_X1 U863 ( .A1(G2084), .A2(n771), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n783), .A2(n779), .ZN(n762) );
  NAND2_X1 U865 ( .A1(G8), .A2(n762), .ZN(n763) );
  XNOR2_X1 U866 ( .A(KEYINPUT30), .B(n763), .ZN(n764) );
  NOR2_X1 U867 ( .A1(G168), .A2(n764), .ZN(n767) );
  NOR2_X1 U868 ( .A1(G171), .A2(n765), .ZN(n766) );
  NOR2_X1 U869 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U870 ( .A(KEYINPUT31), .B(n768), .Z(n769) );
  NAND2_X1 U871 ( .A1(n770), .A2(n769), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n781), .A2(G286), .ZN(n776) );
  NOR2_X1 U873 ( .A1(G1971), .A2(n808), .ZN(n773) );
  NOR2_X1 U874 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U875 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U876 ( .A1(G303), .A2(n774), .ZN(n775) );
  NAND2_X1 U877 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U878 ( .A1(n777), .A2(G8), .ZN(n778) );
  XNOR2_X1 U879 ( .A(n778), .B(KEYINPUT32), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G8), .A2(n779), .ZN(n780) );
  XOR2_X1 U881 ( .A(KEYINPUT93), .B(n780), .Z(n785) );
  INV_X1 U882 ( .A(n781), .ZN(n782) );
  NOR2_X1 U883 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U884 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U885 ( .A1(n787), .A2(n786), .ZN(n806) );
  INV_X1 U886 ( .A(G1971), .ZN(n1012) );
  NAND2_X1 U887 ( .A1(G166), .A2(n1012), .ZN(n788) );
  NAND2_X1 U888 ( .A1(n806), .A2(n788), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n988), .A2(n789), .ZN(n790) );
  NAND2_X1 U890 ( .A1(n998), .A2(n791), .ZN(n792) );
  NOR2_X1 U891 ( .A1(KEYINPUT99), .A2(n792), .ZN(n793) );
  NOR2_X1 U892 ( .A1(KEYINPUT33), .A2(n793), .ZN(n800) );
  INV_X1 U893 ( .A(KEYINPUT99), .ZN(n795) );
  NAND2_X1 U894 ( .A1(n988), .A2(KEYINPUT33), .ZN(n794) );
  NAND2_X1 U895 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n988), .A2(KEYINPUT99), .ZN(n796) );
  NAND2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U898 ( .A1(n808), .A2(n798), .ZN(n799) );
  XOR2_X1 U899 ( .A(G1981), .B(G305), .Z(n980) );
  NAND2_X1 U900 ( .A1(n801), .A2(n980), .ZN(n814) );
  NOR2_X1 U901 ( .A1(G1981), .A2(G305), .ZN(n802) );
  XOR2_X1 U902 ( .A(n802), .B(KEYINPUT24), .Z(n803) );
  OR2_X1 U903 ( .A1(n808), .A2(n803), .ZN(n812) );
  NOR2_X1 U904 ( .A1(G2090), .A2(G303), .ZN(n804) );
  NAND2_X1 U905 ( .A1(G8), .A2(n804), .ZN(n805) );
  NAND2_X1 U906 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U907 ( .A(n807), .B(KEYINPUT100), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U909 ( .A(KEYINPUT101), .B(n810), .Z(n811) );
  AND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  AND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n833) );
  AND2_X1 U913 ( .A1(n904), .A2(n819), .ZN(n820) );
  XNOR2_X1 U914 ( .A(KEYINPUT103), .B(n820), .ZN(n942) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n871), .ZN(n928) );
  AND2_X1 U916 ( .A1(n960), .A2(n899), .ZN(n936) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n936), .A2(n821), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n823), .A2(n822), .ZN(n824) );
  NOR2_X1 U920 ( .A1(n928), .A2(n824), .ZN(n825) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n825), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n826), .B(KEYINPUT102), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n942), .A2(n829), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n835) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(KEYINPUT104), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  XOR2_X1 U933 ( .A(KEYINPUT107), .B(n838), .Z(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  INV_X1 U941 ( .A(n843), .ZN(G319) );
  XOR2_X1 U942 ( .A(G2100), .B(G2096), .Z(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(G2678), .B(G2090), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1966), .Z(n853) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1981), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n854), .B(KEYINPUT109), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(G1956), .B(G1961), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1976), .B(G1971), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U961 ( .A(KEYINPUT108), .B(G2474), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U963 ( .A1(n887), .A2(G100), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G112), .A2(n891), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G136), .A2(n886), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n894), .A2(G124), .ZN(n865) );
  XOR2_X1 U968 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n870), .Z(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n873) );
  XOR2_X1 U973 ( .A(n871), .B(KEYINPUT46), .Z(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n885) );
  NAND2_X1 U975 ( .A1(G139), .A2(n886), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G103), .A2(n887), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G127), .A2(n894), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G115), .A2(n891), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n878), .Z(n879) );
  XNOR2_X1 U982 ( .A(KEYINPUT47), .B(n879), .ZN(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n882), .Z(n945) );
  XOR2_X1 U985 ( .A(G164), .B(n945), .Z(n883) );
  XNOR2_X1 U986 ( .A(G162), .B(n883), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n903) );
  NAND2_X1 U988 ( .A1(G142), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G106), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(KEYINPUT45), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G130), .A2(n894), .ZN(n895) );
  XNOR2_X1 U995 ( .A(KEYINPUT111), .B(n895), .ZN(n896) );
  NOR2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n898), .B(n935), .Z(n901) );
  XNOR2_X1 U998 ( .A(G160), .B(n899), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1001 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(G171), .B(n996), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n907), .B(G286), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2427), .ZN(n920) );
  XOR2_X1 U1008 ( .A(G2430), .B(KEYINPUT106), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G2443), .B(G2451), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1011 ( .A(G2446), .B(KEYINPUT105), .Z(n914) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G1348), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(n916), .B(n915), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2435), .B(G2438), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(n927), .ZN(G401) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n941) );
  XOR2_X1 U1032 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1035 ( .A(KEYINPUT115), .B(n937), .Z(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT116), .B(n944), .ZN(n950) );
  XOR2_X1 U1040 ( .A(G2072), .B(n945), .Z(n947) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT50), .B(n948), .Z(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n976), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n953), .A2(G29), .ZN(n1047) );
  XNOR2_X1 U1049 ( .A(G2090), .B(G35), .ZN(n971) );
  XNOR2_X1 U1050 ( .A(n954), .B(G32), .ZN(n958) );
  XOR2_X1 U1051 ( .A(n955), .B(KEYINPUT117), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G27), .B(n956), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT118), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G25), .B(n960), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G26), .B(n961), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(n962), .A2(G28), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1068 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n979), .ZN(n1045) );
  XNOR2_X1 U1071 ( .A(G16), .B(KEYINPUT56), .ZN(n1011) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n982), .B(KEYINPUT57), .ZN(n1009) );
  XNOR2_X1 U1075 ( .A(n983), .B(G1341), .ZN(n1007) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G303), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n995) );
  XNOR2_X1 U1078 ( .A(n986), .B(G1956), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(KEYINPUT119), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(KEYINPUT120), .A2(n988), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n988), .A2(KEYINPUT120), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n998), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(n996), .B(G1348), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(n1030), .B(G171), .ZN(n1000) );
  INV_X1 U1088 ( .A(KEYINPUT120), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(KEYINPUT121), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1043) );
  INV_X1 U1097 ( .A(G16), .ZN(n1041) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1014) );
  XNOR2_X1 U1099 ( .A(n1012), .B(G22), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G24), .B(G1986), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1017), .Z(n1038) );
  XOR2_X1 U1104 ( .A(G1341), .B(G19), .Z(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT123), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G6), .B(G1981), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT124), .B(n1021), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(G4), .B(KEYINPUT125), .Z(n1023) );
  XNOR2_X1 U1110 ( .A(G1348), .B(KEYINPUT59), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(n1023), .B(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT122), .B(G1956), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(G20), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(KEYINPUT60), .B(n1029), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(n1030), .B(G5), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1035) );
  XNOR2_X1 U1119 ( .A(KEYINPUT126), .B(G1966), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(G21), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1122 ( .A(KEYINPUT127), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XNOR2_X1 U1124 ( .A(KEYINPUT61), .B(n1039), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1126 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U1127 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1128 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1048), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

