//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  XOR2_X1   g000(.A(KEYINPUT75), .B(G902), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT79), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT68), .B(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT76), .B1(new_n190), .B2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT68), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n195), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n197), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G110), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n196), .B1(new_n192), .B2(G128), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT24), .B(G110), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G125), .B(G140), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT16), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n214), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(G146), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT78), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n218), .A3(new_n215), .A4(G146), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n209), .A2(new_n212), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n202), .A2(new_n204), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n202), .A2(KEYINPUT77), .A3(new_n204), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n223), .A2(G110), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n215), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n216), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n206), .A2(new_n207), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n189), .B(new_n220), .C1(new_n225), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n203), .B1(new_n221), .B2(new_n222), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n232), .B2(new_n224), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n212), .A3(new_n219), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n205), .B2(new_n208), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G137), .ZN(new_n237));
  INV_X1    g051(.A(G953), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n238), .A2(G221), .A3(G234), .ZN(new_n239));
  XOR2_X1   g053(.A(new_n237), .B(new_n239), .Z(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(KEYINPUT79), .B(new_n240), .C1(new_n233), .C2(new_n235), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n188), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT80), .B(KEYINPUT25), .Z(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n187), .B2(G234), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n244), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n250), .A2(G902), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT81), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n242), .A2(new_n243), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n248), .A2(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT32), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  INV_X1    g073(.A(G210), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n260), .A2(G237), .A3(G953), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n268), .A2(new_n270), .A3(new_n275), .A4(new_n271), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  OR2_X1    g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  INV_X1    g093(.A(G143), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G146), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n211), .A2(G143), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n278), .B(new_n279), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT65), .B1(new_n280), .B2(G146), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT65), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n211), .A3(G143), .ZN(new_n286));
  INV_X1    g100(.A(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(G146), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n272), .A2(KEYINPUT66), .A3(G131), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n277), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT1), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n293), .B1(G143), .B2(new_n211), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n294), .A2(new_n200), .B1(new_n281), .B2(new_n282), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n284), .A2(new_n286), .A3(new_n288), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n271), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n267), .A2(G137), .ZN(new_n300));
  OAI21_X1  g114(.A(G131), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT69), .ZN(new_n303));
  OR2_X1    g117(.A1(KEYINPUT2), .A2(G113), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n193), .A2(new_n195), .A3(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT2), .A2(G113), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT67), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT2), .A3(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n304), .A2(new_n305), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n305), .A2(new_n312), .B1(new_n310), .B2(new_n304), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n303), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n305), .A2(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n304), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n305), .A2(new_n310), .A3(new_n304), .A4(new_n312), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(KEYINPUT69), .A3(new_n319), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n292), .A2(new_n302), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n265), .B1(new_n321), .B2(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n292), .A2(new_n302), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n292), .A2(new_n315), .A3(new_n320), .A4(new_n302), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(KEYINPUT74), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n292), .A2(new_n332), .A3(new_n302), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n265), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n264), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n292), .A2(KEYINPUT30), .A3(new_n302), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n292), .A2(new_n340), .A3(KEYINPUT30), .A4(new_n302), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XOR2_X1   g156(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n323), .A2(new_n344), .B1(new_n315), .B2(new_n320), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n327), .A2(new_n264), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n337), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n350));
  AOI211_X1 g164(.A(new_n350), .B(new_n347), .C1(new_n342), .C2(new_n345), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n336), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G472), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n258), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n329), .A2(new_n335), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n324), .B1(KEYINPUT74), .B2(new_n323), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT28), .B1(new_n358), .B2(new_n333), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n265), .B1(new_n325), .B2(new_n327), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT29), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n357), .A2(new_n361), .A3(new_n264), .ZN(new_n362));
  INV_X1    g176(.A(new_n264), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n346), .A2(new_n363), .A3(new_n327), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n187), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n365));
  OAI21_X1  g179(.A(G472), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n329), .A2(new_n335), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n363), .ZN(new_n368));
  INV_X1    g182(.A(new_n351), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n342), .A2(new_n345), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT31), .B1(new_n370), .B2(new_n347), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  INV_X1    g195(.A(G227), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G953), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n381), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  AND4_X1   g200(.A1(new_n284), .A2(new_n286), .A3(new_n288), .A4(new_n296), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n281), .B2(new_n293), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT82), .B(KEYINPUT1), .C1(new_n280), .C2(G146), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(G128), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n284), .A2(new_n286), .A3(new_n288), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n394), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n394), .A2(G107), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(G104), .ZN(new_n403));
  OAI21_X1  g217(.A(G101), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n386), .B1(new_n393), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G101), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n410), .A3(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n290), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n405), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT10), .A3(new_n298), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n277), .A2(new_n291), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n406), .A2(new_n416), .A3(new_n412), .A4(new_n414), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n385), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n413), .A2(new_n298), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n390), .A2(G128), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n211), .A2(G143), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT82), .B1(new_n424), .B2(KEYINPUT1), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n392), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n405), .B1(new_n426), .B2(new_n297), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT12), .B1(new_n428), .B2(new_n416), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT12), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n417), .B(new_n430), .C1(new_n427), .C2(new_n422), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n429), .A2(new_n419), .A3(new_n385), .A4(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n188), .B1(new_n421), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n380), .B1(new_n433), .B2(new_n378), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n418), .A2(new_n419), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n384), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(new_n419), .A3(new_n431), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n385), .B1(new_n437), .B2(KEYINPUT83), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n429), .A2(new_n419), .A3(new_n439), .A4(new_n431), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n436), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G469), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n377), .B1(new_n434), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n257), .A2(new_n374), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  NOR2_X1   g259(.A1(G237), .A2(G953), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(G143), .A3(G214), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(G143), .B1(new_n446), .B2(G214), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT17), .B(G131), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n227), .A2(new_n216), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  INV_X1    g267(.A(new_n449), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n275), .A3(new_n447), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n452), .B1(new_n456), .B2(KEYINPUT17), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT17), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(KEYINPUT91), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G113), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(new_n394), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n210), .B(new_n211), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT18), .B(G131), .C1(new_n448), .C2(new_n449), .ZN(new_n464));
  NAND2_X1  g278(.A1(KEYINPUT18), .A2(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n454), .A2(new_n447), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n456), .A2(new_n217), .A3(new_n219), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n210), .A2(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n211), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT90), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n210), .B(KEYINPUT19), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(new_n211), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n462), .B1(new_n478), .B2(new_n467), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n445), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT20), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n460), .A2(new_n462), .A3(new_n467), .ZN(new_n482));
  INV_X1    g296(.A(new_n467), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n469), .B2(new_n477), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n462), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT20), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n445), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n462), .B1(new_n460), .B2(new_n467), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n379), .B1(new_n468), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G475), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n375), .A2(new_n249), .A3(G953), .ZN(new_n493));
  INV_X1    g307(.A(G122), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(new_n494), .B2(G116), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT93), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n494), .A2(G116), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(KEYINPUT94), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(G116), .B2(new_n494), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n494), .A2(KEYINPUT14), .A3(G116), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G107), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n280), .A2(G128), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n200), .A2(G143), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G134), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n267), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n311), .A2(G122), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n497), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n508), .A2(new_n509), .B1(new_n511), .B2(new_n397), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n504), .A2(KEYINPUT95), .A3(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n397), .ZN(new_n518));
  OAI21_X1  g332(.A(G107), .B1(new_n497), .B2(new_n510), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT13), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(G134), .C1(KEYINPUT13), .C2(new_n505), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n509), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n509), .A2(new_n523), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n520), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n493), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n493), .ZN(new_n528));
  INV_X1    g342(.A(new_n526), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n528), .B(new_n529), .C1(new_n515), .C2(new_n516), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n187), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G478), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n531), .B(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n238), .A2(G952), .ZN(new_n539));
  INV_X1    g353(.A(G234), .ZN(new_n540));
  INV_X1    g354(.A(G237), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n238), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT21), .B(G898), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n492), .A2(new_n538), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n283), .A2(new_n289), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G125), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT84), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(KEYINPUT84), .A3(G125), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT85), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT85), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT84), .B1(new_n548), .B2(G125), .ZN(new_n555));
  AOI211_X1 g369(.A(new_n550), .B(new_n214), .C1(new_n283), .C2(new_n289), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n295), .A2(new_n214), .A3(new_n297), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n553), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G224), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(G953), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n561), .A2(KEYINPUT88), .A3(KEYINPUT7), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT88), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n553), .A2(new_n557), .A3(new_n564), .A4(new_n560), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n551), .A3(new_n552), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n563), .B1(KEYINPUT87), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(KEYINPUT87), .B2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G110), .B(G122), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT8), .Z(new_n575));
  INV_X1    g389(.A(KEYINPUT5), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n190), .A2(new_n576), .A3(G116), .ZN(new_n577));
  OAI211_X1 g391(.A(G113), .B(new_n577), .C1(new_n316), .C2(new_n576), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n319), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n405), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n319), .A3(new_n413), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n409), .A2(new_n411), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n324), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n585), .B2(new_n574), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n565), .A2(new_n569), .A3(new_n573), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n553), .A2(new_n557), .A3(new_n560), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n563), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n567), .ZN(new_n590));
  INV_X1    g404(.A(new_n574), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n409), .A2(new_n411), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n315), .B2(new_n320), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(new_n583), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n313), .A2(new_n314), .A3(new_n303), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT69), .B1(new_n318), .B2(new_n319), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n584), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n581), .A3(new_n574), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT6), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT6), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n591), .C1(new_n593), .C2(new_n583), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n587), .A2(new_n379), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G210), .B1(G237), .B2(G902), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT89), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n587), .A2(new_n602), .A3(new_n379), .A4(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n608), .A2(new_n607), .ZN(new_n610));
  OAI21_X1  g424(.A(G214), .B1(G237), .B2(G902), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n547), .A2(new_n609), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n444), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT97), .B(G101), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  NAND2_X1  g429(.A1(new_n606), .A2(new_n608), .ZN(new_n616));
  AOI21_X1  g430(.A(KEYINPUT98), .B1(new_n616), .B2(new_n611), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n618));
  INV_X1    g432(.A(new_n611), .ZN(new_n619));
  AOI211_X1 g433(.A(new_n618), .B(new_n619), .C1(new_n606), .C2(new_n608), .ZN(new_n620));
  INV_X1    g434(.A(new_n527), .ZN(new_n621));
  INV_X1    g435(.A(new_n530), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT33), .B1(new_n527), .B2(new_n530), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n188), .A2(new_n532), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n626), .A2(new_n627), .B1(new_n532), .B2(new_n531), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n481), .A2(new_n487), .B1(G475), .B2(new_n490), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n617), .A2(new_n620), .A3(new_n631), .A4(new_n546), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n328), .A2(new_n322), .B1(new_n334), .B2(new_n265), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n347), .B1(new_n342), .B2(new_n345), .ZN(new_n634));
  OAI22_X1  g448(.A1(new_n633), .A2(new_n264), .B1(new_n337), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n187), .B1(new_n635), .B2(new_n351), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n636), .A2(G472), .B1(new_n353), .B2(new_n372), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n257), .A2(new_n443), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  NOR2_X1   g455(.A1(new_n617), .A2(new_n620), .ZN(new_n642));
  INV_X1    g456(.A(new_n546), .ZN(new_n643));
  INV_X1    g457(.A(new_n537), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n531), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n492), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n638), .A2(new_n637), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  OR2_X1    g465(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n652));
  OR3_X1    g466(.A1(new_n233), .A2(new_n235), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n233), .B2(new_n235), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n255), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n256), .A2(new_n252), .A3(new_n187), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n250), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n657), .B1(new_n659), .B2(new_n247), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n637), .A3(new_n443), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n612), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT37), .B(G110), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT100), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n616), .A2(new_n611), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n618), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n611), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n538), .A2(new_n629), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n543), .B1(new_n544), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n668), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n374), .A2(new_n443), .A3(new_n660), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n666), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n672), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n646), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n617), .A2(new_n620), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n374), .A2(new_n443), .A3(new_n660), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(KEYINPUT101), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT102), .B(G128), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G30));
  NAND2_X1  g498(.A1(new_n609), .A2(new_n610), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n645), .A2(new_n629), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n672), .B(KEYINPUT39), .Z(new_n690));
  NAND2_X1  g504(.A1(new_n443), .A2(new_n690), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n619), .B(new_n689), .C1(new_n691), .C2(KEYINPUT40), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n363), .B1(new_n346), .B2(new_n327), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n325), .A2(new_n327), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n379), .B1(new_n694), .B2(new_n264), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n355), .A2(new_n373), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n655), .B(KEYINPUT99), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n248), .B2(new_n253), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n687), .A2(new_n692), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR3_X1   g517(.A1(new_n628), .A2(new_n629), .A3(new_n672), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n680), .A2(new_n642), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  OAI21_X1  g520(.A(new_n433), .B1(KEYINPUT104), .B2(new_n378), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n378), .A2(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(new_n432), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n420), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n708), .B1(new_n710), .B2(new_n188), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n377), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n257), .A2(new_n374), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n642), .A3(new_n643), .A4(new_n630), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT105), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n715), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n714), .A2(new_n642), .A3(new_n643), .A4(new_n646), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  INV_X1    g534(.A(new_n712), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n376), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n617), .A3(new_n620), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n374), .A2(new_n547), .A3(new_n660), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT106), .B(G119), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G21));
  NOR3_X1   g541(.A1(new_n617), .A2(new_n620), .A3(new_n689), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n712), .A2(new_n546), .A3(new_n377), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n694), .A2(KEYINPUT28), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n264), .B1(new_n335), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n730), .B1(new_n349), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n363), .B1(new_n359), .B2(new_n360), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n734), .B(KEYINPUT108), .C1(new_n337), .C2(new_n634), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n735), .A3(new_n369), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n353), .B(KEYINPUT107), .Z(new_n737));
  AOI22_X1  g551(.A1(new_n736), .A2(new_n737), .B1(new_n636), .B2(G472), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n729), .A2(new_n257), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n728), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  AND3_X1   g555(.A1(new_n738), .A2(new_n660), .A3(new_n704), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n642), .A3(new_n713), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n258), .C1(new_n352), .C2(new_n354), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n373), .A3(new_n366), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n372), .A2(new_n353), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n745), .B1(new_n748), .B2(new_n258), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n257), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n437), .A2(KEYINPUT83), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n384), .A3(new_n440), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT109), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n441), .C2(KEYINPUT109), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n377), .B1(new_n754), .B2(new_n434), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n685), .A2(new_n611), .A3(new_n755), .A4(new_n704), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT42), .B1(new_n750), .B2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n685), .A2(new_n611), .A3(new_n755), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n257), .A2(new_n374), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n630), .A2(new_n677), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n275), .ZN(G33));
  AOI21_X1  g578(.A(new_n619), .B1(new_n609), .B2(new_n610), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n257), .A3(new_n374), .A4(new_n755), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n678), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT111), .B(G134), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G36));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n628), .A2(new_n492), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT114), .A3(KEYINPUT43), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n628), .B2(new_n492), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT113), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT115), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n699), .A2(new_n637), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT115), .B1(new_n776), .B2(new_n779), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n770), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n776), .A2(new_n779), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n780), .A4(new_n781), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n433), .A2(new_n378), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n752), .B1(new_n435), .B2(new_n384), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n378), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n753), .B1(new_n441), .B2(KEYINPUT109), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n380), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n789), .B1(new_n796), .B2(KEYINPUT46), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n795), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n376), .B(new_n690), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n784), .A2(new_n765), .A3(new_n788), .A4(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(KEYINPUT116), .B(G137), .Z(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(G39));
  OAI21_X1  g617(.A(new_n376), .B1(new_n797), .B2(new_n798), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(KEYINPUT47), .B(new_n376), .C1(new_n797), .C2(new_n798), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n765), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n257), .A3(new_n374), .A4(new_n760), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  INV_X1    g626(.A(new_n687), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n257), .A2(new_n355), .A3(new_n373), .A4(new_n696), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n712), .A2(KEYINPUT49), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n771), .A3(new_n611), .A4(new_n376), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n721), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n674), .A2(new_n666), .A3(new_n675), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT101), .B1(new_n679), .B2(new_n680), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n755), .A2(new_n677), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n700), .A2(new_n642), .A3(new_n688), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n705), .A3(new_n743), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT52), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n758), .B2(new_n742), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n765), .A2(new_n755), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n738), .A2(new_n660), .A3(new_n704), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n830), .A3(KEYINPUT117), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n492), .A2(new_n538), .A3(new_n672), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n765), .A2(new_n833), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n766), .A2(new_n678), .B1(new_n834), .B2(new_n675), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n832), .A2(new_n763), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n612), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n257), .A2(new_n374), .A3(new_n443), .ZN(new_n838));
  INV_X1    g652(.A(new_n661), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n715), .A2(new_n840), .A3(new_n719), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n546), .B1(new_n631), .B2(new_n670), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n685), .A2(new_n619), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n638), .A2(new_n842), .A3(new_n843), .A4(new_n637), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n725), .A2(new_n740), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n699), .A2(new_n697), .A3(new_n677), .A4(new_n755), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n617), .A2(new_n760), .A3(new_n620), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n728), .A2(new_n847), .B1(new_n848), .B2(new_n680), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n682), .A2(new_n849), .A3(new_n850), .A4(new_n743), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n826), .A2(new_n836), .A3(new_n846), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n612), .B1(new_n444), .B2(new_n661), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n632), .B2(new_n714), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n723), .A2(new_n724), .B1(new_n728), .B2(new_n739), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n719), .A3(new_n857), .A4(new_n844), .ZN(new_n858));
  INV_X1    g672(.A(new_n835), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n758), .A2(new_n742), .A3(new_n827), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT117), .B1(new_n829), .B2(new_n830), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n859), .A2(new_n862), .A3(new_n757), .A4(new_n762), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n824), .A2(new_n705), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n853), .B1(new_n865), .B2(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n864), .A2(new_n826), .A3(new_n866), .A4(new_n851), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n854), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT119), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n854), .A2(new_n867), .A3(new_n868), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n865), .B2(KEYINPUT52), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n854), .B1(new_n852), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n809), .A2(new_n542), .A3(new_n722), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n629), .A3(new_n628), .A4(new_n814), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n785), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n738), .A2(new_n660), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n687), .A2(new_n611), .A3(new_n722), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n257), .A2(new_n738), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n785), .A2(new_n543), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(KEYINPUT50), .A3(new_n885), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n883), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n712), .A2(new_n376), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n765), .B(new_n890), .C1(new_n808), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n878), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n881), .A2(new_n750), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT48), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n630), .A3(new_n814), .ZN(new_n900));
  INV_X1    g714(.A(new_n723), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n539), .B(new_n900), .C1(new_n888), .C2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n899), .B(new_n903), .C1(new_n895), .C2(new_n896), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n877), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n819), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NAND2_X1  g721(.A1(new_n599), .A2(new_n601), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(new_n590), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n187), .B1(new_n854), .B2(new_n867), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n605), .ZN(new_n912));
  OR2_X1    g726(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n238), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n912), .A2(new_n910), .A3(new_n913), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(G51));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n187), .B(new_n794), .C1(new_n854), .C2(new_n867), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n380), .B(KEYINPUT57), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n868), .B1(new_n854), .B2(new_n867), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n869), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n710), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  INV_X1    g741(.A(new_n868), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n825), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n824), .A2(new_n705), .A3(new_n743), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n850), .B1(new_n930), .B2(new_n682), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n932), .B2(new_n864), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n826), .A2(new_n851), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n715), .A2(new_n840), .A3(new_n719), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n835), .B1(new_n861), .B2(new_n860), .ZN(new_n936));
  INV_X1    g750(.A(new_n845), .ZN(new_n937));
  INV_X1    g751(.A(new_n763), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n866), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n928), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n871), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n710), .B1(new_n943), .B2(new_n922), .ZN(new_n944));
  OAI211_X1 g758(.A(KEYINPUT122), .B(new_n916), .C1(new_n944), .C2(new_n921), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n927), .A2(new_n945), .ZN(G54));
  AND2_X1   g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n911), .A2(new_n485), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n485), .B1(new_n911), .B2(new_n947), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(new_n915), .ZN(G60));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT59), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n626), .B1(new_n877), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n626), .A3(new_n953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n916), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(new_n854), .A2(new_n867), .ZN(new_n958));
  NAND2_X1  g772(.A1(G217), .A2(G902), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT123), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n256), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n915), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT124), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT61), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n958), .A2(new_n653), .A3(new_n654), .A4(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n963), .B(new_n966), .C1(new_n964), .C2(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(G66));
  OAI21_X1  g784(.A(G953), .B1(new_n545), .B2(new_n562), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n846), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n908), .B1(G898), .B2(new_n238), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  NAND2_X1  g788(.A1(new_n801), .A2(new_n811), .ZN(new_n975));
  INV_X1    g789(.A(new_n759), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n630), .A2(new_n646), .ZN(new_n977));
  NOR4_X1   g791(.A1(new_n976), .A2(new_n691), .A3(new_n809), .A4(new_n977), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n682), .A2(new_n705), .A3(new_n743), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n702), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n983), .A3(new_n702), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n238), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n323), .A2(new_n344), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n342), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(new_n474), .ZN(new_n989));
  INV_X1    g803(.A(new_n728), .ZN(new_n990));
  OR3_X1    g804(.A1(new_n799), .A2(new_n990), .A3(new_n750), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n991), .A2(new_n980), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n763), .A2(new_n767), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n992), .A2(new_n801), .A3(new_n811), .A4(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n996));
  AOI22_X1  g810(.A1(new_n986), .A2(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n382), .B2(new_n671), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G72));
  NOR4_X1   g813(.A1(new_n985), .A2(new_n975), .A3(new_n858), .A4(new_n978), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT63), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n693), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n991), .A2(new_n980), .A3(new_n993), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n975), .A2(new_n1006), .A3(new_n858), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(new_n1003), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1003), .ZN(new_n1009));
  OAI211_X1 g823(.A(KEYINPUT126), .B(new_n1009), .C1(new_n994), .C2(new_n858), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n346), .A2(new_n363), .A3(new_n327), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1011), .A2(new_n693), .A3(new_n1002), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n915), .B1(new_n875), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1004), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(KEYINPUT127), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT127), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1004), .A2(new_n1012), .A3(new_n1017), .A4(new_n1014), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(G57));
endmodule


