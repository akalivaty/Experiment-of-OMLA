//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT34), .ZN(new_n204));
  OR2_X1    g003(.A1(G113gat), .A2(G120gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  NAND2_X1  g005(.A1(G113gat), .A2(G120gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G127gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT69), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n208), .B(new_n213), .C1(KEYINPUT69), .C2(new_n210), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n205), .A2(new_n215), .A3(new_n207), .ZN(new_n216));
  AND2_X1   g015(.A1(G113gat), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G113gat), .A2(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT70), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n206), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n225));
  AND3_X1   g024(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(KEYINPUT23), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(KEYINPUT24), .ZN(new_n236));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT64), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n237), .A2(KEYINPUT24), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(G183gat), .A3(G190gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n234), .A2(new_n240), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n243), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n247), .A2(new_n248), .B1(new_n234), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G190gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n235), .A2(KEYINPUT27), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT27), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G183gat), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT26), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n230), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n267), .B(new_n268), .C1(new_n227), .C2(new_n226), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n237), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n268), .ZN(new_n277));
  NOR3_X1   g076(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n276), .A2(new_n279), .B1(new_n261), .B2(KEYINPUT28), .ZN(new_n280));
  INV_X1    g079(.A(new_n237), .ZN(new_n281));
  AND4_X1   g080(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n260), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(new_n264), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n271), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n222), .B1(new_n253), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n231), .A2(new_n233), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n274), .A2(new_n275), .B1(KEYINPUT23), .B2(new_n230), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n288), .B(new_n289), .C1(new_n244), .C2(new_n245), .ZN(new_n290));
  INV_X1    g089(.A(new_n246), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n248), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n252), .A2(new_n234), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n214), .A2(new_n221), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n271), .A4(new_n285), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G227gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n204), .B1(new_n297), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(KEYINPUT34), .B(new_n300), .C1(new_n287), .C2(new_n296), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n300), .A3(new_n296), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT33), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(KEYINPUT32), .ZN(new_n308));
  XOR2_X1   g107(.A(G71gat), .B(G99gat), .Z(new_n309));
  XNOR2_X1  g108(.A(G15gat), .B(G43gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n307), .A2(new_n308), .A3(new_n314), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(KEYINPUT33), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n316), .ZN(new_n317));
  AND4_X1   g116(.A1(new_n304), .A2(new_n313), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n312), .B2(KEYINPUT71), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n304), .B1(new_n320), .B2(new_n315), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n203), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n323));
  INV_X1    g122(.A(new_n304), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n304), .A3(new_n315), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(KEYINPUT36), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G8gat), .B(G36gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G64gat), .ZN(new_n329));
  INV_X1    g128(.A(G92gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n270), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n332), .B(new_n334), .C1(new_n253), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(new_n292), .B2(new_n293), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n337), .B2(new_n333), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n271), .A2(new_n285), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n339), .B2(new_n294), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n336), .B(new_n338), .C1(new_n340), .C2(new_n334), .ZN(new_n341));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n343));
  INV_X1    g142(.A(G211gat), .ZN(new_n344));
  INV_X1    g143(.A(G218gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n342), .A3(new_n346), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n350), .A2(KEYINPUT72), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT72), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n341), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n351), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n358), .B(new_n333), .C1(new_n253), .C2(new_n335), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n294), .A2(new_n334), .A3(new_n271), .A4(new_n285), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n331), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n331), .ZN(new_n364));
  AOI211_X1 g163(.A(new_n364), .B(new_n361), .C1(new_n341), .C2(new_n354), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(KEYINPUT30), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT2), .ZN(new_n368));
  OR2_X1    g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n377));
  XNOR2_X1  g176(.A(G141gat), .B(G148gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT2), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(G155gat), .B2(G162gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n373), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n372), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n387), .A3(new_n295), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n222), .A2(new_n385), .A3(KEYINPUT4), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n376), .A2(new_n295), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n385), .B(new_n295), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(KEYINPUT5), .C1(new_n391), .C2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n392), .A2(KEYINPUT5), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT77), .B1(new_n376), .B2(new_n295), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n222), .A2(new_n385), .A3(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n398), .A2(new_n390), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n390), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n388), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(KEYINPUT76), .B(KEYINPUT0), .Z(new_n405));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G57gat), .B(G85gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n403), .A3(new_n409), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(KEYINPUT6), .A3(new_n410), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT74), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n361), .B1(new_n341), .B2(new_n354), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n331), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT74), .B(KEYINPUT30), .C1(new_n418), .C2(new_n331), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n366), .B(new_n416), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(G50gat), .ZN(new_n425));
  XOR2_X1   g224(.A(G78gat), .B(G106gat), .Z(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n350), .B2(new_n351), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n386), .B1(new_n428), .B2(KEYINPUT80), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n356), .A2(KEYINPUT80), .A3(new_n358), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n376), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n376), .A2(KEYINPUT3), .ZN(new_n432));
  OAI22_X1  g231(.A1(new_n432), .A2(KEYINPUT29), .B1(new_n352), .B2(new_n353), .ZN(new_n433));
  INV_X1    g232(.A(G228gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n299), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT79), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n347), .A2(new_n437), .A3(new_n349), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n358), .B(new_n438), .C1(new_n356), .C2(new_n437), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n385), .B1(new_n439), .B2(new_n386), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n356), .B1(new_n387), .B2(new_n358), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n440), .A2(new_n441), .B1(new_n434), .B2(new_n299), .ZN(new_n442));
  INV_X1    g241(.A(G22gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(KEYINPUT82), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n436), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n436), .B2(new_n442), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n427), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT83), .B(new_n427), .C1(new_n445), .C2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT81), .B1(new_n436), .B2(new_n442), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n427), .B1(new_n452), .B2(new_n443), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(new_n443), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n436), .A2(new_n442), .A3(KEYINPUT81), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n322), .A2(new_n327), .B1(new_n423), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n331), .B1(new_n418), .B2(KEYINPUT38), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n459), .A2(new_n414), .A3(new_n415), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT37), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n331), .B1(new_n418), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n359), .A2(new_n360), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n341), .A2(new_n354), .B1(new_n356), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT38), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n418), .A2(new_n461), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT37), .B(new_n361), .C1(new_n341), .C2(new_n354), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n355), .A2(new_n362), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n364), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n420), .B2(new_n419), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT74), .B1(new_n365), .B2(KEYINPUT30), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n419), .A2(new_n417), .A3(new_n420), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  INV_X1    g278(.A(new_n388), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n376), .A2(new_n295), .A3(KEYINPUT77), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n399), .B1(new_n222), .B2(new_n385), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT4), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n398), .A2(new_n400), .A3(new_n390), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT84), .B1(new_n485), .B2(new_n391), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n388), .B1(new_n401), .B2(new_n402), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(new_n392), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n395), .B2(new_n391), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n486), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n409), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT39), .B1(new_n486), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n479), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n486), .A2(new_n489), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n490), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n497), .A2(KEYINPUT40), .A3(new_n409), .A4(new_n492), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n411), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n471), .B(new_n472), .C1(new_n478), .C2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n458), .A2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n472), .A2(new_n326), .A3(new_n325), .ZN(new_n502));
  INV_X1    g301(.A(new_n423), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(KEYINPUT35), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n472), .A2(new_n326), .A3(new_n325), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n423), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n202), .B1(new_n501), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n458), .A2(new_n500), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n507), .A4(new_n504), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT87), .B(G29gat), .ZN(new_n512));
  INV_X1    g311(.A(G36gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT14), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  OR2_X1    g318(.A1(G43gat), .A2(G50gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n515), .A2(KEYINPUT14), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n515), .A2(KEYINPUT14), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(new_n528), .C1(new_n512), .C2(new_n513), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT15), .A3(new_n518), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(new_n523), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT88), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(G1gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G1gat), .B2(new_n536), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G8gat), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n541), .C1(G1gat), .C2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n532), .A3(KEYINPUT17), .A4(new_n530), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n533), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(G229gat), .A2(G233gat), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n546), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n533), .B(new_n543), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n548), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(KEYINPUT18), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n543), .B1(new_n533), .B2(new_n534), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n560), .A2(new_n545), .B1(new_n533), .B2(new_n543), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n548), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT89), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n554), .A2(new_n557), .A3(new_n559), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G169gat), .B(G197gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT86), .B(KEYINPUT11), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT18), .B1(new_n561), .B2(new_n548), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n553), .A2(new_n573), .A3(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G57gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(G64gat), .ZN(new_n577));
  INV_X1    g376(.A(G64gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(G57gat), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT9), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  OR2_X1    g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n578), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(G57gat), .B2(new_n578), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n577), .A2(KEYINPUT91), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT7), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n592), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n596), .A2(new_n598), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n603), .B2(new_n595), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n590), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n601), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n600), .A3(new_n595), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n607), .A2(new_n583), .A3(new_n589), .A4(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(new_n609), .B2(new_n606), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n602), .A2(new_n604), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n583), .A2(new_n589), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(KEYINPUT95), .A3(KEYINPUT10), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT96), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(G176gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n605), .A2(new_n609), .ZN(new_n626));
  INV_X1    g425(.A(new_n617), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n619), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n619), .A2(new_n628), .A3(KEYINPUT98), .A4(new_n621), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n625), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G127gat), .B(G155gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT21), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n590), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(G211gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n344), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n235), .B1(new_n544), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n544), .A2(new_n651), .A3(new_n235), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(new_n652), .A3(new_n649), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n646), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n649), .B1(new_n656), .B2(new_n652), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n653), .A2(new_n654), .A3(new_n650), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(new_n660), .A3(new_n644), .A4(new_n645), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G232gat), .A2(G233gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT92), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n666));
  XNOR2_X1  g465(.A(G190gat), .B(G218gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n613), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n535), .A2(new_n545), .A3(new_n669), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n533), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT93), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n670), .B2(new_n671), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n668), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  INV_X1    g478(.A(new_n668), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n675), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n637), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n509), .A2(new_n511), .A3(new_n575), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n416), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT99), .B(G1gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n684), .A2(new_n478), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n509), .A2(new_n511), .A3(new_n575), .ZN(new_n695));
  INV_X1    g494(.A(new_n478), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n683), .A4(new_n690), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(KEYINPUT100), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G8gat), .B1(new_n684), .B2(new_n478), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n694), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n694), .A2(new_n699), .A3(KEYINPUT101), .A4(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1325gat));
  NAND2_X1  g504(.A1(new_n322), .A2(new_n327), .ZN(new_n706));
  OAI21_X1  g505(.A(G15gat), .B1(new_n684), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n325), .A2(new_n326), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(G15gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n684), .B2(new_n709), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n685), .A2(new_n457), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n637), .A2(new_n662), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n680), .B1(new_n679), .B2(new_n675), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n676), .A2(new_n668), .A3(new_n677), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n509), .A2(new_n511), .A3(new_n575), .A4(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n512), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n416), .A3(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT45), .Z(new_n723));
  INV_X1    g522(.A(new_n718), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n509), .A2(KEYINPUT44), .A3(new_n511), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n510), .A2(new_n507), .A3(new_n504), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n553), .A2(new_n573), .A3(new_n571), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n565), .B2(new_n571), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n686), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n721), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n723), .B1(new_n737), .B2(new_n738), .ZN(G1328gat));
  NAND2_X1  g538(.A1(new_n696), .A2(new_n513), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n720), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n720), .B2(new_n740), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n730), .A2(new_n696), .A3(new_n733), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(new_n513), .ZN(G1329gat));
  INV_X1    g545(.A(new_n706), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n725), .A2(new_n729), .A3(new_n747), .A4(new_n733), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G43gat), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n708), .A2(G43gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n720), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n720), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(KEYINPUT104), .A3(new_n751), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n749), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n751), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT105), .B1(new_n749), .B2(new_n758), .ZN(new_n760));
  OAI22_X1  g559(.A1(KEYINPUT47), .A2(new_n756), .B1(new_n759), .B2(new_n760), .ZN(G1330gat));
  OR3_X1    g560(.A1(new_n720), .A2(G50gat), .A3(new_n472), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT48), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n725), .A2(new_n729), .A3(new_n457), .A4(new_n733), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n762), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n764), .B(new_n767), .ZN(G1331gat));
  AOI22_X1  g567(.A1(new_n631), .A2(new_n632), .B1(new_n625), .B2(new_n635), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n575), .A2(new_n682), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n726), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT107), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n416), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n576), .ZN(G1332gat));
  XOR2_X1   g573(.A(new_n771), .B(KEYINPUT107), .Z(new_n775));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n696), .B1(new_n776), .B2(new_n578), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT108), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT109), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n780), .A2(new_n776), .A3(new_n578), .A4(new_n782), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n775), .A2(new_n781), .A3(new_n778), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n775), .B2(new_n778), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n784), .A2(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(G1333gat));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788));
  OAI21_X1  g587(.A(G71gat), .B1(new_n772), .B2(new_n706), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n772), .A2(G71gat), .A3(new_n708), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(KEYINPUT50), .A3(new_n789), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n775), .A2(new_n457), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n575), .A2(new_n662), .A3(new_n769), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n730), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n416), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n416), .A2(new_n769), .A3(G85gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT111), .ZN(new_n802));
  INV_X1    g601(.A(new_n727), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n575), .A2(new_n662), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(KEYINPUT51), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n807));
  NOR4_X1   g606(.A1(new_n727), .A2(new_n575), .A3(new_n662), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n800), .A2(new_n809), .ZN(G1336gat));
  NOR2_X1   g609(.A1(new_n478), .A2(G92gat), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n637), .B(new_n811), .C1(new_n806), .C2(new_n808), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n725), .A2(new_n729), .A3(new_n696), .A4(new_n798), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G92gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n799), .B2(new_n706), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n708), .A2(G99gat), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n637), .B(new_n818), .C1(new_n806), .C2(new_n808), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n472), .A2(G106gat), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n637), .B(new_n821), .C1(new_n806), .C2(new_n808), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n725), .A2(new_n729), .A3(new_n457), .A4(new_n798), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g625(.A1(new_n683), .A2(new_n732), .ZN(new_n827));
  INV_X1    g626(.A(new_n662), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n561), .A2(new_n548), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n550), .A2(new_n551), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n570), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n574), .B(new_n831), .C1(new_n717), .C2(new_n716), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  INV_X1    g632(.A(new_n621), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n620), .B1(new_n616), .B2(new_n617), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n610), .A2(new_n612), .A3(new_n615), .A4(new_n627), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n625), .B1(new_n618), .B2(KEYINPUT54), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n619), .A2(KEYINPUT54), .A3(new_n621), .A4(new_n836), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n618), .A2(KEYINPUT54), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n625), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n633), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n832), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n574), .A2(new_n831), .ZN(new_n846));
  OAI22_X1  g645(.A1(new_n732), .A2(new_n844), .B1(new_n769), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n847), .B2(new_n718), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n828), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT112), .B(new_n845), .C1(new_n847), .C2(new_n718), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n827), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n696), .A2(new_n416), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n502), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n575), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n575), .A2(G113gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1340gat));
  AOI21_X1  g660(.A(G120gat), .B1(new_n855), .B2(new_n637), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n637), .A2(G120gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n859), .B2(new_n863), .ZN(G1341gat));
  AOI21_X1  g663(.A(new_n209), .B1(new_n859), .B2(new_n662), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n852), .A2(new_n502), .A3(new_n662), .A4(new_n853), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n869));
  AOI21_X1  g668(.A(G127gat), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT115), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n869), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n209), .B1(new_n872), .B2(new_n867), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n828), .B1(new_n857), .B2(new_n858), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n209), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n871), .A2(new_n876), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n855), .A2(new_n724), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n718), .B1(new_n857), .B2(new_n858), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n211), .B2(new_n882), .ZN(G1343gat));
  AND2_X1   g682(.A1(new_n853), .A2(new_n706), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n852), .B2(new_n457), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n472), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n847), .A2(new_n718), .ZN(new_n889));
  INV_X1    g688(.A(new_n845), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n828), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n888), .B1(new_n892), .B2(new_n827), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n575), .B(new_n884), .C1(new_n885), .C2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n747), .A2(new_n472), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n852), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n732), .A2(G141gat), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n853), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT58), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT58), .B1(new_n894), .B2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT117), .B1(new_n897), .B2(new_n416), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n852), .A2(new_n905), .A3(new_n686), .A4(new_n896), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n904), .A2(new_n478), .A3(new_n899), .A4(new_n906), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n902), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n903), .B1(new_n902), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(G1344gat));
  AND3_X1   g709(.A1(new_n904), .A2(new_n478), .A3(new_n906), .ZN(new_n911));
  INV_X1    g710(.A(G148gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n637), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n769), .A2(new_n662), .A3(new_n718), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n575), .A2(new_n915), .A3(KEYINPUT121), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n683), .B2(new_n732), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n662), .B2(new_n848), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n472), .B1(new_n920), .B2(KEYINPUT122), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n892), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n848), .A2(new_n849), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n828), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n888), .B1(new_n927), .B2(new_n827), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n637), .B(new_n884), .C1(new_n924), .C2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n912), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n928), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n921), .A2(new_n923), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(KEYINPUT57), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n934), .A2(KEYINPUT123), .A3(new_n637), .A4(new_n884), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n914), .B1(new_n931), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n637), .B(new_n884), .C1(new_n885), .C2(new_n893), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n912), .A2(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n913), .B1(new_n936), .B2(new_n943), .ZN(G1345gat));
  INV_X1    g743(.A(G155gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n911), .A2(new_n945), .A3(new_n662), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n884), .B1(new_n885), .B2(new_n893), .ZN(new_n947));
  OAI21_X1  g746(.A(G155gat), .B1(new_n947), .B2(new_n828), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1346gat));
  INV_X1    g748(.A(G162gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n911), .A2(new_n950), .A3(new_n724), .ZN(new_n951));
  OAI21_X1  g750(.A(G162gat), .B1(new_n947), .B2(new_n718), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1347gat));
  AOI21_X1  g752(.A(new_n506), .B1(new_n927), .B2(new_n827), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n478), .A2(new_n686), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(new_n223), .A3(new_n732), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n956), .B(KEYINPUT124), .Z(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n575), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n959), .B2(new_n223), .ZN(G1348gat));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n224), .A3(new_n637), .ZN(new_n961));
  OAI21_X1  g760(.A(G176gat), .B1(new_n956), .B2(new_n769), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1349gat));
  OAI21_X1  g762(.A(new_n235), .B1(new_n956), .B2(new_n828), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n954), .A2(new_n662), .A3(new_n955), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n263), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT60), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n249), .A3(new_n724), .ZN(new_n969));
  OAI21_X1  g768(.A(G190gat), .B1(new_n956), .B2(new_n718), .ZN(new_n970));
  NOR2_X1   g769(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n969), .A2(new_n972), .A3(new_n974), .ZN(G1351gat));
  INV_X1    g774(.A(G197gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n898), .A2(new_n955), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n732), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n706), .A2(new_n955), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n934), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n575), .A2(G197gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(KEYINPUT126), .B(new_n978), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1352gat));
  NOR3_X1   g786(.A1(new_n977), .A2(G204gat), .A3(new_n769), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT62), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n934), .A2(new_n637), .A3(new_n980), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G204gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n989), .A2(new_n991), .ZN(G1353gat));
  NOR3_X1   g791(.A1(new_n897), .A2(new_n686), .A3(new_n478), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n993), .A2(new_n344), .A3(new_n662), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n934), .A2(new_n662), .A3(new_n980), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  NOR3_X1   g797(.A1(new_n981), .A2(new_n345), .A3(new_n718), .ZN(new_n999));
  AOI21_X1  g798(.A(G218gat), .B1(new_n993), .B2(new_n724), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(G1355gat));
endmodule


