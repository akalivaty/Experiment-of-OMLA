//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1066, new_n1067;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT86), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT41), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT87), .Z(new_n207));
  XNOR2_X1  g006(.A(G134gat), .B(G162gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  INV_X1    g009(.A(G85gat), .ZN(new_n211));
  INV_X1    g010(.A(G92gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT7), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G85gat), .A3(G92gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G99gat), .B(G106gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(KEYINPUT8), .A2(new_n218), .B1(new_n211), .B2(new_n212), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n217), .B1(new_n216), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n219), .ZN(new_n223));
  INV_X1    g022(.A(new_n217), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(KEYINPUT88), .A3(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G43gat), .ZN(new_n230));
  INV_X1    g029(.A(G43gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G50gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT15), .ZN(new_n233));
  INV_X1    g032(.A(G29gat), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT14), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT14), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n230), .A2(new_n232), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT79), .A2(KEYINPUT15), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT79), .A2(KEYINPUT15), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n234), .A2(KEYINPUT78), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G29gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n241), .A2(new_n244), .B1(new_n248), .B2(G36gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n240), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G43gat), .B(G50gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT79), .B(KEYINPUT15), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT78), .B(G29gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n235), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT15), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n238), .A3(new_n236), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT80), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n239), .A2(KEYINPUT77), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n238), .A3(new_n260), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n259), .B(new_n261), .C1(new_n235), .C2(new_n254), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n251), .A2(new_n258), .B1(new_n262), .B2(new_n233), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n228), .A2(new_n263), .B1(new_n205), .B2(new_n204), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT81), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n233), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT17), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n263), .A2(KEYINPUT81), .A3(KEYINPUT17), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n268), .A2(KEYINPUT17), .A3(new_n269), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n228), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n265), .B(new_n266), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n266), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT81), .B1(new_n263), .B2(KEYINPUT17), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n267), .A3(new_n271), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n281), .B2(new_n264), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n209), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT90), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n282), .A3(new_n209), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n202), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n283), .B(KEYINPUT90), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n286), .B(KEYINPUT89), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT91), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G71gat), .A2(G78gat), .ZN(new_n294));
  OR2_X1    g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT9), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n294), .B(new_n295), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n294), .ZN(new_n299));
  INV_X1    g098(.A(G57gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G64gat), .ZN(new_n301));
  INV_X1    g100(.A(G64gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G57gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n294), .A2(new_n297), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(KEYINPUT85), .A3(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT21), .ZN(new_n312));
  NAND2_X1  g111(.A1(G231gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n312), .B(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G127gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(G15gat), .B(G22gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(G1gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT16), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(G1gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n317), .B1(new_n319), .B2(new_n316), .ZN(new_n320));
  INV_X1    g119(.A(G8gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(KEYINPUT21), .B2(new_n311), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n315), .A2(new_n323), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n326));
  INV_X1    g125(.A(G155gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G183gat), .B(G211gat), .Z(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n324), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n324), .B2(new_n325), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n336), .B1(new_n309), .B2(new_n310), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n222), .A2(new_n227), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n225), .A2(new_n226), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n298), .A2(KEYINPUT85), .A3(new_n306), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT85), .B1(new_n298), .B2(new_n306), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n307), .A2(new_n225), .A3(new_n226), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT10), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n335), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(new_n338), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n307), .A2(new_n225), .A3(new_n226), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n311), .B2(new_n340), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT92), .B(new_n347), .C1(new_n349), .C2(KEYINPUT10), .ZN(new_n350));
  NAND2_X1  g149(.A1(G230gat), .A2(G233gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT93), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n352), .ZN(new_n355));
  XNOR2_X1  g154(.A(G120gat), .B(G148gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(G176gat), .B(G204gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND3_X1  g157(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n353), .B1(new_n339), .B2(new_n345), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(new_n358), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n293), .A2(new_n334), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G113gat), .ZN(new_n369));
  INV_X1    g168(.A(G113gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G120gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT1), .ZN(new_n373));
  INV_X1    g172(.A(G134gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G127gat), .ZN(new_n375));
  INV_X1    g174(.A(G127gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G134gat), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n373), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n377), .ZN(new_n379));
  XNOR2_X1  g178(.A(G113gat), .B(G120gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n379), .B1(new_n380), .B2(KEYINPUT1), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n383));
  AND2_X1   g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  INV_X1    g183(.A(G169gat), .ZN(new_n385));
  INV_X1    g184(.A(G176gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G183gat), .A2(G190gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G183gat), .ZN(new_n393));
  INV_X1    g192(.A(G190gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT23), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n395), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n390), .A2(KEYINPUT65), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT65), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(G183gat), .A3(G190gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n403), .A3(new_n391), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n388), .B1(G169gat), .B2(G176gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407));
  AND4_X1   g206(.A1(KEYINPUT25), .A2(new_n398), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n383), .A2(new_n399), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT26), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT26), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(G169gat), .A2(G176gat), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n390), .B(new_n410), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n393), .A2(KEYINPUT27), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G183gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n417), .A3(new_n394), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT28), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT27), .B(G183gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT28), .A3(new_n394), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n414), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n382), .B1(new_n409), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT64), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n408), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n398), .A2(new_n406), .A3(new_n407), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n383), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n378), .A2(new_n381), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n412), .A2(new_n413), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n410), .A2(new_n390), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT28), .B1(new_n421), .B2(new_n394), .ZN(new_n437));
  AND4_X1   g236(.A1(KEYINPUT28), .A2(new_n415), .A3(new_n417), .A4(new_n394), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n432), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n427), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT34), .B1(new_n426), .B2(KEYINPUT67), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n424), .A2(new_n427), .A3(new_n440), .A4(new_n442), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(G15gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n447), .B(KEYINPUT66), .ZN(new_n451));
  INV_X1    g250(.A(G15gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n231), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n453), .A3(G43gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n409), .A2(new_n382), .A3(new_n423), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n433), .B1(new_n432), .B2(new_n439), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n426), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n424), .A2(new_n440), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT33), .B1(new_n464), .B2(new_n426), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n445), .B(new_n444), .C1(new_n465), .C2(new_n457), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(KEYINPUT32), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n446), .A2(new_n462), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n446), .A2(new_n462), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G228gat), .ZN(new_n475));
  INV_X1    g274(.A(G233gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n478), .A2(G155gat), .A3(G162gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT74), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(G141gat), .A2(G148gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT2), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT75), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT2), .ZN(new_n489));
  NAND2_X1  g288(.A1(G141gat), .A2(G148gat), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n482), .B1(new_n481), .B2(KEYINPUT2), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n485), .A2(new_n490), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n484), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT29), .ZN(new_n495));
  NOR2_X1   g294(.A1(G197gat), .A2(G204gat), .ZN(new_n496));
  AND2_X1   g295(.A1(G197gat), .A2(G204gat), .ZN(new_n497));
  AND2_X1   g296(.A1(G211gat), .A2(G218gat), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(KEYINPUT22), .ZN(new_n499));
  NOR2_X1   g298(.A1(G211gat), .A2(G218gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT69), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G197gat), .ZN(new_n504));
  INV_X1    g303(.A(G204gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G197gat), .A2(G204gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT22), .ZN(new_n508));
  NAND2_X1  g307(.A1(G211gat), .A2(G218gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G211gat), .ZN(new_n511));
  INV_X1    g310(.A(G218gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT69), .A3(new_n509), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n495), .B1(new_n503), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n494), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n502), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n510), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n480), .A2(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n481), .A2(new_n483), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n491), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n482), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n485), .B(new_n490), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(new_n517), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n521), .B1(new_n528), .B2(new_n495), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n477), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G22gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n495), .ZN(new_n532));
  INV_X1    g331(.A(new_n521), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n498), .A2(new_n500), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n495), .B1(new_n510), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n509), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n499), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n517), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AND4_X1   g338(.A1(new_n485), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n478), .B1(G155gat), .B2(G162gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n522), .B1(new_n541), .B2(new_n480), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n527), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n477), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n531), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n531), .B1(new_n530), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n474), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G22gat), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT76), .A3(new_n546), .A4(new_n473), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G50gat), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n549), .B2(new_n552), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n469), .B(new_n472), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n543), .A2(KEYINPUT3), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n528), .A3(new_n382), .ZN(new_n558));
  NAND2_X1  g357(.A1(G225gat), .A2(G233gat), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n524), .A2(new_n527), .A3(new_n378), .A4(new_n381), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n433), .A2(new_n494), .A3(KEYINPUT4), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n558), .A2(new_n559), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT5), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n382), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n560), .ZN(new_n567));
  INV_X1    g366(.A(new_n559), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n562), .A2(new_n563), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n571), .A2(new_n565), .A3(new_n559), .A4(new_n558), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G1gat), .B(G29gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT0), .ZN(new_n575));
  XNOR2_X1  g374(.A(G57gat), .B(G85gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT6), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(new_n572), .A3(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G226gat), .A2(G233gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n430), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT25), .B1(new_n587), .B2(new_n397), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n398), .A2(new_n406), .A3(KEYINPUT25), .A4(new_n407), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n400), .B2(new_n404), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n439), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n586), .B1(new_n591), .B2(new_n495), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n585), .B1(new_n432), .B2(new_n439), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n533), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n420), .A2(new_n422), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n428), .A2(new_n431), .B1(new_n595), .B2(new_n436), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n585), .B1(new_n596), .B2(KEYINPUT29), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n591), .A2(new_n586), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(new_n521), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G8gat), .B(G36gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT71), .ZN(new_n601));
  XNOR2_X1  g400(.A(G64gat), .B(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n594), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT30), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(KEYINPUT73), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n594), .A2(new_n599), .A3(KEYINPUT30), .A4(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n594), .A2(KEYINPUT70), .A3(new_n599), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT70), .B1(new_n594), .B2(new_n599), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n603), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n584), .A2(new_n611), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT35), .B1(new_n556), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g418(.A1(new_n584), .A2(new_n611), .A3(new_n614), .A4(new_n617), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT35), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n549), .A2(new_n552), .ZN(new_n622));
  INV_X1    g421(.A(new_n553), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n472), .A2(new_n469), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n620), .A2(new_n621), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n554), .A2(new_n555), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT68), .B(KEYINPUT36), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n472), .A2(new_n469), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(KEYINPUT68), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n468), .B1(new_n463), .B2(new_n466), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n630), .A2(new_n618), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT70), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n592), .A2(new_n533), .A3(new_n593), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n521), .B1(new_n597), .B2(new_n598), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n594), .A2(KEYINPUT70), .A3(new_n599), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n594), .A2(new_n641), .A3(new_n599), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n603), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT38), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n605), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n594), .A2(new_n599), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT38), .B1(new_n653), .B2(KEYINPUT37), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n650), .A2(new_n655), .A3(new_n583), .A4(new_n582), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n558), .A2(new_n562), .A3(new_n563), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT39), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n568), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n577), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT39), .B1(new_n567), .B2(new_n568), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n568), .B2(new_n658), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n568), .ZN(new_n665));
  INV_X1    g464(.A(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(KEYINPUT40), .A3(new_n577), .A4(new_n660), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n668), .A3(new_n579), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n605), .A2(KEYINPUT73), .A3(new_n606), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT73), .B1(new_n605), .B2(new_n606), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n617), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n612), .B(KEYINPUT72), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n656), .A2(new_n675), .A3(new_n626), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n619), .A2(new_n629), .B1(new_n640), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G113gat), .B(G141gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G197gat), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT11), .B(G169gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT12), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT83), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n320), .B(G8gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n275), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n279), .B2(new_n280), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n322), .A2(new_n270), .ZN(new_n687));
  NAND2_X1  g486(.A1(G229gat), .A2(G233gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(KEYINPUT18), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n683), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n322), .B1(KEYINPUT17), .B2(new_n263), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n272), .B2(new_n273), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n687), .A2(KEYINPUT18), .A3(new_n688), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT83), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n684), .A2(new_n263), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n688), .B(KEYINPUT13), .Z(new_n697));
  AOI22_X1  g496(.A1(new_n690), .A2(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT82), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n687), .A2(new_n688), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n692), .A2(KEYINPUT82), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT18), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n682), .B1(new_n698), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n696), .A2(new_n697), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n682), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n690), .B2(new_n694), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT84), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(KEYINPUT84), .A3(new_n705), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n706), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n677), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT94), .B1(new_n367), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n367), .A2(KEYINPUT94), .A3(new_n715), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n584), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g521(.A1(new_n673), .A2(new_n674), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n717), .B2(new_n718), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT16), .B(G8gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT97), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n724), .B2(new_n321), .ZN(new_n734));
  INV_X1    g533(.A(new_n718), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n716), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT97), .B(G8gat), .C1(new_n736), .C2(new_n723), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n723), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT95), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n740), .B(new_n741), .C1(new_n735), .C2(new_n716), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(KEYINPUT96), .A3(new_n726), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT96), .B1(new_n742), .B2(new_n726), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT99), .B1(new_n739), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT99), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n748), .A2(new_n749), .A3(new_n732), .A4(new_n738), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1325gat));
  NAND2_X1  g550(.A1(new_n639), .A2(new_n633), .ZN(new_n752));
  OAI21_X1  g551(.A(G15gat), .B1(new_n736), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n719), .A2(new_n452), .A3(new_n628), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1326gat));
  NAND2_X1  g554(.A1(new_n719), .A2(new_n630), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT43), .B(G22gat), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1327gat));
  NOR2_X1   g557(.A1(new_n334), .A2(new_n364), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n289), .A2(new_n292), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT100), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n715), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n720), .A3(new_n254), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n627), .B1(new_n625), .B2(new_n624), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n621), .B1(new_n766), .B2(new_n620), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n556), .A2(KEYINPUT35), .A3(new_n618), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n752), .B1(new_n620), .B2(new_n626), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT37), .B1(new_n643), .B2(new_n644), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT38), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n770), .A2(new_n771), .A3(new_n603), .A4(new_n648), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n582), .A2(new_n583), .A3(new_n772), .A4(new_n605), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT37), .B1(new_n615), .B2(new_n616), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n652), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n773), .A2(new_n775), .B1(new_n554), .B2(new_n555), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n604), .B1(new_n645), .B2(new_n646), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n609), .B2(new_n610), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n669), .B1(new_n778), .B2(new_n614), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT102), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n677), .A2(KEYINPUT102), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n760), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n760), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT101), .B1(new_n787), .B2(KEYINPUT44), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT101), .B(KEYINPUT44), .C1(new_n677), .C2(new_n293), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n786), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n714), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n759), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n720), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n765), .B1(new_n254), .B2(new_n794), .ZN(G1328gat));
  NAND4_X1  g594(.A1(new_n762), .A2(new_n235), .A3(new_n740), .A4(new_n715), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT46), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT104), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n793), .A2(new_n740), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n799), .C1(new_n235), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n235), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT104), .B1(new_n802), .B2(new_n797), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1329gat));
  NAND4_X1  g603(.A1(new_n762), .A2(new_n231), .A3(new_n628), .A4(new_n715), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT105), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n807));
  INV_X1    g606(.A(new_n752), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n231), .B1(new_n793), .B2(new_n808), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n806), .B2(new_n809), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1330gat));
  NOR2_X1   g611(.A1(new_n626), .A2(G50gat), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT106), .B1(new_n763), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n814), .A2(KEYINPUT48), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n793), .A2(new_n630), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n816), .A2(G50gat), .B1(new_n763), .B2(new_n813), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n815), .B(new_n817), .ZN(G1331gat));
  NAND4_X1  g617(.A1(new_n293), .A2(new_n334), .A3(new_n714), .A4(new_n364), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n783), .A2(new_n784), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n720), .ZN(new_n822));
  XNOR2_X1  g621(.A(KEYINPUT107), .B(G57gat), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n822), .B(new_n823), .ZN(G1332gat));
  AOI21_X1  g623(.A(new_n723), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT108), .ZN(new_n827));
  NOR2_X1   g626(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n827), .B(new_n828), .ZN(G1333gat));
  INV_X1    g628(.A(G71gat), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n821), .A2(new_n830), .A3(new_n628), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n820), .A2(new_n752), .A3(new_n819), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n830), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g633(.A1(new_n821), .A2(new_n630), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(G78gat), .ZN(G1335gat));
  INV_X1    g635(.A(KEYINPUT109), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n333), .A2(new_n714), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n365), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n791), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n840), .B2(new_n584), .ZN(new_n841));
  INV_X1    g640(.A(new_n839), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT44), .B1(new_n677), .B2(new_n293), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n789), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n846), .B2(new_n786), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(KEYINPUT109), .A3(new_n720), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n841), .A2(G85gat), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n781), .A2(new_n760), .A3(new_n714), .A4(new_n333), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n850), .A2(KEYINPUT110), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT110), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n850), .A2(new_n851), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n855), .A2(new_n211), .A3(new_n720), .A4(new_n364), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n849), .A2(new_n856), .ZN(G1336gat));
  NOR3_X1   g656(.A1(new_n723), .A2(G92gat), .A3(new_n365), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT52), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n791), .A2(new_n740), .A3(new_n839), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G92gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n863));
  NOR2_X1   g662(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n850), .B(new_n864), .Z(new_n865));
  INV_X1    g664(.A(new_n858), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n860), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n870));
  AOI211_X1 g669(.A(KEYINPUT113), .B(new_n863), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n723), .B(new_n842), .C1(new_n846), .C2(new_n786), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n868), .B1(new_n873), .B2(new_n212), .ZN(new_n874));
  INV_X1    g673(.A(new_n867), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n872), .B1(new_n876), .B2(KEYINPUT52), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n862), .B1(new_n871), .B2(new_n877), .ZN(G1337gat));
  XOR2_X1   g677(.A(KEYINPUT115), .B(G99gat), .Z(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n627), .A2(new_n365), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n855), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT114), .B1(new_n840), .B2(new_n752), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n847), .A2(new_n884), .A3(new_n808), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n882), .B1(new_n886), .B2(new_n880), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT116), .ZN(G1338gat));
  NAND3_X1  g687(.A1(new_n791), .A2(new_n630), .A3(new_n839), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G106gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n626), .A2(G106gat), .A3(new_n365), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n855), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n896));
  INV_X1    g695(.A(new_n891), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n865), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n890), .B2(KEYINPUT117), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n889), .A2(new_n900), .A3(G106gat), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n895), .B(new_n896), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n626), .B(new_n842), .C1(new_n846), .C2(new_n786), .ZN(new_n903));
  INV_X1    g702(.A(G106gat), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT117), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n898), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT118), .B1(new_n907), .B2(KEYINPUT53), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n894), .B1(new_n902), .B2(new_n908), .ZN(G1339gat));
  NAND2_X1  g708(.A1(new_n367), .A2(new_n714), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n362), .B1(new_n360), .B2(KEYINPUT54), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT54), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n339), .A2(new_n345), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n352), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n354), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n354), .A2(new_n914), .A3(KEYINPUT120), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT55), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT55), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n911), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n918), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT120), .B1(new_n354), .B2(new_n914), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n359), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n712), .A2(new_n713), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n688), .B1(new_n692), .B2(new_n687), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n696), .A2(new_n697), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n681), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n920), .A2(new_n926), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n293), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n709), .A2(KEYINPUT84), .A3(new_n705), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT84), .B1(new_n709), .B2(new_n705), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n364), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n925), .B(new_n359), .C1(new_n919), .C2(KEYINPUT55), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n714), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n937), .A2(KEYINPUT121), .B1(new_n292), .B2(new_n289), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n935), .B(new_n939), .C1(new_n714), .C2(new_n936), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n932), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n910), .B1(new_n941), .B2(new_n334), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n740), .A2(new_n584), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n942), .A2(new_n626), .A3(new_n628), .A4(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n370), .A3(new_n714), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n937), .A2(KEYINPUT121), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(new_n293), .A3(new_n940), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n293), .A2(new_n931), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n334), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n366), .A2(new_n792), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n584), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n740), .A2(new_n556), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n792), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n945), .B1(new_n956), .B2(new_n370), .ZN(G1340gat));
  NOR3_X1   g756(.A1(new_n944), .A2(new_n368), .A3(new_n365), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n364), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n368), .ZN(G1341gat));
  OAI21_X1  g759(.A(G127gat), .B1(new_n944), .B2(new_n333), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n334), .A2(new_n376), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n954), .B2(new_n962), .ZN(G1342gat));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n374), .A3(new_n760), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(KEYINPUT56), .ZN(new_n965));
  OAI21_X1  g764(.A(G134gat), .B1(new_n944), .B2(new_n293), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(KEYINPUT56), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(G1343gat));
  NOR3_X1   g767(.A1(new_n808), .A2(new_n740), .A3(new_n626), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n969), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n970), .A2(G141gat), .A3(new_n714), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT58), .ZN(new_n972));
  INV_X1    g771(.A(new_n943), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n973), .A2(new_n808), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT57), .B1(new_n942), .B2(new_n630), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n630), .A2(KEYINPUT57), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n293), .A2(new_n937), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n333), .B1(new_n977), .B2(new_n932), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n978), .B2(new_n910), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n974), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(G141gat), .B1(new_n980), .B2(new_n714), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n630), .B1(new_n949), .B2(new_n950), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT57), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(new_n974), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT122), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n988), .B(new_n974), .C1(new_n975), .C2(new_n979), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(new_n792), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n971), .B1(new_n990), .B2(G141gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT58), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n982), .B1(new_n991), .B2(new_n992), .ZN(G1344gat));
  INV_X1    g792(.A(KEYINPUT59), .ZN(new_n994));
  INV_X1    g793(.A(new_n970), .ZN(new_n995));
  AOI211_X1 g794(.A(new_n994), .B(G148gat), .C1(new_n995), .C2(new_n364), .ZN(new_n996));
  INV_X1    g795(.A(G148gat), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n978), .A2(new_n910), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n984), .B1(new_n998), .B2(new_n626), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n942), .A2(KEYINPUT57), .A3(new_n630), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n1001), .A2(new_n364), .A3(new_n974), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n997), .B1(new_n1002), .B2(KEYINPUT59), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n987), .A2(new_n989), .A3(new_n994), .A4(new_n364), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n996), .B1(new_n1003), .B2(new_n1004), .ZN(G1345gat));
  NAND3_X1  g804(.A1(new_n987), .A2(new_n334), .A3(new_n989), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G155gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n995), .A2(new_n327), .A3(new_n334), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1346gat));
  AOI21_X1  g808(.A(G162gat), .B1(new_n995), .B2(new_n760), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n987), .A2(new_n989), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n760), .A2(G162gat), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(G1347gat));
  NOR2_X1   g812(.A1(new_n723), .A2(new_n720), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n942), .A2(new_n626), .A3(new_n628), .A4(new_n1014), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1015), .A2(new_n385), .A3(new_n714), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n951), .A2(new_n720), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n556), .A2(new_n723), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(KEYINPUT123), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n1017), .A2(new_n792), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1016), .B1(new_n385), .B2(new_n1020), .ZN(G1348gat));
  OAI21_X1  g820(.A(G176gat), .B1(new_n1015), .B2(new_n365), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n942), .A2(new_n584), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n364), .A2(new_n386), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(G1349gat));
  OAI21_X1  g824(.A(G183gat), .B1(new_n1015), .B2(new_n333), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n334), .A2(new_n421), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1026), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g827(.A(new_n1028), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g828(.A(KEYINPUT124), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n760), .A2(new_n394), .ZN(new_n1031));
  OR3_X1    g830(.A1(new_n1023), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1030), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g833(.A(KEYINPUT61), .B(G190gat), .C1(new_n1015), .C2(new_n293), .ZN(new_n1035));
  OAI21_X1  g834(.A(G190gat), .B1(new_n1015), .B2(new_n293), .ZN(new_n1036));
  INV_X1    g835(.A(KEYINPUT61), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1039), .A2(KEYINPUT125), .ZN(new_n1040));
  INV_X1    g839(.A(KEYINPUT125), .ZN(new_n1041));
  NAND4_X1  g840(.A1(new_n1034), .A2(new_n1041), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1040), .A2(new_n1042), .ZN(G1351gat));
  NOR3_X1   g842(.A1(new_n808), .A2(new_n723), .A3(new_n626), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n1017), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g844(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1046), .A2(new_n504), .A3(new_n792), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1014), .A2(new_n752), .ZN(new_n1048));
  AOI211_X1 g847(.A(new_n714), .B(new_n1048), .C1(new_n999), .C2(new_n1000), .ZN(new_n1049));
  AND2_X1   g848(.A1(new_n1049), .A2(KEYINPUT126), .ZN(new_n1050));
  OAI21_X1  g849(.A(G197gat), .B1(new_n1049), .B2(KEYINPUT126), .ZN(new_n1051));
  OAI21_X1  g850(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(G1352gat));
  NAND4_X1  g851(.A1(new_n1017), .A2(new_n505), .A3(new_n364), .A4(new_n1044), .ZN(new_n1053));
  XOR2_X1   g852(.A(new_n1053), .B(KEYINPUT62), .Z(new_n1054));
  AOI211_X1 g853(.A(new_n365), .B(new_n1048), .C1(new_n999), .C2(new_n1000), .ZN(new_n1055));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1056));
  OAI21_X1  g855(.A(G204gat), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g857(.A(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(G1353gat));
  NAND3_X1  g858(.A1(new_n1046), .A2(new_n511), .A3(new_n334), .ZN(new_n1060));
  AOI21_X1  g859(.A(new_n1048), .B1(new_n999), .B2(new_n1000), .ZN(new_n1061));
  NAND2_X1  g860(.A1(new_n1061), .A2(new_n334), .ZN(new_n1062));
  AND3_X1   g861(.A1(new_n1062), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1063));
  AOI21_X1  g862(.A(KEYINPUT63), .B1(new_n1062), .B2(G211gat), .ZN(new_n1064));
  OAI21_X1  g863(.A(new_n1060), .B1(new_n1063), .B2(new_n1064), .ZN(G1354gat));
  NAND3_X1  g864(.A1(new_n1046), .A2(new_n512), .A3(new_n760), .ZN(new_n1066));
  AND2_X1   g865(.A1(new_n1061), .A2(new_n760), .ZN(new_n1067));
  OAI21_X1  g866(.A(new_n1066), .B1(new_n1067), .B2(new_n512), .ZN(G1355gat));
endmodule


