

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  NOR2_X1 U322 ( .A1(n513), .A2(n524), .ZN(n392) );
  NOR2_X1 U323 ( .A1(n390), .A2(n389), .ZN(n391) );
  XOR2_X2 U324 ( .A(n417), .B(n361), .Z(n571) );
  NOR2_X1 U325 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U326 ( .A(n416), .B(KEYINPUT65), .ZN(n566) );
  XNOR2_X1 U327 ( .A(n391), .B(KEYINPUT48), .ZN(n524) );
  OR2_X1 U328 ( .A1(n383), .A2(n382), .ZN(n385) );
  XOR2_X1 U329 ( .A(G92GAT), .B(G64GAT), .Z(n348) );
  XNOR2_X1 U330 ( .A(n358), .B(KEYINPUT73), .ZN(n359) );
  XNOR2_X1 U331 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U332 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT75), .B(KEYINPUT71), .Z(n291) );
  XNOR2_X1 U335 ( .A(G218GAT), .B(G92GAT), .ZN(n290) );
  XNOR2_X1 U336 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U337 ( .A(n292), .B(KEYINPUT11), .Z(n294) );
  XOR2_X1 U338 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n342) );
  XNOR2_X1 U339 ( .A(n342), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U341 ( .A(G29GAT), .B(KEYINPUT76), .Z(n396) );
  XOR2_X1 U342 ( .A(G50GAT), .B(G162GAT), .Z(n423) );
  XOR2_X1 U343 ( .A(n396), .B(n423), .Z(n296) );
  NAND2_X1 U344 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U346 ( .A(KEYINPUT67), .B(KEYINPUT74), .Z(n298) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G85GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U349 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U350 ( .A(G43GAT), .B(G134GAT), .Z(n440) );
  XOR2_X1 U351 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n302) );
  XNOR2_X1 U352 ( .A(G190GAT), .B(G106GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n440), .B(n303), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n551) );
  XOR2_X1 U357 ( .A(G183GAT), .B(KEYINPUT84), .Z(n309) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n311) );
  XNOR2_X1 U361 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(n313), .B(n312), .Z(n438) );
  XOR2_X1 U364 ( .A(n348), .B(KEYINPUT77), .Z(n315) );
  NAND2_X1 U365 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U367 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n317) );
  XNOR2_X1 U368 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n326) );
  XOR2_X1 U371 ( .A(G36GAT), .B(G8GAT), .Z(n341) );
  XOR2_X1 U372 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n321) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(KEYINPUT91), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n322), .B(KEYINPUT90), .Z(n324) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n428) );
  XNOR2_X1 U378 ( .A(n341), .B(n428), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n438), .B(n327), .ZN(n513) );
  XOR2_X1 U381 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n329) );
  NAND2_X1 U382 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(n330), .B(KEYINPUT69), .Z(n338) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G29GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(G43GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U388 ( .A(KEYINPUT30), .B(G197GAT), .Z(n334) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G141GAT), .ZN(n333) );
  XNOR2_X1 U390 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n340) );
  XNOR2_X1 U393 ( .A(G15GAT), .B(G22GAT), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n339), .B(G1GAT), .ZN(n369) );
  XOR2_X1 U395 ( .A(n340), .B(n369), .Z(n344) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n568) );
  INV_X1 U398 ( .A(n568), .ZN(n529) );
  XNOR2_X1 U399 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n362) );
  XOR2_X1 U400 ( .A(G148GAT), .B(G106GAT), .Z(n346) );
  XNOR2_X1 U401 ( .A(G204GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U403 ( .A(KEYINPUT70), .B(n347), .Z(n417) );
  XOR2_X1 U404 ( .A(KEYINPUT71), .B(n348), .Z(n350) );
  XOR2_X1 U405 ( .A(G85GAT), .B(G57GAT), .Z(n397) );
  XNOR2_X1 U406 ( .A(G120GAT), .B(n397), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U408 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n352) );
  XNOR2_X1 U409 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n351) );
  XOR2_X1 U410 ( .A(n352), .B(n351), .Z(n353) );
  XNOR2_X1 U411 ( .A(n354), .B(n353), .ZN(n356) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n360) );
  XNOR2_X1 U414 ( .A(G99GAT), .B(G71GAT), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n357), .B(G176GAT), .ZN(n439) );
  XOR2_X1 U416 ( .A(n439), .B(KEYINPUT33), .Z(n358) );
  XNOR2_X1 U417 ( .A(n362), .B(n571), .ZN(n495) );
  AND2_X1 U418 ( .A1(n529), .A2(n495), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n363), .B(KEYINPUT46), .ZN(n383) );
  XOR2_X1 U420 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n365) );
  XNOR2_X1 U421 ( .A(KEYINPUT13), .B(KEYINPUT78), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n373) );
  XOR2_X1 U423 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n371) );
  XOR2_X1 U424 ( .A(KEYINPUT77), .B(G64GAT), .Z(n367) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G57GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n381) );
  NAND2_X1 U430 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XOR2_X1 U431 ( .A(G78GAT), .B(G211GAT), .Z(n375) );
  XNOR2_X1 U432 ( .A(G183GAT), .B(G155GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U434 ( .A(G127GAT), .B(G71GAT), .Z(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n533) );
  INV_X1 U438 ( .A(n533), .ZN(n574) );
  NAND2_X1 U439 ( .A1(n574), .A2(n551), .ZN(n382) );
  XOR2_X1 U440 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n390) );
  INV_X1 U442 ( .A(n551), .ZN(n538) );
  XNOR2_X1 U443 ( .A(n538), .B(KEYINPUT36), .ZN(n577) );
  NAND2_X1 U444 ( .A1(n533), .A2(n577), .ZN(n386) );
  XNOR2_X1 U445 ( .A(KEYINPUT45), .B(n386), .ZN(n388) );
  NAND2_X1 U446 ( .A1(n571), .A2(n568), .ZN(n387) );
  NOR2_X1 U447 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n392), .B(KEYINPUT54), .ZN(n415) );
  XOR2_X1 U449 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT92), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U452 ( .A(G141GAT), .B(n395), .Z(n432) );
  XOR2_X1 U453 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(G162GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U456 ( .A(n432), .B(n400), .Z(n402) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U459 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n404) );
  XNOR2_X1 U460 ( .A(G148GAT), .B(KEYINPUT1), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U462 ( .A(n406), .B(n405), .Z(n414) );
  XOR2_X1 U463 ( .A(KEYINPUT81), .B(G127GAT), .Z(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U466 ( .A(G113GAT), .B(n409), .Z(n446) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n411) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n446), .B(n412), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n467) );
  XNOR2_X1 U472 ( .A(KEYINPUT96), .B(n467), .ZN(n510) );
  NAND2_X1 U473 ( .A1(n415), .A2(n510), .ZN(n416) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n419) );
  XNOR2_X1 U475 ( .A(n417), .B(KEYINPUT87), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n427) );
  XOR2_X1 U477 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n421) );
  XNOR2_X1 U478 ( .A(KEYINPUT93), .B(KEYINPUT88), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n430) );
  XNOR2_X1 U484 ( .A(G22GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n461) );
  NAND2_X1 U487 ( .A1(n566), .A2(n461), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n447) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT66), .Z(n436) );
  XNOR2_X1 U491 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n442) );
  NAND2_X1 U495 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n516) );
  NOR2_X1 U499 ( .A1(n447), .A2(n516), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n448), .B(KEYINPUT121), .ZN(n560) );
  NOR2_X1 U501 ( .A1(n551), .A2(n560), .ZN(n452) );
  XNOR2_X1 U502 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n450) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n449) );
  AND2_X1 U504 ( .A1(n529), .A2(n571), .ZN(n484) );
  XOR2_X1 U505 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n454) );
  NAND2_X1 U506 ( .A1(n533), .A2(n551), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n470) );
  INV_X1 U508 ( .A(n510), .ZN(n543) );
  XNOR2_X1 U509 ( .A(KEYINPUT28), .B(n461), .ZN(n520) );
  AND2_X1 U510 ( .A1(n543), .A2(n520), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n513), .Z(n463) );
  NAND2_X1 U512 ( .A1(n455), .A2(n463), .ZN(n525) );
  XNOR2_X1 U513 ( .A(KEYINPUT85), .B(n516), .ZN(n456) );
  NOR2_X1 U514 ( .A1(n525), .A2(n456), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n457), .B(KEYINPUT99), .ZN(n469) );
  OR2_X1 U516 ( .A1(n513), .A2(n516), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n458), .A2(n461), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U519 ( .A(KEYINPUT101), .B(n460), .ZN(n465) );
  INV_X1 U520 ( .A(n516), .ZN(n526) );
  NOR2_X1 U521 ( .A1(n526), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(KEYINPUT26), .B(n462), .ZN(n565) );
  NAND2_X1 U523 ( .A1(n565), .A2(n463), .ZN(n541) );
  XNOR2_X1 U524 ( .A(n541), .B(KEYINPUT100), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n481) );
  AND2_X1 U528 ( .A1(n470), .A2(n481), .ZN(n496) );
  NAND2_X1 U529 ( .A1(n484), .A2(n496), .ZN(n479) );
  NOR2_X1 U530 ( .A1(n510), .A2(n479), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U533 ( .A(G1GAT), .B(n473), .Z(G1324GAT) );
  NOR2_X1 U534 ( .A1(n513), .A2(n479), .ZN(n475) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1325GAT) );
  NOR2_X1 U537 ( .A1(n516), .A2(n479), .ZN(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n478), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n520), .A2(n479), .ZN(n480) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n480), .Z(G1327GAT) );
  NAND2_X1 U543 ( .A1(n577), .A2(n481), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n533), .A2(n482), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n483), .Z(n507) );
  NAND2_X1 U546 ( .A1(n484), .A2(n507), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n485), .B(KEYINPUT38), .ZN(n493) );
  NOR2_X1 U548 ( .A1(n510), .A2(n493), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n487) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT106), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n493), .A2(n513), .ZN(n490) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n493), .A2(n516), .ZN(n491) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(n491), .Z(n492) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n520), .A2(n493), .ZN(n494) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n494), .Z(G1331GAT) );
  INV_X1 U560 ( .A(n495), .ZN(n557) );
  NOR2_X1 U561 ( .A1(n529), .A2(n557), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n496), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n510), .A2(n503), .ZN(n498) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U565 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n513), .A2(n503), .ZN(n500) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n500), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n516), .A2(n503), .ZN(n501) );
  XOR2_X1 U570 ( .A(KEYINPUT108), .B(n501), .Z(n502) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n502), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n520), .A2(n503), .ZN(n505) );
  XNOR2_X1 U573 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n506), .Z(G1335GAT) );
  NAND2_X1 U576 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U577 ( .A(n509), .B(KEYINPUT110), .ZN(n519) );
  NOR2_X1 U578 ( .A1(n519), .A2(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NOR2_X1 U581 ( .A1(n519), .A2(n513), .ZN(n514) );
  XOR2_X1 U582 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n515), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(G1338GAT) );
  XNOR2_X1 U587 ( .A(KEYINPUT114), .B(KEYINPUT44), .ZN(n522) );
  NOR2_X1 U588 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n523), .Z(G1339GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n525), .ZN(n527) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT116), .B(n528), .Z(n537) );
  NAND2_X1 U594 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U597 ( .A1(n495), .A2(n537), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U600 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n524), .A2(n541), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n568), .A2(n550), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  NOR2_X1 U613 ( .A1(n557), .A2(n550), .ZN(n547) );
  XOR2_X1 U614 ( .A(n548), .B(n547), .Z(G1345GAT) );
  NOR2_X1 U615 ( .A1(n574), .A2(n550), .ZN(n549) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n568), .A2(n560), .ZN(n554) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n559) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1349GAT) );
  NOR2_X1 U626 ( .A1(n574), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(n567), .Z(n576) );
  NOR2_X1 U634 ( .A1(n568), .A2(n576), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n576), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n576), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  INV_X1 U642 ( .A(n576), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

