//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT68), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  OR3_X1    g036(.A1(new_n455), .A2(KEYINPUT68), .A3(new_n460), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(G319));
  AND2_X1   g039(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  INV_X1    g054(.A(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(new_n469), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(KEYINPUT71), .A3(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n485), .A2(new_n486), .B1(G136), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT4), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n467), .A2(new_n474), .A3(new_n469), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT72), .B1(new_n474), .B2(G114), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n498), .A3(G2105), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n496), .A2(new_n499), .A3(G2104), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT3), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(new_n503), .A3(G138), .A4(new_n474), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n493), .A2(new_n495), .A3(new_n501), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT73), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n510), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  INV_X1    g098(.A(new_n514), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n518), .A2(new_n523), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n522), .A2(G51), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n525), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n532), .B2(new_n514), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n525), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n526), .A2(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n526), .A2(new_n545), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT74), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n549), .B2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n522), .A2(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT77), .B1(new_n559), .B2(KEYINPUT76), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT79), .B(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n514), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n558), .A2(new_n561), .B1(new_n564), .B2(G651), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n560), .B1(KEYINPUT77), .B2(new_n559), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n527), .B2(G91), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  NOR3_X1   g144(.A1(new_n526), .A2(KEYINPUT78), .A3(new_n569), .ZN(new_n570));
  OAI221_X1 g145(.A(new_n565), .B1(new_n558), .B2(new_n566), .C1(new_n568), .C2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  OAI21_X1  g148(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n522), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n524), .A2(new_n525), .A3(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n514), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(G48), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n514), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(new_n525), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n590), .A2(G651), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n526), .A2(new_n593), .B1(new_n541), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n524), .A2(new_n525), .A3(G92), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n522), .A2(G54), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n538), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n598), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(new_n608), .B2(G168), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n549), .A2(G651), .ZN(new_n614));
  INV_X1    g189(.A(new_n547), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n608), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n604), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g195(.A1(new_n471), .A2(new_n475), .A3(new_n474), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n482), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n487), .A2(G135), .ZN(new_n626));
  NOR2_X1   g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(new_n474), .B2(G111), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2443), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  AND2_X1   g219(.A1(new_n644), .A2(G14), .ZN(G401));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT82), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT17), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2096), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  INV_X1    g231(.A(new_n652), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n656), .B1(new_n649), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(KEYINPUT20), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n661), .A3(new_n664), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n668), .B(new_n670), .C1(KEYINPUT20), .C2(new_n665), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1986), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1991), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n678), .A2(G24), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(G290), .B2(G16), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT35), .B(G1991), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n482), .A2(G119), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n487), .A2(G131), .ZN(new_n686));
  NOR2_X1   g261(.A1(G95), .A2(G2105), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(new_n474), .B2(G107), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n685), .B(new_n686), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(KEYINPUT84), .A2(G29), .ZN(new_n690));
  NOR2_X1   g265(.A1(KEYINPUT84), .A2(G29), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n689), .S(new_n692), .Z(new_n693));
  OAI211_X1 g268(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n678), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n678), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT33), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1976), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n678), .A2(G6), .ZN(new_n700));
  INV_X1    g275(.A(G305), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n678), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT85), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n678), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n678), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n705), .B1(new_n707), .B2(G1971), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n699), .B(new_n708), .C1(G1971), .C2(new_n707), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n694), .B1(new_n709), .B2(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n693), .A2(new_n684), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n710), .B(new_n711), .C1(KEYINPUT34), .C2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT36), .ZN(new_n713));
  NOR2_X1   g288(.A1(G29), .A2(G33), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n487), .A2(G139), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT87), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  AOI22_X1  g293(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n718), .C1(new_n474), .C2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(G29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2072), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n678), .A2(G4), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n605), .B2(new_n678), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT86), .B(G1348), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n678), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n550), .B2(new_n678), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(new_n727), .B1(G1341), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n692), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT24), .B(G34), .ZN(new_n732));
  AOI22_X1  g307(.A1(G160), .A2(G29), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n730), .B1(G1341), .B2(new_n729), .C1(G2084), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G2084), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT89), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n731), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n731), .ZN(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT28), .B1(new_n731), .B2(G26), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n731), .A2(KEYINPUT28), .A3(G26), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G128), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n487), .A2(G140), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n742), .B(new_n744), .C1(new_n749), .C2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n678), .A2(G21), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G168), .B2(new_n678), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G5), .A2(G16), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G171), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  INV_X1    g334(.A(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT90), .B(G28), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT30), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n629), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n757), .A2(G1961), .B1(new_n764), .B2(new_n692), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n755), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n482), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT26), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n471), .A2(G105), .A3(new_n474), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n767), .A2(new_n768), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G32), .B(new_n772), .S(G29), .Z(new_n773));
  XOR2_X1   g348(.A(KEYINPUT27), .B(G1996), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR3_X1   g351(.A1(new_n766), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n737), .A2(new_n741), .A3(new_n751), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2090), .ZN(new_n779));
  INV_X1    g354(.A(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT91), .B1(new_n692), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g356(.A1(new_n692), .A2(KEYINPUT91), .A3(new_n780), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G162), .C2(new_n731), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n724), .B(new_n778), .C1(new_n779), .C2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n726), .A2(new_n727), .ZN(new_n787));
  NAND2_X1  g362(.A1(G299), .A2(G16), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT93), .B(KEYINPUT23), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n678), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  INV_X1    g368(.A(new_n785), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n713), .A2(new_n786), .A3(new_n787), .A4(new_n796), .ZN(G150));
  INV_X1    g372(.A(G150), .ZN(G311));
  INV_X1    g373(.A(G93), .ZN(new_n799));
  INV_X1    g374(.A(G55), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n526), .A2(new_n799), .B1(new_n541), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  INV_X1    g380(.A(G67), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n514), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G651), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT96), .B(G860), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n809), .A2(new_n550), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n802), .A2(new_n803), .B1(G651), .B2(new_n807), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n616), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT39), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n605), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n812), .B1(new_n820), .B2(new_n810), .ZN(G145));
  XOR2_X1   g396(.A(new_n491), .B(G160), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n772), .B(new_n749), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n495), .A2(new_n506), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n493), .A2(KEYINPUT97), .A3(new_n501), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT97), .B1(new_n493), .B2(new_n501), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n823), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(new_n720), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT98), .ZN(new_n831));
  INV_X1    g406(.A(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n722), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n834), .A3(new_n720), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n482), .A2(G130), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n487), .A2(G142), .ZN(new_n838));
  NOR2_X1   g413(.A1(G106), .A2(G2105), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(new_n474), .B2(G118), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n622), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n836), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n629), .B(new_n689), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n831), .A2(new_n833), .A3(new_n845), .A4(new_n835), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n844), .B1(new_n843), .B2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n822), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  INV_X1    g426(.A(new_n822), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g431(.A1(new_n809), .A2(new_n608), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n816), .B(new_n618), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n604), .A2(G299), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n604), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT99), .Z(new_n864));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n866), .B2(new_n858), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  XNOR2_X1  g443(.A(G290), .B(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(G288), .B(G305), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  OAI21_X1  g448(.A(G303), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n869), .A2(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n871), .A3(G166), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT101), .B1(new_n874), .B2(new_n876), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT101), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n882), .B2(KEYINPUT42), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n867), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n857), .B1(new_n884), .B2(new_n608), .ZN(G295));
  OAI21_X1  g460(.A(new_n857), .B1(new_n884), .B2(new_n608), .ZN(G331));
  NAND3_X1  g461(.A1(new_n813), .A2(new_n815), .A3(G301), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G301), .B1(new_n813), .B2(new_n815), .ZN(new_n889));
  OAI21_X1  g464(.A(G286), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(G168), .A3(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n866), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n892), .A3(new_n862), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n854), .B1(new_n897), .B2(new_n882), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n899));
  INV_X1    g474(.A(new_n881), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n879), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT102), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n895), .A2(KEYINPUT103), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n866), .B1(new_n890), .B2(new_n892), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n907), .A3(new_n896), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n898), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT104), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n907), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n901), .B(new_n902), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n895), .A2(new_n896), .ZN(new_n915));
  INV_X1    g490(.A(new_n882), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n898), .B1(new_n903), .B2(new_n897), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n910), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n911), .A2(new_n920), .A3(KEYINPUT44), .A4(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n903), .A2(new_n897), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n910), .B1(new_n926), .B2(new_n917), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(G397));
  NOR2_X1   g504(.A1(new_n749), .A2(G2067), .ZN(new_n930));
  INV_X1    g505(.A(G2067), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n749), .B(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n772), .B(G1996), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n689), .A2(new_n684), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n828), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n828), .A2(KEYINPUT105), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G40), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n473), .A2(new_n945), .A3(new_n478), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n937), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(G1996), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n948), .B1(new_n772), .B2(new_n933), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(KEYINPUT46), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  INV_X1    g531(.A(new_n935), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n689), .B(new_n684), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n948), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n592), .A2(new_n681), .A3(new_n596), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT48), .Z(new_n962));
  AOI211_X1 g537(.A(new_n950), .B(new_n956), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT63), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT55), .Z(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n947), .B1(new_n939), .B2(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n507), .A2(new_n938), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(KEYINPUT50), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G2090), .ZN(new_n971));
  INV_X1    g546(.A(G1971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n828), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n942), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n946), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n971), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G8), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n967), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n969), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n947), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n828), .A2(new_n986), .A3(new_n938), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n779), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n975), .A2(new_n989), .A3(new_n972), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n980), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n966), .A3(G8), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n828), .A2(new_n938), .A3(new_n946), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(G288), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n696), .A2(KEYINPUT110), .A3(G1976), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(G8), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(G288), .A2(new_n995), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n998), .A2(KEYINPUT52), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n998), .A2(KEYINPUT52), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT111), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n998), .A2(KEYINPUT52), .A3(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G305), .A2(G1981), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n581), .B2(new_n585), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(KEYINPUT49), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n993), .A4(G8), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1003), .A2(new_n1006), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n978), .A2(new_n992), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT109), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n982), .B(new_n986), .C1(new_n507), .C2(new_n938), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n987), .B(new_n946), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(G2084), .ZN(new_n1024));
  INV_X1    g599(.A(G2084), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n985), .A2(KEYINPUT115), .A3(new_n1025), .A4(new_n987), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n969), .A2(new_n942), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n493), .A2(new_n501), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT97), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n493), .A2(KEYINPUT97), .A3(new_n501), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n1032), .B2(new_n825), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n946), .B(new_n1027), .C1(new_n1033), .C2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n754), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1024), .A2(new_n1026), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(G8), .A3(G168), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n964), .B1(new_n1019), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  INV_X1    g614(.A(new_n992), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1003), .A2(new_n1006), .A3(new_n1017), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n1037), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n991), .A2(G8), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n964), .B1(new_n1043), .B2(new_n967), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1039), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1037), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1018), .A2(new_n1046), .A3(new_n992), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n967), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT63), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1047), .A2(new_n1049), .A3(KEYINPUT116), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1038), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1018), .A2(new_n1040), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1007), .B(KEYINPUT113), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(G1976), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1017), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(new_n1055), .B(KEYINPUT114), .Z(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(G8), .A3(new_n993), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1024), .A2(new_n1026), .A3(G168), .A4(new_n1035), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1036), .A2(G286), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1060), .B2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1059), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1036), .B2(G286), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1061), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1071), .A2(KEYINPUT124), .A3(new_n1067), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT62), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n973), .A2(new_n740), .A3(new_n974), .A4(new_n946), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(KEYINPUT126), .A3(new_n1075), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1023), .A2(new_n759), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT125), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1034), .B2(G2078), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT45), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n947), .B1(new_n939), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT125), .A3(new_n740), .A4(new_n1027), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(KEYINPUT53), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G301), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1065), .A2(new_n1059), .A3(new_n1068), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT124), .B1(new_n1071), .B2(new_n1067), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1073), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  NAND2_X1  g670(.A1(G299), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT57), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n973), .A2(new_n974), .A3(new_n946), .A4(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT117), .B(G1956), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n970), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1097), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n605), .ZN(new_n1105));
  INV_X1    g680(.A(new_n727), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1023), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1033), .A2(new_n1108), .A3(new_n946), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n993), .A2(KEYINPUT120), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n931), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1103), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1107), .A2(new_n1111), .A3(KEYINPUT60), .A4(new_n605), .ZN(new_n1117));
  AOI22_X1  g692(.A1(KEYINPUT61), .A2(new_n1104), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT58), .B(G1341), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT121), .B(G1996), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n975), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n975), .A2(new_n1124), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT122), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1119), .B1(new_n1129), .B2(new_n550), .ZN(new_n1130));
  AOI211_X1 g705(.A(KEYINPUT59), .B(new_n616), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1118), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n1104), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1113), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n947), .B1(new_n1033), .B2(KEYINPUT45), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n944), .A2(KEYINPUT53), .A3(new_n740), .A4(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1078), .A2(new_n1139), .A3(new_n1081), .A4(new_n1079), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1137), .B1(new_n1140), .B2(G171), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1080), .A2(G301), .A3(new_n1081), .A4(new_n1088), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1140), .A2(G171), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1137), .B1(new_n1089), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1135), .A2(new_n1136), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1094), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1019), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1058), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n960), .A2(KEYINPUT107), .ZN(new_n1153));
  NAND2_X1  g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1153), .B(new_n1154), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n959), .B1(new_n949), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n963), .B1(new_n1152), .B2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g732(.A1(G229), .A2(new_n463), .ZN(new_n1159));
  OAI21_X1  g733(.A(new_n1159), .B1(new_n925), .B2(new_n927), .ZN(new_n1160));
  NOR2_X1   g734(.A1(G401), .A2(G227), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n855), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1162), .ZN(G308));
  NAND2_X1  g737(.A1(new_n909), .A2(new_n910), .ZN(new_n1164));
  OAI21_X1  g738(.A(new_n1164), .B1(new_n910), .B2(new_n921), .ZN(new_n1165));
  NAND4_X1  g739(.A1(new_n1165), .A2(new_n855), .A3(new_n1159), .A4(new_n1161), .ZN(G225));
endmodule


