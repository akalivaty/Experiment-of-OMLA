//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898;
  NAND3_X1  g000(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT7), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT8), .ZN(new_n205));
  AND2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206));
  OAI221_X1 g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(G85gat), .C2(G92gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G99gat), .B(G106gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n210), .A2(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NOR3_X1   g013(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT104), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n213), .B(new_n214), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n219), .A2(new_n215), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n202), .B(new_n226), .C1(new_n228), .C2(new_n209), .ZN(new_n229));
  XOR2_X1   g028(.A(G190gat), .B(G218gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT110), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G134gat), .B(G162gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n233), .B(new_n234), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n232), .B(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n230), .A2(KEYINPUT110), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G71gat), .A2(G78gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT108), .B1(G71gat), .B2(G78gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(KEYINPUT108), .A2(G71gat), .A3(G78gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n244), .A2(KEYINPUT109), .ZN(new_n245));
  XOR2_X1   g044(.A(G57gat), .B(G64gat), .Z(new_n246));
  INV_X1    g045(.A(new_n240), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(KEYINPUT9), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(KEYINPUT109), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT9), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n251), .A2(G71gat), .A3(G78gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n246), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT21), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G15gat), .B(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT16), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(G1gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G1gat), .B2(new_n257), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(G8gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G183gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n254), .A2(new_n255), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n266), .B(G211gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n265), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G155gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(G231gat), .A2(G233gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n272), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n239), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n209), .A2(new_n253), .A3(new_n250), .ZN(new_n276));
  INV_X1    g075(.A(new_n208), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n207), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n254), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT10), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(KEYINPUT111), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n281), .A3(new_n279), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT111), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n276), .A2(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G230gat), .A2(G233gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G120gat), .B(G148gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G176gat), .B(G204gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n289), .B(new_n293), .C1(new_n280), .C2(new_n288), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n287), .A2(KEYINPUT112), .A3(new_n288), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT112), .B1(new_n287), .B2(new_n288), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n288), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n298), .B2(new_n293), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n275), .A2(KEYINPUT113), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT113), .B1(new_n275), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(KEYINPUT88), .B(KEYINPUT2), .Z(new_n307));
  XNOR2_X1  g106(.A(G141gat), .B(G148gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT89), .ZN(new_n310));
  INV_X1    g109(.A(new_n308), .ZN(new_n311));
  NOR3_X1   g110(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT85), .B(KEYINPUT29), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT84), .B(G211gat), .Z(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G218gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G211gat), .B(G218gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n321), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n315), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n313), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n317), .B1(new_n330), .B2(KEYINPUT96), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n326), .A2(new_n329), .A3(new_n327), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(KEYINPUT96), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n315), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT92), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n333), .B(new_n342), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n341), .A2(new_n343), .B1(new_n330), .B2(new_n319), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n335), .B(KEYINPUT95), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G22gat), .ZN(new_n347));
  INV_X1    g146(.A(G22gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n337), .B(new_n348), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n346), .B2(G22gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT31), .B(G50gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n350), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n347), .A2(new_n349), .A3(new_n351), .A4(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  INV_X1    g159(.A(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT78), .B(G71gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G169gat), .ZN(new_n366));
  INV_X1    g165(.A(G176gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT23), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT67), .B(G176gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI22_X1  g178(.A1(KEYINPUT66), .A2(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n380));
  OAI221_X1 g179(.A(new_n371), .B1(new_n372), .B2(new_n373), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n371), .B1(G176gat), .B2(new_n373), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT69), .B1(new_n374), .B2(KEYINPUT68), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT69), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(new_n376), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n376), .A2(new_n385), .B1(new_n388), .B2(new_n374), .ZN(new_n389));
  INV_X1    g188(.A(G190gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT70), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT70), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G190gat), .ZN(new_n393));
  AOI21_X1  g192(.A(G183gat), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT25), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n383), .B1(new_n384), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n370), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n374), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT71), .A2(G183gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT27), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT71), .A3(G183gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n392), .A2(G190gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT70), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n402), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT28), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n391), .B2(new_n393), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT27), .B(G183gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n400), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n369), .A2(KEYINPUT26), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n397), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n407), .A2(new_n408), .B1(new_n411), .B2(new_n410), .ZN(new_n416));
  INV_X1    g215(.A(new_n414), .ZN(new_n417));
  NOR4_X1   g216(.A1(new_n416), .A2(KEYINPUT72), .A3(new_n417), .A4(new_n400), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n396), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G113gat), .B(G120gat), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT73), .B1(new_n420), .B2(KEYINPUT1), .ZN(new_n421));
  XNOR2_X1  g220(.A(G127gat), .B(G134gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT73), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n425));
  INV_X1    g224(.A(G120gat), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n426), .A2(G113gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(G113gat), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n424), .B(new_n425), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n423), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT73), .B(new_n422), .C1(new_n420), .C2(KEYINPUT1), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT74), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT74), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n435), .A3(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n436), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT75), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n419), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT64), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n409), .A2(new_n412), .ZN(new_n445));
  INV_X1    g244(.A(new_n400), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n414), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT72), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n413), .A2(new_n397), .A3(new_n414), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n434), .B1(new_n433), .B2(new_n436), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n396), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n441), .A2(new_n444), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n441), .A2(new_n452), .A3(KEYINPUT76), .A4(new_n444), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n365), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n457), .B2(KEYINPUT32), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT32), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT77), .B(new_n462), .C1(new_n455), .C2(new_n456), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n466), .B(new_n459), .C1(new_n461), .C2(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n457), .B(KEYINPUT32), .C1(new_n458), .C2(new_n365), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n441), .A2(new_n452), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n443), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n442), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT80), .B(KEYINPUT34), .Z(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n474), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT82), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n470), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n486), .A2(new_n468), .A3(new_n469), .A4(new_n482), .ZN(new_n487));
  INV_X1    g286(.A(new_n469), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n465), .B2(new_n467), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n489), .B2(new_n482), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n359), .B(new_n485), .C1(new_n487), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n396), .A2(new_n447), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G226gat), .A2(G233gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(KEYINPUT29), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n495), .A2(new_n498), .B1(new_n419), .B2(new_n496), .ZN(new_n499));
  INV_X1    g298(.A(new_n330), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n497), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n419), .A2(new_n496), .A3(new_n318), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n330), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT86), .ZN(new_n506));
  XNOR2_X1  g305(.A(G64gat), .B(G92gat), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n506), .B(new_n507), .Z(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(KEYINPUT87), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n509), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n508), .B1(new_n501), .B2(new_n504), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(KEYINPUT87), .B2(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n433), .A2(new_n436), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n343), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g317(.A1(G225gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT91), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n314), .A2(new_n432), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n432), .B(KEYINPUT90), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n316), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n518), .A2(new_n521), .A3(new_n524), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n333), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n528), .B(KEYINPUT5), .C1(new_n521), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n517), .A2(new_n523), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n523), .B1(new_n314), .B2(new_n432), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT94), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n527), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT93), .B(KEYINPUT0), .Z(new_n538));
  XNOR2_X1  g337(.A(G1gat), .B(G29gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G85gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n531), .A2(new_n537), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT6), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n543), .B1(new_n531), .B2(new_n537), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n515), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n468), .A2(new_n469), .A3(new_n482), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT83), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n489), .A2(new_n486), .A3(new_n482), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n470), .A2(new_n480), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n551), .A3(new_n359), .A4(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n493), .A2(new_n551), .B1(new_n557), .B2(new_n492), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n485), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT36), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n531), .A2(new_n537), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n542), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n545), .B2(new_n544), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(new_n548), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n501), .B2(new_n504), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT101), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n566), .A2(new_n567), .A3(new_n508), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n566), .B2(new_n508), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n570));
  NAND3_X1  g369(.A1(new_n501), .A2(new_n565), .A3(new_n504), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n508), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n502), .A2(new_n503), .A3(new_n500), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n565), .B1(new_n499), .B2(new_n330), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n572), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n564), .A2(new_n578), .A3(new_n509), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n521), .B1(new_n535), .B2(new_n527), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT39), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n530), .A2(new_n521), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n542), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT99), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT40), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n547), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n587), .B(new_n515), .C1(new_n586), .C2(new_n585), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n579), .A2(new_n588), .A3(new_n359), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n357), .A2(new_n358), .ZN(new_n590));
  INV_X1    g389(.A(new_n515), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n563), .B2(new_n548), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n594), .B(new_n556), .C1(new_n487), .C2(new_n490), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n560), .A2(new_n589), .A3(new_n593), .A4(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n303), .B1(new_n558), .B2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G113gat), .B(G141gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT103), .ZN(new_n599));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT102), .B(KEYINPUT11), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT12), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n228), .A2(new_n261), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n261), .A2(new_n225), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT106), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT105), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n606), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT18), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n608), .B1(new_n225), .B2(new_n261), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n610), .B(KEYINPUT13), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT107), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT107), .A3(new_n615), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n605), .B1(new_n613), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n612), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n619), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n604), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n597), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n564), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n515), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(KEYINPUT42), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(G8gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(KEYINPUT42), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(G1325gat));
  NAND2_X1  g436(.A1(new_n560), .A2(new_n595), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(G15gat), .B1(new_n627), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n555), .A2(new_n556), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n642), .B2(G15gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT114), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n627), .A2(new_n359), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  OAI211_X1 g446(.A(new_n359), .B(new_n556), .C1(new_n487), .C2(new_n490), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n492), .B1(new_n648), .B2(new_n592), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n468), .A2(new_n469), .B1(new_n483), .B2(new_n482), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n553), .A2(new_n554), .B1(new_n650), .B2(new_n481), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n651), .A2(KEYINPUT35), .A3(new_n359), .A4(new_n551), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n595), .B(new_n593), .C1(new_n651), .C2(new_n594), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n579), .A2(new_n588), .A3(new_n359), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n649), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n273), .A2(new_n274), .ZN(new_n656));
  INV_X1    g455(.A(new_n626), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n656), .A2(new_n657), .A3(new_n299), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n655), .A2(new_n239), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n221), .A3(new_n564), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n655), .A2(new_n239), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n655), .A2(new_n664), .A3(new_n239), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n564), .A3(new_n658), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n661), .B1(new_n668), .B2(new_n221), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n659), .A2(new_n222), .A3(new_n515), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT115), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT115), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT46), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n666), .A2(new_n515), .A3(new_n658), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(G36gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(KEYINPUT46), .A3(new_n672), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(G1329gat));
  AND3_X1   g478(.A1(new_n655), .A2(new_n664), .A3(new_n239), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n664), .B1(new_n655), .B2(new_n239), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n638), .B(new_n658), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G43gat), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT116), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT47), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(G43gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n659), .A2(new_n686), .A3(new_n641), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n683), .B(new_n687), .C1(new_n684), .C2(KEYINPUT47), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  OAI211_X1 g490(.A(new_n590), .B(new_n658), .C1(new_n680), .C2(new_n681), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G50gat), .ZN(new_n693));
  INV_X1    g492(.A(G50gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n659), .A2(new_n694), .A3(new_n590), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT117), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT48), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT117), .B(new_n699), .C1(new_n693), .C2(new_n695), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(G1331gat));
  AND3_X1   g500(.A1(new_n275), .A2(new_n657), .A3(new_n299), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n655), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n564), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g505(.A(new_n591), .B(new_n703), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1333gat));
  OAI21_X1  g508(.A(G71gat), .B1(new_n703), .B2(new_n639), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n704), .A2(new_n641), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(G71gat), .ZN(new_n712));
  XOR2_X1   g511(.A(new_n712), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g512(.A1(new_n704), .A2(new_n590), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n656), .A2(new_n626), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n299), .B(new_n716), .C1(new_n680), .C2(new_n681), .ZN(new_n717));
  INV_X1    g516(.A(new_n564), .ZN(new_n718));
  OAI21_X1  g517(.A(G85gat), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n653), .A2(new_n654), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n649), .A2(new_n652), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n239), .B(new_n716), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n655), .A2(KEYINPUT51), .A3(new_n239), .A4(new_n716), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(KEYINPUT118), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n725), .A2(KEYINPUT118), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT119), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G85gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n726), .A2(KEYINPUT119), .A3(new_n727), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n299), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n719), .B1(new_n733), .B2(new_n718), .ZN(G1336gat));
  OAI21_X1  g533(.A(G92gat), .B1(new_n717), .B2(new_n591), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n300), .A2(new_n591), .A3(G92gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n239), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n558), .B2(new_n596), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n738), .B2(new_n716), .ZN(new_n739));
  INV_X1    g538(.A(new_n725), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT120), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT120), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(new_n736), .C1(new_n739), .C2(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n735), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT52), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n727), .A3(new_n736), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT121), .A4(new_n736), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n735), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n746), .A2(new_n752), .ZN(G1337gat));
  OAI21_X1  g552(.A(G99gat), .B1(new_n717), .B2(new_n639), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n730), .A2(new_n361), .A3(new_n299), .A4(new_n732), .ZN(new_n755));
  INV_X1    g554(.A(new_n641), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(G1338gat));
  OAI21_X1  g556(.A(G106gat), .B1(new_n717), .B2(new_n359), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n359), .A2(new_n300), .A3(G106gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n739), .B2(new_n740), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT122), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(new_n717), .B2(new_n359), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n300), .B1(new_n663), .B2(new_n665), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(KEYINPUT122), .A3(new_n590), .A4(new_n716), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n766), .A3(G106gat), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  INV_X1    g567(.A(new_n759), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n728), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n762), .B1(new_n767), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n656), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n295), .B2(new_n296), .ZN(new_n774));
  OR2_X1    g573(.A1(new_n287), .A2(new_n288), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT54), .A3(new_n289), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n292), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n776), .A4(new_n292), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n626), .A3(new_n294), .A4(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n614), .A2(new_n615), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n611), .B1(new_n606), .B2(new_n608), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n603), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n299), .A2(new_n625), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n239), .B1(new_n781), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n779), .A2(new_n294), .A3(new_n780), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n239), .A2(new_n625), .A3(new_n785), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n772), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n275), .A2(new_n657), .A3(new_n300), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n718), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n648), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n591), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795), .B2(new_n657), .ZN(new_n796));
  INV_X1    g595(.A(new_n491), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n591), .ZN(new_n799));
  OR2_X1    g598(.A1(new_n799), .A2(G113gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n800), .B2(new_n657), .ZN(G1340gat));
  NOR2_X1   g600(.A1(new_n300), .A2(new_n515), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n426), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G120gat), .B1(new_n795), .B2(new_n300), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1341gat));
  INV_X1    g604(.A(G127gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n795), .A2(new_n806), .A3(new_n772), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n799), .A2(new_n772), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT123), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n806), .ZN(G1342gat));
  NOR3_X1   g609(.A1(new_n799), .A2(G134gat), .A3(new_n737), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT56), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n795), .B2(new_n737), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n639), .A2(new_n564), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n791), .A2(new_n792), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n590), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(G141gat), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n626), .A4(new_n591), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(KEYINPUT57), .A3(new_n590), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n825), .A2(new_n657), .A3(new_n515), .A4(new_n815), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g627(.A(G148gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n829), .A3(new_n802), .ZN(new_n830));
  INV_X1    g629(.A(new_n815), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n824), .A2(new_n831), .A3(new_n299), .A4(new_n591), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n832), .A2(new_n833), .A3(G148gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n657), .B1(new_n301), .B2(new_n302), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n359), .B1(new_n835), .B2(new_n791), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n823), .B1(new_n836), .B2(KEYINPUT57), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n837), .A3(new_n802), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(G148gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n830), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT124), .B(new_n830), .C1(new_n834), .C2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1345gat));
  NAND2_X1  g643(.A1(new_n818), .A2(new_n591), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n772), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n825), .A2(new_n515), .A3(new_n815), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n656), .ZN(new_n848));
  MUX2_X1   g647(.A(new_n846), .B(new_n848), .S(G155gat), .Z(G1346gat));
  NOR2_X1   g648(.A1(new_n845), .A2(new_n737), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n239), .ZN(new_n851));
  MUX2_X1   g650(.A(new_n850), .B(new_n851), .S(G162gat), .Z(G1347gat));
  NOR2_X1   g651(.A1(new_n564), .A2(new_n591), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n816), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n797), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n366), .A3(new_n626), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n794), .ZN(new_n857));
  OAI21_X1  g656(.A(G169gat), .B1(new_n857), .B2(new_n657), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1348gat));
  AOI21_X1  g658(.A(G176gat), .B1(new_n855), .B2(new_n299), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT125), .Z(new_n861));
  INV_X1    g660(.A(new_n372), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n857), .A2(new_n300), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n863), .ZN(G1349gat));
  NAND3_X1  g663(.A1(new_n855), .A2(new_n656), .A3(new_n411), .ZN(new_n865));
  OAI21_X1  g664(.A(G183gat), .B1(new_n857), .B2(new_n772), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g667(.A(G190gat), .B1(new_n857), .B2(new_n737), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT61), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n855), .B(new_n239), .C1(new_n405), .C2(new_n406), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1351gat));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n837), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n639), .A2(new_n853), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n823), .B(KEYINPUT126), .C1(new_n836), .C2(KEYINPUT57), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n874), .A2(new_n626), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G197gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n875), .A2(new_n817), .ZN(new_n880));
  INV_X1    g679(.A(G197gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n626), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n883), .B(new_n884), .ZN(G1352gat));
  NOR4_X1   g684(.A1(new_n875), .A2(G204gat), .A3(new_n300), .A4(new_n817), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT62), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n888));
  OAI21_X1  g687(.A(G204gat), .B1(new_n888), .B2(new_n300), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1353gat));
  NAND3_X1  g689(.A1(new_n880), .A2(new_n656), .A3(new_n324), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n837), .A3(new_n656), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT63), .B1(new_n892), .B2(G211gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(G1354gat));
  OAI21_X1  g695(.A(G218gat), .B1(new_n888), .B2(new_n737), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n325), .A3(new_n239), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1355gat));
endmodule


