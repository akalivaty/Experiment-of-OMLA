//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n545, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n476), .A2(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n478), .B2(G112), .ZN(new_n482));
  NOR3_X1   g057(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n481), .A2(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n464), .A2(G126), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n490), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n479), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n472), .A2(new_n497), .A3(G138), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n493), .A2(new_n494), .B1(new_n496), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT72), .B1(new_n501), .B2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(G543), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n502), .A2(new_n505), .B1(KEYINPUT5), .B2(new_n501), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n507), .A2(new_n508), .B1(G75), .B2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n506), .A2(KEYINPUT74), .A3(G62), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT73), .B(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n514), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AND2_X1   g098(.A1(new_n512), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(G51), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n525), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(new_n524), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OAI221_X1 g106(.A(new_n529), .B1(new_n513), .B2(new_n530), .C1(new_n531), .C2(new_n500), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(new_n506), .A2(G56), .ZN(new_n534));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n500), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n502), .A2(new_n505), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n537), .A2(G81), .A3(new_n538), .A4(new_n512), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n545));
  XOR2_X1   g120(.A(new_n545), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT6), .A2(G651), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT6), .A2(G651), .ZN(new_n552));
  OAI211_X1 g127(.A(G53), .B(G543), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n554));
  OAI211_X1 g129(.A(KEYINPUT77), .B(new_n550), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  INV_X1    g131(.A(new_n553), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(KEYINPUT78), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n553), .B2(KEYINPUT77), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(G78), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n506), .B2(G65), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n500), .B1(new_n513), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n560), .A2(new_n564), .ZN(G299));
  NAND2_X1  g140(.A1(new_n537), .A2(new_n538), .ZN(new_n566));
  INV_X1    g141(.A(G62), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n508), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G75), .A2(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(new_n510), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n514), .A2(new_n515), .B1(G50), .B2(new_n524), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n524), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n506), .A2(G87), .A3(new_n512), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n506), .A2(G86), .A3(new_n512), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n524), .A2(G48), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n500), .ZN(G305));
  AOI22_X1  g156(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n500), .ZN(new_n583));
  INV_X1    g158(.A(G85), .ZN(new_n584));
  INV_X1    g159(.A(G47), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n513), .A2(new_n584), .B1(new_n585), .B2(new_n518), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n583), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT81), .B(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n566), .B2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n518), .A2(KEYINPUT80), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n518), .B2(KEYINPUT80), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n591), .A2(G651), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n537), .A2(G92), .A3(new_n538), .A4(new_n512), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT79), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n506), .A2(new_n599), .A3(G92), .A4(new_n512), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n598), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n588), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n588), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n560), .A2(new_n564), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  XOR2_X1   g184(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g191(.A(new_n477), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G123), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT83), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n472), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n478), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n464), .A2(new_n473), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(G2096), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n624), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NOR2_X1   g223(.A1(G2072), .A2(G2078), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n442), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n648), .B1(new_n651), .B2(KEYINPUT84), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(KEYINPUT84), .B2(new_n651), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n650), .B(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(new_n648), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n648), .A3(new_n654), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT18), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n657), .A3(new_n654), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT85), .Z(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  OR3_X1    g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n683));
  AND3_X1   g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n682), .B1(new_n681), .B2(new_n683), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  NAND2_X1  g262(.A1(new_n472), .A2(G131), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT86), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n617), .A2(G119), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n478), .A2(G107), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G25), .B(new_n693), .S(G29), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT35), .B(G1991), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n694), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G24), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n583), .A2(new_n586), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(G16), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G1971), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n698), .A2(G23), .ZN(new_n708));
  NAND2_X1  g283(.A1(G288), .A2(KEYINPUT88), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n574), .A2(new_n575), .A3(new_n576), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n708), .B1(new_n712), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT33), .B(G1976), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n706), .A2(G1971), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n707), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G305), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT32), .B(G1981), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n713), .B2(new_n714), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n717), .B2(new_n723), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n704), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n730));
  AOI21_X1  g305(.A(KEYINPUT91), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(KEYINPUT90), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT36), .B1(new_n729), .B2(KEYINPUT90), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n729), .A2(KEYINPUT90), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n736), .A2(new_n732), .A3(KEYINPUT91), .A4(KEYINPUT36), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n623), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(KEYINPUT97), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G11), .Z(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT98), .B(G28), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT99), .Z(new_n744));
  AOI211_X1 g319(.A(G29), .B(new_n744), .C1(KEYINPUT30), .C2(new_n742), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n740), .A2(new_n741), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2084), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G34), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(new_n738), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(new_n738), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n739), .A2(KEYINPUT97), .B1(new_n747), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n738), .A2(G35), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT100), .Z(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n738), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT29), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n746), .B(new_n753), .C1(G2090), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n738), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n738), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n698), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n698), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n738), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n617), .A2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n472), .A2(G140), .ZN(new_n769));
  OR2_X1    g344(.A1(G104), .A2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n770), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n738), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n738), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n617), .A2(G129), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n473), .A2(G105), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(G141), .C2(new_n472), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n765), .B(new_n776), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n758), .A2(new_n761), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n698), .A2(G5), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G171), .B2(new_n698), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1961), .ZN(new_n792));
  NOR2_X1   g367(.A1(G16), .A2(G19), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n542), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT92), .B(G1341), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  NAND4_X1  g371(.A1(new_n788), .A2(new_n791), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n785), .A2(new_n786), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n738), .A2(G33), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT25), .Z(new_n803));
  INV_X1    g378(.A(G139), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n479), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n464), .A2(G127), .ZN(new_n806));
  NAND2_X1  g381(.A1(G115), .A2(G2104), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n478), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n801), .B1(new_n809), .B2(new_n738), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G2072), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(G2072), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n752), .A2(new_n747), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n800), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT96), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n604), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G4), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n815), .B1(G1348), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n698), .A2(G20), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT23), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n608), .B2(new_n698), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G1956), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n757), .A2(G2090), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT101), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n818), .A2(G1348), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n814), .B2(KEYINPUT96), .ZN(new_n828));
  NOR4_X1   g403(.A1(new_n797), .A2(new_n819), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n735), .A2(new_n737), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(new_n604), .A2(G559), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n537), .A2(G56), .A3(new_n538), .ZN(new_n835));
  INV_X1    g410(.A(new_n535), .ZN(new_n836));
  OAI21_X1  g411(.A(G651), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n537), .A2(G67), .A3(new_n538), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  INV_X1    g416(.A(new_n541), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n537), .A2(G93), .A3(new_n538), .A4(new_n512), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n512), .A2(G55), .A3(G543), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n837), .A2(new_n841), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n500), .B1(new_n838), .B2(new_n839), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n844), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n536), .A2(new_n541), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n834), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n784), .B(new_n772), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n491), .B1(new_n496), .B2(new_n498), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n784), .B(new_n773), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n496), .A2(new_n498), .ZN(new_n863));
  INV_X1    g438(.A(new_n491), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n861), .A2(new_n866), .B1(new_n808), .B2(new_n805), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n859), .A2(new_n860), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n869), .A3(new_n809), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n693), .B(new_n626), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n472), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n478), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n873), .B1(new_n874), .B2(new_n875), .C1(new_n876), .C2(new_n477), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT104), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n867), .A2(new_n878), .A3(new_n870), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G160), .B(G162), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT103), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n623), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n867), .A2(KEYINPUT104), .A3(new_n878), .A4(new_n870), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n871), .B2(new_n879), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n888), .B2(new_n881), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g466(.A1(new_n603), .A2(G299), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n597), .A2(new_n600), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT10), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n608), .A3(new_n595), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n892), .A2(new_n897), .A3(KEYINPUT41), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n892), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n604), .A2(new_n611), .A3(new_n850), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n613), .A2(new_n851), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n897), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n700), .A2(new_n709), .A3(new_n711), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n700), .B1(new_n709), .B2(new_n711), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT105), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n712), .A2(G290), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n907), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n511), .A2(new_n519), .A3(G305), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n719), .B1(new_n571), .B2(new_n572), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G303), .A2(G305), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n719), .A2(new_n571), .A3(new_n572), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(new_n912), .A3(new_n911), .A4(new_n907), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n906), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n923), .B(new_n922), .C1(new_n903), .C2(new_n905), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G868), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n927), .A3(new_n926), .A4(new_n928), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n847), .B2(new_n848), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n931), .B2(new_n932), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n934), .A2(new_n937), .ZN(G295));
  NOR2_X1   g513(.A1(new_n934), .A2(new_n937), .ZN(G331));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n846), .A2(G301), .A3(new_n849), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n846), .B2(new_n849), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n941), .A2(new_n942), .A3(G286), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n850), .A2(G171), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n846), .A2(G301), .A3(new_n849), .ZN(new_n945));
  AOI21_X1  g520(.A(G168), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n900), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n603), .A2(G299), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n608), .B1(new_n896), .B2(new_n595), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n892), .A2(new_n897), .A3(KEYINPUT41), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(G168), .A3(new_n945), .ZN(new_n955));
  OAI21_X1  g530(.A(G286), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT109), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n904), .B1(new_n956), .B2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n922), .ZN(new_n962));
  INV_X1    g537(.A(G37), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n917), .A2(new_n921), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n949), .A2(new_n958), .A3(new_n964), .A4(new_n960), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n957), .B1(new_n959), .B2(KEYINPUT110), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  AOI211_X1 g544(.A(new_n969), .B(new_n904), .C1(new_n956), .C2(new_n955), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n922), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n971), .A2(new_n963), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT43), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n940), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n971), .A2(new_n965), .A3(new_n963), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n962), .A2(new_n973), .A3(new_n963), .A4(new_n965), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n978), .A2(KEYINPUT44), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT111), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT44), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n966), .A2(KEYINPUT43), .B1(new_n972), .B2(new_n974), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n940), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n865), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n988), .A2(KEYINPUT112), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n467), .A2(G40), .A3(new_n474), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n988), .B2(KEYINPUT112), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n772), .B(G2067), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n784), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n997), .B1(new_n996), .B2(new_n999), .ZN(new_n1001));
  INV_X1    g576(.A(new_n784), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1002), .B2(new_n994), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n992), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n992), .A2(new_n994), .A3(new_n1002), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(KEYINPUT113), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n693), .A2(new_n696), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n693), .A2(new_n696), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n993), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n700), .A2(new_n702), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n992), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1000), .A2(new_n1001), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1008), .A2(new_n1009), .B1(new_n775), .B2(new_n773), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT126), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n992), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT71), .B1(new_n488), .B2(new_n490), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n490), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n863), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n987), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n467), .A2(G40), .A3(new_n474), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n863), .B2(new_n864), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1961), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n860), .B2(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2078), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1035), .A2(new_n990), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1036), .B1(G164), .B2(G1384), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1038), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G171), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n989), .A2(new_n991), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1028), .A2(KEYINPUT124), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1039), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1028), .B2(KEYINPUT124), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1049), .A2(new_n1054), .B1(new_n1045), .B2(new_n1038), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1961), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1048), .B1(new_n1060), .B2(G171), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G303), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1971), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1067), .A2(KEYINPUT114), .B1(new_n1032), .B2(G2090), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(G1971), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1066), .B(G8), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1028), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n1072));
  INV_X1    g647(.A(G2090), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1025), .A2(new_n1030), .A3(new_n987), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1075), .B2(new_n1067), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1064), .B(KEYINPUT55), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1029), .B2(new_n990), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n712), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT52), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n1084));
  AND2_X1   g659(.A1(G305), .A2(G1981), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G305), .A2(G1981), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n580), .A2(new_n500), .ZN(new_n1088));
  INV_X1    g663(.A(G1981), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n578), .A4(new_n579), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1080), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1080), .B(new_n1094), .C1(new_n712), .C2(new_n1081), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1083), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1071), .A2(new_n1078), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1062), .B1(new_n1099), .B2(G301), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1060), .A2(G171), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(G164), .A2(new_n1036), .A3(G1384), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1037), .A2(new_n990), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n764), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1027), .A2(new_n747), .A3(new_n1031), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(G168), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G8), .ZN(new_n1108));
  AOI21_X1  g683(.A(G168), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1111), .A3(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1063), .A2(new_n1098), .A3(new_n1102), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1029), .A2(new_n990), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT120), .B1(new_n1115), .B2(G2067), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1029), .A2(new_n990), .A3(new_n1117), .A4(new_n775), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1348), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n604), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n604), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT60), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(G1956), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1042), .A2(new_n1043), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT119), .B1(G299), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n608), .A2(new_n1131), .A3(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n560), .B2(new_n564), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1133), .B(new_n1136), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(KEYINPUT61), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1124), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1042), .A2(new_n1043), .A3(new_n994), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT121), .A4(new_n994), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT58), .B(G1341), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1115), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1142), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1149), .ZN(new_n1151));
  AOI211_X1 g726(.A(KEYINPUT122), .B(new_n1151), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n542), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(KEYINPUT59), .B(new_n542), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1157));
  NOR4_X1   g732(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT60), .A4(new_n603), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1141), .A2(new_n1155), .A3(new_n1156), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1139), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1122), .B2(new_n1138), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1114), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G288), .A2(G1976), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1086), .B1(new_n1093), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1080), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g742(.A(KEYINPUT115), .B(new_n1086), .C1(new_n1093), .C2(new_n1164), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1083), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1167), .A2(new_n1168), .B1(new_n1071), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1067), .A2(KEYINPUT114), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1070), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1032), .A2(G2090), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1176), .A2(new_n1096), .A3(G8), .A4(new_n1066), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1177), .B(KEYINPUT116), .C1(new_n1168), .C2(new_n1167), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1040), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1056), .ZN(new_n1181));
  AOI21_X1  g756(.A(G301), .B1(new_n1181), .B2(new_n1046), .ZN(new_n1182));
  AND4_X1   g757(.A1(new_n1071), .A2(new_n1078), .A3(new_n1182), .A4(new_n1096), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1110), .A2(new_n1184), .A3(new_n1112), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1184), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1183), .B(new_n1185), .C1(new_n1186), .C2(KEYINPUT125), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1186), .A2(KEYINPUT125), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1179), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1079), .B(G286), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1071), .A2(KEYINPUT63), .A3(new_n1096), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1066), .B1(new_n1176), .B2(G8), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AND4_X1   g768(.A1(new_n1071), .A2(new_n1078), .A3(new_n1096), .A4(new_n1190), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n1194), .B2(KEYINPUT117), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT117), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1190), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1196), .B1(new_n1097), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1193), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1163), .A2(new_n1189), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(G290), .A2(G1986), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n992), .B1(new_n1013), .B2(new_n1201), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1012), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1022), .B1(new_n1200), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g779(.A(new_n984), .ZN(new_n1206));
  NOR3_X1   g780(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1207));
  AND4_X1   g781(.A1(new_n686), .A2(new_n1206), .A3(new_n890), .A4(new_n1207), .ZN(G308));
  NAND4_X1  g782(.A1(new_n686), .A2(new_n1206), .A3(new_n890), .A4(new_n1207), .ZN(G225));
endmodule


