

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740;

  XNOR2_X1 U371 ( .A(n541), .B(n540), .ZN(n552) );
  XNOR2_X1 U372 ( .A(n445), .B(n718), .ZN(n460) );
  XOR2_X1 U373 ( .A(n379), .B(n378), .Z(n350) );
  XNOR2_X2 U374 ( .A(n367), .B(n543), .ZN(n681) );
  OR2_X2 U375 ( .A1(n539), .A2(n662), .ZN(n541) );
  XNOR2_X2 U376 ( .A(n512), .B(KEYINPUT1), .ZN(n539) );
  XNOR2_X1 U377 ( .A(KEYINPUT82), .B(G104), .ZN(n442) );
  INV_X1 U378 ( .A(G953), .ZN(n736) );
  NOR2_X1 U379 ( .A1(G237), .A2(G953), .ZN(n377) );
  XNOR2_X1 U380 ( .A(n442), .B(G110), .ZN(n468) );
  OR2_X1 U381 ( .A1(n688), .A2(n575), .ZN(n516) );
  XNOR2_X1 U382 ( .A(n498), .B(KEYINPUT22), .ZN(n535) );
  INV_X1 U383 ( .A(n351), .ZN(n485) );
  OR2_X1 U384 ( .A1(n499), .A2(n495), .ZN(n662) );
  OR2_X1 U385 ( .A1(n699), .A2(G902), .ZN(n452) );
  XNOR2_X1 U386 ( .A(n731), .B(G146), .ZN(n450) );
  XNOR2_X1 U387 ( .A(n471), .B(n470), .ZN(n720) );
  XNOR2_X1 U388 ( .A(n419), .B(n374), .ZN(n731) );
  XNOR2_X1 U389 ( .A(G137), .B(G140), .ZN(n441) );
  XNOR2_X1 U390 ( .A(n352), .B(n475), .ZN(n351) );
  NOR2_X1 U391 ( .A1(n631), .A2(n604), .ZN(n352) );
  BUF_X1 U392 ( .A(n551), .Z(n353) );
  XNOR2_X1 U393 ( .A(n358), .B(n359), .ZN(n551) );
  BUF_X1 U394 ( .A(n596), .Z(n354) );
  XNOR2_X1 U395 ( .A(n613), .B(KEYINPUT71), .ZN(n355) );
  XNOR2_X1 U396 ( .A(n613), .B(KEYINPUT71), .ZN(n607) );
  INV_X1 U397 ( .A(n524), .ZN(n356) );
  INV_X1 U398 ( .A(n503), .ZN(n357) );
  NOR2_X1 U399 ( .A1(n616), .A2(G902), .ZN(n358) );
  XOR2_X1 U400 ( .A(G472), .B(KEYINPUT96), .Z(n359) );
  NAND2_X2 U401 ( .A1(n601), .A2(n600), .ZN(n613) );
  XNOR2_X1 U402 ( .A(n486), .B(KEYINPUT79), .ZN(n522) );
  NAND2_X1 U403 ( .A1(n552), .A2(n500), .ZN(n367) );
  NAND2_X1 U404 ( .A1(n523), .A2(n522), .ZN(n366) );
  XNOR2_X1 U405 ( .A(n521), .B(n520), .ZN(n523) );
  INV_X1 U406 ( .A(KEYINPUT110), .ZN(n520) );
  INV_X1 U407 ( .A(KEYINPUT104), .ZN(n370) );
  XNOR2_X1 U408 ( .A(n397), .B(G128), .ZN(n398) );
  XNOR2_X1 U409 ( .A(G119), .B(KEYINPUT90), .ZN(n397) );
  OR2_X1 U410 ( .A1(n542), .A2(n508), .ZN(n418) );
  AND2_X1 U411 ( .A1(n620), .A2(G953), .ZN(n712) );
  XNOR2_X1 U412 ( .A(n364), .B(n525), .ZN(n591) );
  NAND2_X1 U413 ( .A1(n365), .A2(n524), .ZN(n364) );
  XNOR2_X1 U414 ( .A(n366), .B(n363), .ZN(n365) );
  INV_X1 U415 ( .A(KEYINPUT34), .ZN(n544) );
  NAND2_X1 U416 ( .A1(n518), .A2(n369), .ZN(n519) );
  AND2_X1 U417 ( .A1(n480), .A2(n479), .ZN(n360) );
  XOR2_X1 U418 ( .A(n511), .B(KEYINPUT28), .Z(n361) );
  NAND2_X1 U419 ( .A1(n473), .A2(G214), .ZN(n362) );
  XOR2_X1 U420 ( .A(KEYINPUT78), .B(KEYINPUT36), .Z(n363) );
  XNOR2_X1 U421 ( .A(n353), .B(KEYINPUT6), .ZN(n542) );
  XNOR2_X2 U422 ( .A(KEYINPUT65), .B(G101), .ZN(n445) );
  XNOR2_X1 U423 ( .A(n368), .B(n450), .ZN(n616) );
  XNOR2_X1 U424 ( .A(n350), .B(n380), .ZN(n368) );
  INV_X1 U425 ( .A(n510), .ZN(n369) );
  XNOR2_X2 U426 ( .A(n558), .B(n370), .ZN(n510) );
  BUF_X1 U427 ( .A(n696), .Z(n707) );
  OR2_X1 U428 ( .A1(KEYINPUT44), .A2(KEYINPUT67), .ZN(n371) );
  OR2_X1 U429 ( .A1(n490), .A2(n489), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n550), .B(n371), .ZN(n569) );
  NAND2_X1 U431 ( .A1(n351), .A2(n362), .ZN(n486) );
  INV_X1 U432 ( .A(KEYINPUT30), .ZN(n477) );
  XNOR2_X2 U433 ( .A(G143), .B(G128), .ZN(n463) );
  INV_X1 U434 ( .A(G134), .ZN(n373) );
  XNOR2_X2 U435 ( .A(n463), .B(n373), .ZN(n419) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(G131), .ZN(n374) );
  XNOR2_X2 U437 ( .A(KEYINPUT3), .B(G119), .ZN(n718) );
  XNOR2_X1 U438 ( .A(G113), .B(G116), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n375), .B(KEYINPUT95), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n460), .B(n376), .ZN(n380) );
  XNOR2_X1 U441 ( .A(KEYINPUT72), .B(n377), .ZN(n433) );
  NAND2_X1 U442 ( .A1(n433), .A2(G210), .ZN(n379) );
  XNOR2_X1 U443 ( .A(KEYINPUT5), .B(G137), .ZN(n378) );
  XOR2_X1 U444 ( .A(KEYINPUT14), .B(KEYINPUT85), .Z(n382) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n387) );
  NAND2_X1 U447 ( .A1(n387), .A2(G902), .ZN(n383) );
  XOR2_X1 U448 ( .A(KEYINPUT87), .B(n383), .Z(n488) );
  OR2_X1 U449 ( .A1(n736), .A2(n488), .ZN(n384) );
  NOR2_X1 U450 ( .A1(G900), .A2(n384), .ZN(n386) );
  INV_X1 U451 ( .A(KEYINPUT106), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n389) );
  NAND2_X1 U453 ( .A1(G952), .A2(n387), .ZN(n687) );
  NOR2_X1 U454 ( .A1(n687), .A2(G953), .ZN(n489) );
  INV_X1 U455 ( .A(n489), .ZN(n388) );
  NAND2_X1 U456 ( .A1(n389), .A2(n388), .ZN(n479) );
  INV_X1 U457 ( .A(KEYINPUT15), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n390), .B(G902), .ZN(n604) );
  INV_X1 U459 ( .A(n604), .ZN(n606) );
  NAND2_X1 U460 ( .A1(n606), .A2(G234), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n391), .B(KEYINPUT20), .ZN(n410) );
  INV_X1 U462 ( .A(n410), .ZN(n393) );
  INV_X1 U463 ( .A(G221), .ZN(n392) );
  OR2_X1 U464 ( .A1(n393), .A2(n392), .ZN(n396) );
  INV_X1 U465 ( .A(KEYINPUT93), .ZN(n394) );
  XNOR2_X1 U466 ( .A(n394), .B(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n396), .B(n395), .ZN(n495) );
  INV_X1 U468 ( .A(n495), .ZN(n658) );
  AND2_X1 U469 ( .A1(n479), .A2(n658), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n398), .B(n441), .ZN(n402) );
  XOR2_X1 U471 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n400) );
  NAND2_X1 U472 ( .A1(G234), .A2(n736), .ZN(n399) );
  XNOR2_X1 U473 ( .A(n400), .B(n399), .ZN(n422) );
  NAND2_X1 U474 ( .A1(n422), .A2(G221), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n409) );
  XNOR2_X1 U476 ( .A(G146), .B(G125), .ZN(n458) );
  INV_X1 U477 ( .A(KEYINPUT10), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n458), .B(n403), .ZN(n728) );
  INV_X1 U479 ( .A(n728), .ZN(n407) );
  XNOR2_X1 U480 ( .A(G110), .B(KEYINPUT23), .ZN(n405) );
  XNOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n404) );
  XNOR2_X1 U482 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U483 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U484 ( .A(n409), .B(n408), .ZN(n708) );
  INV_X1 U485 ( .A(G902), .ZN(n454) );
  NAND2_X1 U486 ( .A1(n708), .A2(n454), .ZN(n416) );
  AND2_X1 U487 ( .A1(n410), .A2(G217), .ZN(n414) );
  XNOR2_X1 U488 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n412) );
  XNOR2_X1 U489 ( .A(KEYINPUT25), .B(KEYINPUT74), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U491 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U492 ( .A(n416), .B(n415), .ZN(n499) );
  NAND2_X1 U493 ( .A1(n417), .A2(n499), .ZN(n508) );
  XNOR2_X1 U494 ( .A(n418), .B(KEYINPUT107), .ZN(n440) );
  XNOR2_X1 U495 ( .A(KEYINPUT97), .B(KEYINPUT7), .ZN(n426) );
  XNOR2_X1 U496 ( .A(G116), .B(G107), .ZN(n467) );
  XOR2_X1 U497 ( .A(G122), .B(KEYINPUT9), .Z(n420) );
  XNOR2_X1 U498 ( .A(n467), .B(n420), .ZN(n421) );
  XNOR2_X1 U499 ( .A(n419), .B(n421), .ZN(n424) );
  NAND2_X1 U500 ( .A1(G217), .A2(n422), .ZN(n423) );
  XOR2_X1 U501 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U502 ( .A(n426), .B(n425), .ZN(n703) );
  NOR2_X1 U503 ( .A1(G902), .A2(n703), .ZN(n428) );
  XOR2_X1 U504 ( .A(KEYINPUT98), .B(G478), .Z(n427) );
  XNOR2_X1 U505 ( .A(n428), .B(n427), .ZN(n561) );
  XNOR2_X1 U506 ( .A(G113), .B(G122), .ZN(n469) );
  XNOR2_X1 U507 ( .A(G143), .B(G131), .ZN(n429) );
  XNOR2_X1 U508 ( .A(n469), .B(n429), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n728), .B(n430), .ZN(n437) );
  XOR2_X1 U510 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n432) );
  XNOR2_X1 U511 ( .A(G140), .B(G104), .ZN(n431) );
  XNOR2_X1 U512 ( .A(n432), .B(n431), .ZN(n435) );
  NAND2_X1 U513 ( .A1(n433), .A2(G214), .ZN(n434) );
  XNOR2_X1 U514 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U515 ( .A(n437), .B(n436), .ZN(n625) );
  NAND2_X1 U516 ( .A1(n625), .A2(n454), .ZN(n439) );
  XNOR2_X1 U517 ( .A(KEYINPUT13), .B(G475), .ZN(n438) );
  XNOR2_X1 U518 ( .A(n439), .B(n438), .ZN(n560) );
  OR2_X1 U519 ( .A1(n561), .A2(n560), .ZN(n650) );
  INV_X1 U520 ( .A(n650), .ZN(n647) );
  NAND2_X1 U521 ( .A1(n440), .A2(n647), .ZN(n521) );
  XNOR2_X1 U522 ( .A(n441), .B(KEYINPUT88), .ZN(n729) );
  XNOR2_X1 U523 ( .A(n729), .B(n468), .ZN(n448) );
  XNOR2_X1 U524 ( .A(G107), .B(KEYINPUT75), .ZN(n444) );
  NAND2_X1 U525 ( .A1(n736), .A2(G227), .ZN(n443) );
  XNOR2_X1 U526 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U527 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U528 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n450), .B(n449), .ZN(n699) );
  INV_X1 U530 ( .A(G469), .ZN(n451) );
  XNOR2_X2 U531 ( .A(n452), .B(n451), .ZN(n512) );
  INV_X1 U532 ( .A(n539), .ZN(n524) );
  INV_X1 U533 ( .A(G237), .ZN(n453) );
  NAND2_X1 U534 ( .A1(n454), .A2(n453), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n356), .A2(n362), .ZN(n455) );
  OR2_X1 U536 ( .A1(n521), .A2(n455), .ZN(n456) );
  XNOR2_X1 U537 ( .A(n456), .B(KEYINPUT43), .ZN(n476) );
  XNOR2_X1 U538 ( .A(KEYINPUT83), .B(KEYINPUT4), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U540 ( .A(n460), .B(n459), .ZN(n466) );
  XNOR2_X1 U541 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n462) );
  NAND2_X1 U542 ( .A1(n736), .A2(G224), .ZN(n461) );
  XNOR2_X1 U543 ( .A(n462), .B(n461), .ZN(n464) );
  XNOR2_X1 U544 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U545 ( .A(n466), .B(n465), .ZN(n472) );
  XNOR2_X1 U546 ( .A(n468), .B(n467), .ZN(n471) );
  XNOR2_X1 U547 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U548 ( .A(n472), .B(n720), .ZN(n631) );
  NAND2_X1 U549 ( .A1(n473), .A2(G210), .ZN(n474) );
  XNOR2_X1 U550 ( .A(n474), .B(KEYINPUT84), .ZN(n475) );
  NAND2_X1 U551 ( .A1(n476), .A2(n485), .ZN(n599) );
  XNOR2_X1 U552 ( .A(n599), .B(G140), .ZN(G42) );
  INV_X1 U553 ( .A(n551), .ZN(n558) );
  NAND2_X1 U554 ( .A1(n510), .A2(n362), .ZN(n478) );
  XNOR2_X1 U555 ( .A(n478), .B(n477), .ZN(n481) );
  OR2_X1 U556 ( .A1(n662), .A2(n512), .ZN(n554) );
  INV_X1 U557 ( .A(n554), .ZN(n480) );
  NAND2_X1 U558 ( .A1(n481), .A2(n360), .ZN(n482) );
  XNOR2_X1 U559 ( .A(n482), .B(KEYINPUT73), .ZN(n527) );
  INV_X1 U560 ( .A(n561), .ZN(n483) );
  OR2_X1 U561 ( .A1(n483), .A2(n560), .ZN(n546) );
  NOR2_X1 U562 ( .A1(n546), .A2(n485), .ZN(n484) );
  AND2_X1 U563 ( .A1(n527), .A2(n484), .ZN(n574) );
  XOR2_X1 U564 ( .A(G143), .B(n574), .Z(G45) );
  XNOR2_X1 U565 ( .A(n522), .B(KEYINPUT19), .ZN(n487) );
  INV_X1 U566 ( .A(n487), .ZN(n577) );
  XOR2_X1 U567 ( .A(G898), .B(KEYINPUT86), .Z(n715) );
  NAND2_X1 U568 ( .A1(G953), .A2(n715), .ZN(n722) );
  NOR2_X1 U569 ( .A1(n488), .A2(n722), .ZN(n490) );
  NAND2_X1 U570 ( .A1(n577), .A2(n372), .ZN(n492) );
  XNOR2_X1 U571 ( .A(KEYINPUT64), .B(KEYINPUT0), .ZN(n491) );
  XNOR2_X1 U572 ( .A(n492), .B(n491), .ZN(n555) );
  INV_X1 U573 ( .A(n560), .ZN(n493) );
  OR2_X1 U574 ( .A1(n561), .A2(n493), .ZN(n494) );
  XNOR2_X1 U575 ( .A(n494), .B(KEYINPUT100), .ZN(n677) );
  NOR2_X1 U576 ( .A1(n677), .A2(n495), .ZN(n496) );
  XNOR2_X1 U577 ( .A(n496), .B(KEYINPUT101), .ZN(n497) );
  OR2_X2 U578 ( .A1(n555), .A2(n497), .ZN(n498) );
  INV_X1 U579 ( .A(n535), .ZN(n503) );
  INV_X1 U580 ( .A(n499), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(KEYINPUT102), .ZN(n659) );
  NAND2_X1 U582 ( .A1(n356), .A2(n659), .ZN(n501) );
  INV_X1 U583 ( .A(n542), .ZN(n500) );
  NOR2_X1 U584 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U585 ( .A1(n503), .A2(n502), .ZN(n563) );
  XNOR2_X1 U586 ( .A(n563), .B(G101), .ZN(G3) );
  INV_X1 U587 ( .A(n677), .ZN(n504) );
  AND2_X1 U588 ( .A1(n504), .A2(n362), .ZN(n505) );
  XNOR2_X1 U589 ( .A(n485), .B(KEYINPUT38), .ZN(n675) );
  NAND2_X1 U590 ( .A1(n505), .A2(n675), .ZN(n507) );
  INV_X1 U591 ( .A(KEYINPUT41), .ZN(n506) );
  XNOR2_X1 U592 ( .A(n507), .B(n506), .ZN(n688) );
  INV_X1 U593 ( .A(n508), .ZN(n509) );
  NAND2_X1 U594 ( .A1(n510), .A2(n509), .ZN(n511) );
  INV_X1 U595 ( .A(n512), .ZN(n513) );
  NAND2_X1 U596 ( .A1(n361), .A2(n513), .ZN(n514) );
  XNOR2_X1 U597 ( .A(n514), .B(KEYINPUT108), .ZN(n575) );
  XNOR2_X1 U598 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n515) );
  XNOR2_X1 U599 ( .A(n516), .B(n515), .ZN(n571) );
  XOR2_X1 U600 ( .A(G137), .B(n571), .Z(G39) );
  NOR2_X1 U601 ( .A1(n524), .A2(n517), .ZN(n518) );
  NOR2_X1 U602 ( .A1(n357), .A2(n519), .ZN(n537) );
  XOR2_X1 U603 ( .A(G110), .B(n537), .Z(G12) );
  INV_X1 U604 ( .A(KEYINPUT111), .ZN(n525) );
  XOR2_X1 U605 ( .A(G125), .B(KEYINPUT37), .Z(n526) );
  XNOR2_X1 U606 ( .A(n591), .B(n526), .ZN(G27) );
  NAND2_X1 U607 ( .A1(n527), .A2(n675), .ZN(n529) );
  XNOR2_X1 U608 ( .A(KEYINPUT68), .B(KEYINPUT39), .ZN(n528) );
  XNOR2_X2 U609 ( .A(n529), .B(n528), .ZN(n596) );
  NAND2_X1 U610 ( .A1(n596), .A2(n647), .ZN(n531) );
  INV_X1 U611 ( .A(KEYINPUT40), .ZN(n530) );
  XNOR2_X1 U612 ( .A(n531), .B(n530), .ZN(n572) );
  BUF_X1 U613 ( .A(n572), .Z(n532) );
  XOR2_X1 U614 ( .A(G131), .B(n532), .Z(G33) );
  NOR2_X1 U615 ( .A1(n539), .A2(n659), .ZN(n533) );
  NAND2_X1 U616 ( .A1(n533), .A2(n542), .ZN(n534) );
  NOR2_X1 U617 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U618 ( .A(n536), .B(KEYINPUT32), .ZN(n538) );
  XOR2_X1 U619 ( .A(n538), .B(G119), .Z(G21) );
  NOR2_X1 U620 ( .A1(n538), .A2(n537), .ZN(n549) );
  INV_X1 U621 ( .A(KEYINPUT70), .ZN(n540) );
  XNOR2_X1 U622 ( .A(KEYINPUT105), .B(KEYINPUT33), .ZN(n543) );
  NOR2_X1 U623 ( .A1(n681), .A2(n555), .ZN(n545) );
  XNOR2_X1 U624 ( .A(n545), .B(n544), .ZN(n547) );
  NOR2_X1 U625 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U626 ( .A(n548), .B(KEYINPUT35), .ZN(n637) );
  NAND2_X1 U627 ( .A1(n549), .A2(n637), .ZN(n550) );
  NAND2_X1 U628 ( .A1(n552), .A2(n353), .ZN(n667) );
  NOR2_X1 U629 ( .A1(n555), .A2(n667), .ZN(n553) );
  XNOR2_X1 U630 ( .A(n553), .B(KEYINPUT31), .ZN(n652) );
  OR2_X1 U631 ( .A1(n555), .A2(n554), .ZN(n557) );
  INV_X1 U632 ( .A(KEYINPUT94), .ZN(n556) );
  XNOR2_X1 U633 ( .A(n557), .B(n556), .ZN(n559) );
  NAND2_X1 U634 ( .A1(n559), .A2(n558), .ZN(n640) );
  NAND2_X1 U635 ( .A1(n652), .A2(n640), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n561), .A2(n560), .ZN(n653) );
  XNOR2_X1 U637 ( .A(n653), .B(KEYINPUT99), .ZN(n597) );
  OR2_X1 U638 ( .A1(n597), .A2(n647), .ZN(n672) );
  NAND2_X1 U639 ( .A1(n562), .A2(n672), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U641 ( .A(n565), .B(KEYINPUT103), .ZN(n567) );
  NAND2_X1 U642 ( .A1(KEYINPUT44), .A2(KEYINPUT67), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X2 U644 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X2 U645 ( .A(n570), .B(KEYINPUT45), .ZN(n612) );
  NOR2_X2 U646 ( .A1(n612), .A2(KEYINPUT77), .ZN(n602) );
  NOR2_X2 U647 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n573), .B(KEYINPUT46), .ZN(n593) );
  XNOR2_X1 U649 ( .A(n574), .B(KEYINPUT76), .ZN(n589) );
  INV_X1 U650 ( .A(n575), .ZN(n576) );
  AND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n648) );
  INV_X1 U652 ( .A(KEYINPUT69), .ZN(n578) );
  AND2_X1 U653 ( .A1(n672), .A2(n578), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n648), .A2(n579), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n580), .A2(KEYINPUT47), .ZN(n587) );
  INV_X1 U656 ( .A(n672), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n581), .A2(KEYINPUT69), .ZN(n584) );
  NOR2_X1 U658 ( .A1(KEYINPUT69), .A2(KEYINPUT47), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n672), .A2(n582), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n648), .A2(n585), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  AND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n595) );
  INV_X1 U666 ( .A(KEYINPUT48), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n595), .B(n594), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n354), .A2(n597), .ZN(n598) );
  XNOR2_X1 U669 ( .A(n598), .B(KEYINPUT112), .ZN(n740) );
  AND2_X1 U670 ( .A1(n740), .A2(n599), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n607), .A2(n602), .ZN(n603) );
  INV_X1 U672 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U673 ( .A1(n603), .A2(n656), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n612), .A2(n606), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n608), .A2(n355), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n609), .A2(KEYINPUT77), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n612), .A2(n613), .ZN(n657) );
  NAND2_X1 U680 ( .A1(n657), .A2(KEYINPUT2), .ZN(n614) );
  AND2_X2 U681 ( .A1(n615), .A2(n614), .ZN(n696) );
  NAND2_X1 U682 ( .A1(n696), .A2(G472), .ZN(n619) );
  XNOR2_X1 U683 ( .A(KEYINPUT80), .B(KEYINPUT62), .ZN(n617) );
  XNOR2_X1 U684 ( .A(n616), .B(n617), .ZN(n618) );
  XNOR2_X1 U685 ( .A(n619), .B(n618), .ZN(n621) );
  INV_X1 U686 ( .A(G952), .ZN(n620) );
  NOR2_X2 U687 ( .A1(n621), .A2(n712), .ZN(n623) );
  XNOR2_X1 U688 ( .A(KEYINPUT113), .B(KEYINPUT63), .ZN(n622) );
  XNOR2_X1 U689 ( .A(n623), .B(n622), .ZN(G57) );
  NAND2_X1 U690 ( .A1(n696), .A2(G475), .ZN(n627) );
  XOR2_X1 U691 ( .A(KEYINPUT81), .B(KEYINPUT59), .Z(n624) );
  XNOR2_X1 U692 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U693 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U694 ( .A1(n628), .A2(n712), .ZN(n630) );
  XOR2_X1 U695 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n629) );
  XNOR2_X1 U696 ( .A(n630), .B(n629), .ZN(G60) );
  NAND2_X1 U697 ( .A1(n696), .A2(G210), .ZN(n634) );
  XOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n632) );
  XNOR2_X1 U699 ( .A(n631), .B(n632), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X2 U701 ( .A1(n635), .A2(n712), .ZN(n636) );
  XNOR2_X1 U702 ( .A(n636), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U703 ( .A(n637), .B(G122), .ZN(G24) );
  NOR2_X1 U704 ( .A1(n640), .A2(n650), .ZN(n638) );
  XOR2_X1 U705 ( .A(KEYINPUT114), .B(n638), .Z(n639) );
  XNOR2_X1 U706 ( .A(G104), .B(n639), .ZN(G6) );
  NOR2_X1 U707 ( .A1(n640), .A2(n653), .ZN(n642) );
  XNOR2_X1 U708 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U710 ( .A(G107), .B(n643), .ZN(G9) );
  XOR2_X1 U711 ( .A(G128), .B(KEYINPUT29), .Z(n646) );
  INV_X1 U712 ( .A(n653), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n648), .A2(n644), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(G30) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(G146), .B(n649), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n650), .A2(n652), .ZN(n651) );
  XOR2_X1 U718 ( .A(G113), .B(n651), .Z(G15) );
  NOR2_X1 U719 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U720 ( .A(G116), .B(KEYINPUT115), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(G18) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(n693) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(n660), .Z(n661) );
  NOR2_X1 U725 ( .A1(n661), .A2(n353), .ZN(n666) );
  NAND2_X1 U726 ( .A1(n356), .A2(n662), .ZN(n664) );
  XNOR2_X1 U727 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n668) );
  AND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U731 ( .A(n669), .B(KEYINPUT117), .ZN(n670) );
  XNOR2_X1 U732 ( .A(KEYINPUT51), .B(n670), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n671), .A2(n688), .ZN(n684) );
  NAND2_X1 U734 ( .A1(n672), .A2(n362), .ZN(n674) );
  INV_X1 U735 ( .A(n675), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n679) );
  NOR2_X1 U737 ( .A1(n675), .A2(n362), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n680), .B(KEYINPUT118), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U743 ( .A(n685), .B(KEYINPUT52), .ZN(n686) );
  NOR2_X1 U744 ( .A1(n687), .A2(n686), .ZN(n691) );
  OR2_X1 U745 ( .A1(n681), .A2(n688), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(KEYINPUT119), .ZN(n690) );
  OR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U749 ( .A1(n694), .A2(G953), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n695), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U751 ( .A1(n707), .A2(G469), .ZN(n701) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  XNOR2_X1 U753 ( .A(n697), .B(KEYINPUT120), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U755 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n712), .A2(n702), .ZN(G54) );
  NAND2_X1 U757 ( .A1(n707), .A2(G478), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n703), .B(KEYINPUT122), .ZN(n704) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n712), .A2(n706), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n707), .A2(G217), .ZN(n710) );
  XNOR2_X1 U762 ( .A(n708), .B(KEYINPUT123), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(G66) );
  NOR2_X1 U765 ( .A1(n612), .A2(G953), .ZN(n717) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n713) );
  XOR2_X1 U767 ( .A(KEYINPUT61), .B(n713), .Z(n714) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n727) );
  XNOR2_X1 U770 ( .A(n718), .B(KEYINPUT125), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U772 ( .A(G101), .B(n721), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n724), .B(KEYINPUT124), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT126), .B(n725), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(G69) );
  XOR2_X1 U777 ( .A(n729), .B(n728), .Z(n730) );
  XNOR2_X1 U778 ( .A(n731), .B(n730), .ZN(n735) );
  XOR2_X1 U779 ( .A(n735), .B(KEYINPUT127), .Z(n732) );
  XNOR2_X1 U780 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(G900), .A2(n733), .ZN(n734) );
  NAND2_X1 U782 ( .A1(n734), .A2(G953), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n613), .B(n735), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U786 ( .A(G134), .B(n740), .ZN(G36) );
endmodule

