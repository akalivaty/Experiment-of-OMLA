//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(G101), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .A4(new_n190), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT10), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT69), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT70), .A2(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT70), .A2(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(KEYINPUT65), .A3(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT66), .B1(new_n215), .B2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n203), .A3(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n206), .A2(new_n208), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(G128), .A3(new_n225), .A4(new_n217), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n220), .A2(KEYINPUT74), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT74), .B1(new_n220), .B2(new_n226), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n202), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n221), .A2(new_n223), .B1(new_n215), .B2(G146), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n226), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n193), .A2(new_n199), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n201), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n194), .A2(new_n197), .A3(new_n190), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n238), .A2(KEYINPUT84), .A3(KEYINPUT4), .A4(new_n199), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n230), .A2(new_n241), .B1(new_n219), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT84), .A2(KEYINPUT4), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n237), .A2(G101), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n229), .A2(new_n236), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT11), .A3(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT68), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n252), .A2(new_n249), .A3(KEYINPUT11), .A4(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G137), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n255), .A2(G137), .B1(KEYINPUT67), .B2(KEYINPUT11), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G131), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n249), .A2(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT67), .A2(KEYINPUT11), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n263), .B1(new_n249), .B2(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n264), .B2(new_n258), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n265), .A2(new_n266), .A3(new_n251), .A4(new_n253), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n248), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n261), .A2(new_n267), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n229), .A2(new_n270), .A3(new_n236), .A4(new_n247), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G110), .B(G140), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n273), .B(new_n275), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT12), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n220), .A2(new_n226), .A3(new_n200), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n224), .A2(new_n217), .ZN(new_n280));
  INV_X1    g094(.A(new_n232), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n200), .B1(new_n282), .B2(new_n226), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n278), .B(new_n268), .C1(new_n279), .C2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n268), .B1(new_n279), .B2(new_n283), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT12), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n271), .A2(new_n276), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n272), .A2(new_n277), .B1(new_n287), .B2(KEYINPUT85), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n289), .B(new_n276), .C1(new_n269), .C2(new_n271), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n187), .A2(new_n188), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n269), .A2(new_n271), .A3(new_n276), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n286), .A2(new_n284), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n276), .B1(new_n296), .B2(new_n271), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n291), .B(new_n293), .C1(new_n187), .C2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT9), .B(G234), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n301), .B2(G902), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G217), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n301), .A2(new_n304), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(G107), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT70), .B(G128), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G143), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT91), .B1(new_n231), .B2(G143), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT91), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n215), .A3(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n314), .A3(new_n255), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT13), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(KEYINPUT92), .A3(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT13), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n310), .A4(new_n322), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n308), .B(new_n316), .C1(new_n323), .C2(G134), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n307), .A2(new_n196), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT14), .A3(G122), .ZN(new_n327));
  XOR2_X1   g141(.A(G116), .B(G122), .Z(new_n328));
  OAI211_X1 g142(.A(G107), .B(new_n327), .C1(new_n328), .C2(KEYINPUT14), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n255), .B1(new_n310), .B2(new_n314), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n325), .B(new_n329), .C1(new_n316), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n306), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n308), .B1(new_n323), .B2(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n315), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n331), .A3(new_n305), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT93), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n335), .A2(KEYINPUT93), .A3(new_n331), .A4(new_n305), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n188), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n341));
  NOR2_X1   g155(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n342));
  OAI21_X1  g156(.A(G478), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n340), .B(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n303), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G125), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n346), .A2(KEYINPUT16), .A3(G140), .ZN(new_n347));
  XNOR2_X1  g161(.A(G125), .B(G140), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(KEYINPUT16), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(G146), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT89), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n274), .A3(G214), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(G143), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G131), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n266), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT17), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(KEYINPUT17), .A3(G131), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n350), .A2(new_n363), .A3(new_n351), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n353), .A2(new_n361), .A3(new_n362), .A4(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT18), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n356), .B1(new_n366), .B2(new_n266), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n348), .B(new_n203), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n367), .B(new_n368), .C1(new_n358), .C2(new_n366), .ZN(new_n369));
  XOR2_X1   g183(.A(G113), .B(G122), .Z(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT88), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(new_n189), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n365), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n358), .A2(new_n359), .ZN(new_n375));
  XOR2_X1   g189(.A(new_n348), .B(KEYINPUT19), .Z(new_n376));
  OAI21_X1  g190(.A(new_n351), .B1(new_n376), .B2(G146), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n369), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n372), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G475), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n188), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n374), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n373), .B1(new_n365), .B2(new_n369), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n188), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT90), .B(G475), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(KEYINPUT20), .A3(new_n381), .A4(new_n188), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G214), .B1(G237), .B2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n274), .A2(G952), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(G234), .B2(G237), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(KEYINPUT21), .B(G898), .Z(new_n397));
  NAND2_X1  g211(.A1(G234), .A2(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(G902), .A3(G953), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G224), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G953), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n219), .A2(new_n243), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n280), .B2(new_n240), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G125), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n220), .A2(new_n346), .A3(new_n226), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n403), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n408), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n244), .A2(new_n346), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT86), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(new_n402), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n418));
  INV_X1    g232(.A(G119), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G116), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT72), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n326), .B2(G119), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n326), .A2(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(KEYINPUT72), .A3(G116), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(G113), .B(new_n420), .C1(new_n425), .C2(new_n418), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT2), .B(G113), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n234), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n239), .A2(new_n246), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n425), .A2(KEYINPUT71), .A3(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n425), .B2(KEYINPUT71), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n437), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n436), .B(new_n429), .C1(new_n430), .C2(new_n433), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n417), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G210), .B1(G237), .B2(G902), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n436), .B(KEYINPUT8), .ZN(new_n444));
  INV_X1    g258(.A(new_n429), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n234), .B1(new_n428), .B2(new_n426), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n403), .A2(KEYINPUT7), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n412), .B2(new_n413), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n406), .A2(KEYINPUT7), .A3(new_n403), .A4(new_n408), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n447), .A2(new_n440), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(new_n188), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n442), .A2(new_n443), .A3(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n443), .B(KEYINPUT87), .Z(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n442), .B2(new_n452), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n393), .B(new_n400), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n345), .A2(new_n392), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G472), .A2(G902), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT76), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n249), .A2(G134), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n256), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n267), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n227), .B2(new_n228), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT73), .B1(new_n268), .B2(new_n244), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n465), .B(new_n433), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(G101), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n354), .A2(new_n274), .A3(G210), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n470), .B(new_n471), .Z(new_n472));
  AND2_X1   g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n465), .B(KEYINPUT30), .C1(new_n466), .C2(new_n467), .ZN(new_n474));
  INV_X1    g288(.A(new_n433), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n476));
  NAND2_X1  g290(.A1(new_n268), .A2(new_n244), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n267), .A2(new_n463), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n220), .B2(new_n226), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n475), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n461), .B1(new_n483), .B2(KEYINPUT31), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT31), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT75), .B(new_n485), .C1(new_n473), .C2(new_n482), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n475), .B1(new_n478), .B2(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n468), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n465), .A2(new_n433), .A3(new_n477), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n492), .A2(new_n489), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n473), .A2(new_n485), .A3(new_n482), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n460), .B1(new_n487), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n474), .A2(new_n475), .A3(new_n481), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n468), .A2(new_n472), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT31), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT75), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n483), .A2(new_n461), .A3(KEYINPUT31), .ZN(new_n502));
  AND4_X1   g316(.A1(new_n460), .A2(new_n496), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n459), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n459), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT76), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n487), .A2(new_n460), .A3(new_n496), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT32), .ZN(new_n512));
  OR3_X1    g326(.A1(new_n491), .A2(new_n493), .A3(new_n488), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n482), .A2(new_n468), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n488), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n475), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n468), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT28), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT78), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n524), .B2(new_n493), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n493), .A2(new_n524), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT29), .A3(new_n472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n518), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n519), .A2(new_n528), .A3(new_n188), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G472), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n506), .A2(new_n512), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n212), .A2(new_n419), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n231), .A2(G119), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT23), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n419), .B2(G128), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n536), .A2(new_n537), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n535), .B1(new_n309), .B2(G119), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n538), .B(new_n540), .C1(new_n542), .C2(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT79), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  OAI211_X1 g359(.A(new_n541), .B(new_n544), .C1(new_n542), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n348), .A2(new_n203), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n351), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n542), .A2(new_n545), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n536), .A2(new_n540), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n352), .B(new_n549), .C1(new_n550), .C2(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(KEYINPUT80), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(KEYINPUT22), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G137), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT80), .B1(new_n548), .B2(new_n551), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n552), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(new_n560), .B2(new_n555), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT82), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n304), .B1(G234), .B2(new_n188), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT81), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT25), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n561), .A2(new_n188), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n552), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n555), .B1(new_n572), .B2(new_n558), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n552), .A2(new_n556), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n188), .A3(new_n574), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n563), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n565), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n532), .A2(new_n533), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n533), .B1(new_n532), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n458), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  OAI21_X1  g397(.A(new_n188), .B1(new_n497), .B2(new_n503), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n511), .B1(new_n584), .B2(G472), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n579), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n338), .A2(new_n588), .A3(new_n339), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n333), .A2(new_n336), .A3(KEYINPUT33), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(G902), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n340), .A2(new_n591), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n391), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n443), .B1(new_n442), .B2(new_n452), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n393), .B1(new_n453), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT95), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n602), .B(new_n393), .C1(new_n453), .C2(new_n599), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n400), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n598), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n587), .A2(new_n303), .A3(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NOR3_X1   g422(.A1(new_n604), .A2(new_n391), .A3(new_n344), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n587), .A2(new_n303), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G107), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NAND2_X1  g426(.A1(new_n548), .A2(new_n551), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n556), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n564), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n577), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n458), .A2(new_n585), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT37), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n538), .ZN(G12));
  NAND2_X1  g434(.A1(new_n442), .A2(new_n452), .ZN(new_n621));
  INV_X1    g435(.A(new_n443), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n442), .A2(new_n443), .A3(new_n452), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n602), .B1(new_n625), .B2(new_n393), .ZN(new_n626));
  INV_X1    g440(.A(new_n603), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n303), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n399), .A2(G900), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n396), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n344), .A2(new_n391), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n532), .A2(new_n617), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  INV_X1    g449(.A(new_n515), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n488), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n188), .B1(new_n522), .B2(new_n472), .ZN(new_n638));
  OAI21_X1  g452(.A(G472), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n506), .A2(new_n512), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n453), .A2(new_n455), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT97), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT38), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n392), .A2(new_n344), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n640), .A2(new_n393), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n631), .B(KEYINPUT39), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n303), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT40), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n645), .A2(new_n649), .A3(new_n617), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n215), .ZN(G45));
  NAND3_X1  g465(.A1(new_n595), .A2(new_n391), .A3(new_n631), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n595), .A2(new_n391), .A3(KEYINPUT98), .A4(new_n631), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n532), .A2(new_n617), .A3(new_n629), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  OAI21_X1  g474(.A(new_n188), .B1(new_n288), .B2(new_n290), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(G469), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n302), .A3(new_n291), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT99), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n302), .A3(new_n291), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n532), .A2(new_n605), .A3(new_n579), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT41), .B(G113), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G15));
  NAND2_X1  g485(.A1(new_n509), .A2(new_n510), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT32), .B1(new_n672), .B2(new_n459), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n505), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n578), .B1(new_n675), .B2(new_n531), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n609), .A4(new_n668), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n532), .A2(new_n579), .A3(new_n609), .A4(new_n668), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT101), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NAND2_X1  g497(.A1(new_n601), .A2(new_n603), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n665), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n532), .A2(new_n344), .A3(new_n617), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n392), .A2(new_n400), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n419), .ZN(G21));
  OAI211_X1 g503(.A(new_n495), .B(new_n500), .C1(new_n527), .C2(new_n472), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n584), .A2(G472), .B1(new_n459), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n604), .B1(new_n664), .B2(new_n667), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n692), .A3(new_n579), .A4(new_n644), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  AND4_X1   g508(.A1(new_n628), .A2(new_n654), .A3(new_n656), .A4(new_n663), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n617), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n690), .A2(new_n459), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n509), .B2(new_n510), .ZN(new_n699));
  INV_X1    g513(.A(G472), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n617), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n628), .A2(new_n654), .A3(new_n663), .A4(new_n656), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT102), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  AND2_X1   g519(.A1(new_n302), .A2(new_n393), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n641), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n295), .B2(new_n297), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n294), .A2(KEYINPUT103), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(G469), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n291), .A3(new_n293), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n655), .A2(new_n714), .A3(new_n657), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n532), .A2(new_n579), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n532), .A2(new_n719), .A3(new_n715), .A4(new_n579), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n673), .B2(new_n674), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n722), .B(new_n531), .C1(KEYINPUT105), .C2(new_n673), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n579), .A4(new_n715), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT106), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  INV_X1    g541(.A(new_n714), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n676), .A2(new_n633), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n255), .ZN(G36));
  INV_X1    g544(.A(new_n595), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n391), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT43), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  INV_X1    g548(.A(new_n617), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n585), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n585), .A2(new_n735), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT108), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n733), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n711), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n298), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(G469), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT107), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n744), .A3(new_n747), .A4(G469), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n292), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n749), .A2(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n291), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n302), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(new_n646), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n741), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n641), .A2(new_n393), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n739), .B2(new_n740), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT109), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(KEYINPUT47), .B(new_n302), .C1(new_n750), .C2(new_n751), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n755), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n532), .A2(new_n655), .A3(new_n657), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n578), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  OAI21_X1  g581(.A(KEYINPUT113), .B1(new_n344), .B2(new_n391), .ZN(new_n768));
  MUX2_X1   g582(.A(KEYINPUT113), .B(new_n768), .S(new_n596), .Z(new_n769));
  NAND4_X1  g583(.A1(new_n587), .A2(new_n303), .A3(new_n457), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n582), .A2(new_n618), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n679), .B(new_n677), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n669), .B(new_n693), .C1(new_n686), .C2(new_n687), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n775), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT112), .B1(new_n777), .B2(new_n681), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n772), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n755), .A2(new_n632), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n532), .A2(new_n345), .A3(new_n392), .A4(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n691), .A2(new_n715), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n617), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n729), .B1(new_n721), .B2(new_n724), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n631), .A2(KEYINPUT114), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n631), .A2(KEYINPUT114), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n577), .A2(new_n616), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n302), .ZN(new_n789));
  INV_X1    g603(.A(new_n713), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n788), .A2(new_n789), .A3(new_n684), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n640), .A3(new_n644), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n704), .A2(new_n634), .A3(new_n659), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n784), .B(new_n785), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n779), .A2(new_n780), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n793), .B(KEYINPUT52), .ZN(new_n799));
  INV_X1    g613(.A(new_n729), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n725), .A2(new_n800), .A3(new_n784), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n777), .A2(new_n681), .A3(KEYINPUT112), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n771), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n780), .B1(new_n779), .B2(new_n797), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n771), .A2(new_n773), .A3(new_n775), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n675), .A2(new_n395), .A3(new_n639), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n662), .A2(new_n291), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n708), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n578), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n813), .A2(new_n598), .A3(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n579), .A2(new_n691), .A3(new_n395), .A4(new_n733), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n394), .B(new_n818), .C1(new_n685), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n733), .A2(new_n395), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n816), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n723), .A2(new_n579), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT48), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n643), .A2(new_n393), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n819), .A2(new_n663), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n819), .A2(KEYINPUT50), .A3(new_n663), .A4(new_n826), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n813), .A2(new_n817), .A3(new_n391), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n731), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n814), .A2(new_n302), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n764), .B(new_n819), .C1(new_n763), .C2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n821), .A2(new_n701), .A3(new_n816), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT115), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n832), .A2(new_n834), .A3(new_n839), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n825), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n807), .A2(new_n812), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  OR2_X1    g661(.A1(G952), .A2(G953), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n807), .A2(new_n845), .A3(new_n849), .A4(new_n812), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n579), .A2(new_n706), .A3(new_n732), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT110), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT49), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n815), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT111), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n640), .B(new_n643), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  OAI221_X1 g671(.A(new_n857), .B1(new_n856), .B2(new_n855), .C1(KEYINPUT49), .C2(new_n814), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n851), .A2(KEYINPUT118), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(G75));
  AND2_X1   g677(.A1(new_n808), .A2(new_n811), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n188), .ZN(new_n865));
  INV_X1    g679(.A(new_n454), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n441), .A2(new_n438), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n417), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT55), .Z(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n865), .A2(KEYINPUT119), .A3(new_n866), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n869), .A2(new_n870), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n865), .A2(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n873), .B1(new_n877), .B2(KEYINPUT56), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n274), .A2(G952), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(G51));
  XNOR2_X1  g695(.A(new_n864), .B(new_n809), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n292), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n883), .A2(new_n292), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n288), .A2(new_n290), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n865), .A2(new_n746), .A3(new_n748), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n879), .B1(new_n888), .B2(new_n889), .ZN(G54));
  NAND3_X1  g704(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(new_n380), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n880), .ZN(G60));
  XNOR2_X1  g707(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n591), .A2(new_n188), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n894), .B(new_n895), .Z(new_n896));
  AND4_X1   g710(.A1(new_n589), .A2(new_n882), .A3(new_n590), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n807), .A2(new_n812), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n898), .A2(new_n896), .B1(new_n589), .B2(new_n590), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n897), .A2(new_n879), .A3(new_n899), .ZN(G63));
  XNOR2_X1  g714(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n901));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n864), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n615), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n880), .C1(new_n562), .C2(new_n904), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(G66));
  INV_X1    g722(.A(new_n397), .ZN(new_n909));
  OAI21_X1  g723(.A(G953), .B1(new_n909), .B2(new_n401), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n805), .B2(G953), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n871), .B1(G898), .B2(new_n274), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT123), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT124), .Z(G69));
  NAND2_X1  g729(.A1(new_n474), .A2(new_n481), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n376), .ZN(new_n917));
  NAND2_X1  g731(.A1(G900), .A2(G953), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n723), .A2(new_n579), .A3(new_n628), .A4(new_n644), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n753), .A2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n920), .A2(new_n785), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT126), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n704), .A2(new_n634), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n659), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n757), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g740(.A(KEYINPUT126), .B(new_n924), .C1(new_n754), .C2(new_n756), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n766), .B(new_n921), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n917), .B(new_n918), .C1(new_n928), .C2(G953), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT127), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n924), .A2(new_n650), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  INV_X1    g747(.A(new_n648), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n769), .A2(new_n764), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n934), .B(new_n935), .C1(new_n580), .C2(new_n581), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n933), .A2(new_n757), .A3(new_n766), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n274), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n917), .B(KEYINPUT125), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n929), .B(new_n931), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n930), .A2(KEYINPUT127), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n940), .B(new_n941), .Z(G72));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n928), .B2(new_n779), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n488), .A3(new_n636), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n937), .B2(new_n779), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n879), .B1(new_n947), .B2(new_n637), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n516), .A2(new_n483), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n944), .B(new_n949), .C1(new_n798), .C2(new_n806), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n946), .A2(new_n948), .A3(new_n950), .ZN(G57));
endmodule


