//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338, new_n1339, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1348, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1409, new_n1410, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT65), .B(G238), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n205), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n208), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G274), .ZN(new_n244));
  AND2_X1   g0044(.A1(G1), .A2(G13), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n248), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n258));
  MUX2_X1   g0058(.A(G222), .B(G223), .S(G1698), .Z(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n258), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G77), .ZN(new_n267));
  OAI221_X1 g0067(.A(new_n251), .B1(new_n256), .B2(new_n257), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G200), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n214), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n277), .B1(new_n248), .B2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n279), .B2(new_n274), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n202), .A2(G20), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n215), .A2(new_n260), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n260), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT68), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(new_n209), .A3(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n281), .B1(new_n282), .B2(new_n283), .C1(new_n285), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n280), .B1(new_n291), .B2(new_n277), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI211_X1 g0094(.A(KEYINPUT9), .B(new_n280), .C1(new_n291), .C2(new_n277), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n271), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT10), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n268), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G179), .B2(new_n268), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n292), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G244), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n251), .B1(new_n256), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n266), .A2(G232), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G107), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(G1698), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n306), .B1(new_n307), .B2(new_n266), .C1(new_n308), .C2(new_n218), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n304), .B1(new_n309), .B2(new_n258), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G20), .A2(G77), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n313), .B1(new_n286), .B2(new_n283), .C1(new_n285), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n277), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n273), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n278), .A2(G77), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n312), .B(new_n320), .C1(G169), .C2(new_n310), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n310), .A2(G190), .ZN(new_n322));
  INV_X1    g0122(.A(new_n320), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n310), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n297), .A2(new_n302), .A3(new_n327), .ZN(new_n328));
  AOI211_X1 g0128(.A(G68), .B(new_n272), .C1(KEYINPUT72), .C2(KEYINPUT12), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n210), .B2(new_n279), .ZN(new_n332));
  INV_X1    g0132(.A(new_n277), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n284), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n334));
  INV_X1    g0134(.A(new_n283), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G50), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT11), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  INV_X1    g0141(.A(G238), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n251), .B1(new_n256), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n257), .A2(G1698), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(new_n261), .A3(new_n263), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT69), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT69), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n266), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n261), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT70), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n254), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n349), .A2(KEYINPUT70), .A3(new_n352), .ZN(new_n356));
  AOI211_X1 g0156(.A(KEYINPUT13), .B(new_n343), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n353), .A2(new_n354), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n356), .A3(new_n258), .ZN(new_n360));
  INV_X1    g0160(.A(new_n343), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n341), .B(G169), .C1(new_n357), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n350), .A2(new_n351), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n348), .B2(new_n346), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n258), .B1(new_n365), .B2(KEYINPUT70), .ZN(new_n366));
  INV_X1    g0166(.A(new_n356), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n360), .A2(new_n358), .A3(new_n361), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(G179), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n341), .B1(new_n373), .B2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n340), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(G190), .A3(new_n370), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n376), .A2(new_n339), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n373), .B2(G200), .ZN(new_n379));
  AOI211_X1 g0179(.A(KEYINPUT71), .B(new_n324), .C1(new_n369), .C2(new_n370), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n215), .A2(KEYINPUT7), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n262), .A2(G33), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT74), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n261), .A2(new_n263), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n266), .B2(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n210), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n211), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G20), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n335), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n383), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n395), .A2(KEYINPUT73), .A3(new_n396), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n215), .B1(new_n211), .B2(new_n393), .ZN(new_n401));
  INV_X1    g0201(.A(G159), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n283), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n264), .B2(new_n215), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n266), .A2(new_n384), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n398), .A2(new_n409), .A3(new_n277), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n290), .A2(new_n278), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n272), .B2(new_n290), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n253), .A2(G232), .A3(new_n254), .A4(new_n255), .ZN(new_n415));
  NOR2_X1   g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n257), .B2(G1698), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n266), .B1(G33), .B2(G87), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n251), .B(new_n415), .C1(new_n418), .C2(new_n254), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(new_n311), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(G169), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n414), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n414), .B2(new_n422), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT75), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n414), .A2(new_n422), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT18), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT75), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n414), .A2(new_n422), .A3(new_n423), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n419), .A2(G200), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n257), .A2(G1698), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G223), .B2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G87), .ZN(new_n435));
  OAI22_X1  g0235(.A1(new_n434), .A2(new_n264), .B1(new_n260), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n258), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n437), .A2(G190), .A3(new_n251), .A4(new_n415), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n439), .A2(new_n410), .A3(new_n413), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT17), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n426), .A2(new_n431), .A3(new_n441), .ZN(new_n442));
  OR3_X1    g0242(.A1(new_n328), .A2(new_n382), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n254), .A2(G274), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n248), .A2(G45), .ZN(new_n452));
  INV_X1    g0252(.A(new_n449), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n258), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n451), .B1(G270), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n261), .A2(new_n263), .A3(G257), .A4(new_n305), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n261), .A2(new_n263), .A3(G264), .A4(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(G303), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n457), .B(new_n458), .C1(new_n459), .C2(new_n266), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n258), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n298), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n276), .A2(new_n214), .B1(G20), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n215), .C1(G33), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n272), .A2(G116), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n248), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n272), .A2(new_n475), .A3(new_n214), .A4(new_n276), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n474), .B1(new_n477), .B2(G116), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n472), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n473), .B1(new_n472), .B2(new_n478), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n462), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n454), .A2(new_n247), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n450), .A2(new_n254), .ZN(new_n485));
  INV_X1    g0285(.A(G270), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(new_n258), .B2(new_n460), .ZN(new_n488));
  OAI211_X1 g0288(.A(G179), .B(new_n488), .C1(new_n479), .C2(new_n480), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n462), .B(KEYINPUT21), .C1(new_n479), .C2(new_n480), .ZN(new_n490));
  AND3_X1   g0290(.A1(new_n483), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n215), .B1(new_n351), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(KEYINPUT83), .B(new_n215), .C1(new_n351), .C2(new_n492), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n435), .A2(new_n466), .A3(new_n307), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n210), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n266), .A2(new_n499), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n333), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n476), .A2(new_n435), .ZN(new_n503));
  INV_X1    g0303(.A(new_n314), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n272), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n303), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(G238), .B2(G1698), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n264), .B1(new_n260), .B2(new_n463), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n452), .B(KEYINPUT81), .ZN(new_n510));
  INV_X1    g0310(.A(G250), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n258), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n509), .A2(new_n258), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT80), .B1(new_n444), .B2(new_n452), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n247), .A2(new_n515), .A3(new_n446), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(G190), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT81), .B1(new_n248), .B2(G45), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n446), .A2(KEYINPUT81), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(G250), .A4(new_n254), .ZN(new_n522));
  AND2_X1   g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G238), .A2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n303), .B2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n523), .B1(new_n525), .B2(new_n266), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n522), .B1(new_n526), .B2(new_n254), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n515), .B1(new_n247), .B2(new_n446), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n515), .A2(new_n254), .A3(G274), .A4(new_n446), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G200), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n506), .A2(new_n518), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n476), .A2(new_n314), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n502), .A2(new_n505), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G169), .B1(new_n527), .B2(new_n530), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n513), .A2(G179), .A3(new_n517), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n534), .B1(new_n537), .B2(KEYINPUT82), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT82), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n532), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n488), .A2(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n456), .A2(new_n461), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G200), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n472), .A2(new_n478), .A3(new_n473), .ZN(new_n545));
  INV_X1    g0345(.A(new_n480), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n491), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n215), .A2(KEYINPUT85), .A3(G87), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n264), .B2(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n215), .A2(KEYINPUT85), .A3(G87), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n266), .A2(KEYINPUT22), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n215), .B2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n307), .A2(KEYINPUT23), .A3(G20), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n555), .A2(new_n556), .B1(new_n215), .B2(new_n523), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n551), .A2(KEYINPUT24), .A3(new_n553), .A4(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n277), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n273), .A2(new_n563), .A3(new_n307), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT25), .B1(new_n272), .B2(G107), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n307), .C2(new_n476), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n333), .A2(G107), .A3(new_n272), .A4(new_n475), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(KEYINPUT86), .A3(new_n564), .A4(new_n565), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n450), .A2(G264), .A3(new_n254), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n260), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G250), .A2(G1698), .ZN(new_n576));
  INV_X1    g0376(.A(G257), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1698), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n578), .B2(new_n266), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n484), .B(new_n573), .C1(new_n579), .C2(new_n254), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT87), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n581), .A3(G169), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n511), .A2(new_n305), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(G1698), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n264), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n258), .B1(new_n586), .B2(new_n575), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n587), .A2(G179), .A3(new_n484), .A4(new_n573), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n581), .B1(new_n580), .B2(G169), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n572), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT88), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n580), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G190), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n580), .A2(G200), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n562), .A3(new_n571), .A4(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n572), .B(KEYINPUT88), .C1(new_n589), .C2(new_n590), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n484), .B1(new_n485), .B2(new_n577), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(new_n305), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(KEYINPUT77), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n465), .B(new_n606), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT77), .B1(new_n602), .B2(new_n603), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n601), .B1(new_n609), .B2(new_n254), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n298), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT76), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n261), .A2(new_n263), .A3(new_n387), .ZN(new_n613));
  OAI211_X1 g0413(.A(KEYINPUT7), .B(new_n215), .C1(new_n261), .C2(new_n387), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(G107), .C1(new_n615), .C2(new_n406), .ZN(new_n616));
  XNOR2_X1  g0416(.A(G97), .B(G107), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT6), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n466), .A3(G107), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n622), .A2(G20), .B1(G77), .B2(new_n335), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n307), .B1(new_n389), .B2(new_n391), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n612), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n277), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n273), .A2(new_n466), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n476), .B2(new_n466), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n607), .A2(new_n608), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n254), .B1(new_n632), .B2(new_n604), .ZN(new_n633));
  NOR4_X1   g0433(.A1(new_n633), .A2(KEYINPUT79), .A3(G179), .A4(new_n600), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT79), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n602), .A2(new_n603), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT77), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n305), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n606), .A2(new_n465), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n638), .A2(new_n604), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n600), .B1(new_n641), .B2(new_n258), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n635), .B1(new_n642), .B2(new_n311), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n611), .B(new_n631), .C1(new_n634), .C2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(G190), .B(new_n601), .C1(new_n609), .C2(new_n254), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT78), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n215), .B1(new_n385), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n390), .A2(new_n648), .B1(new_n386), .B2(new_n388), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT76), .B1(new_n649), .B2(new_n307), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n616), .A3(new_n623), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n629), .B1(new_n651), .B2(new_n277), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT78), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n642), .A2(new_n653), .A3(G190), .ZN(new_n654));
  OAI21_X1  g0454(.A(G200), .B1(new_n633), .B2(new_n600), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n646), .A2(new_n652), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n443), .A2(new_n548), .A3(new_n599), .A4(new_n657), .ZN(G372));
  NOR2_X1   g0458(.A1(new_n424), .A2(new_n425), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n376), .A2(new_n339), .ZN(new_n661));
  OAI21_X1  g0461(.A(G200), .B1(new_n357), .B2(new_n362), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT71), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n373), .A2(new_n378), .A3(G200), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n375), .B1(new_n665), .B2(new_n321), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n660), .B1(new_n666), .B2(new_n441), .ZN(new_n667));
  INV_X1    g0467(.A(new_n297), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n302), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n534), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n537), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n634), .A2(new_n643), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n620), .B1(new_n617), .B2(new_n618), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n674), .A2(new_n215), .B1(new_n317), .B2(new_n283), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n625), .B2(new_n612), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n333), .B1(new_n676), .B2(new_n650), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n611), .B1(new_n677), .B2(new_n629), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n656), .B(new_n597), .C1(new_n673), .C2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n483), .A2(new_n591), .A3(new_n489), .A4(new_n490), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  INV_X1    g0481(.A(new_n503), .ZN(new_n682));
  INV_X1    g0482(.A(new_n505), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n498), .A2(new_n501), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n333), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n324), .B1(new_n513), .B2(new_n517), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n506), .A2(KEYINPUT89), .A3(new_n531), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n518), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n672), .B1(new_n679), .B2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n311), .B(new_n601), .C1(new_n609), .C2(new_n254), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT79), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n642), .A2(new_n635), .A3(new_n311), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n627), .A2(new_n630), .B1(new_n610), .B2(new_n298), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n541), .A2(KEYINPUT26), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT26), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n689), .A2(new_n695), .A3(new_n696), .A4(new_n672), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n697), .A2(KEYINPUT90), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT90), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT26), .A4(new_n541), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n691), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n670), .B1(new_n443), .B2(new_n704), .ZN(G369));
  NAND3_X1  g0505(.A1(new_n248), .A2(new_n215), .A3(G13), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(KEYINPUT27), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G213), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G343), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n591), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n599), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n572), .A2(new_n711), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(KEYINPUT91), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT91), .B1(new_n714), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n546), .A2(new_n545), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n711), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n491), .A2(new_n547), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n483), .A2(new_n489), .A3(new_n490), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n720), .A3(new_n711), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n591), .A2(new_n711), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n714), .A2(new_n715), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n491), .A2(new_n711), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n716), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n206), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n497), .A2(G116), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n212), .B2(new_n738), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT28), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n593), .A2(new_n598), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n491), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n644), .A2(new_n597), .A3(new_n656), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n689), .A2(new_n672), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n527), .A2(new_n530), .A3(new_n311), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n298), .B1(new_n513), .B2(new_n517), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT82), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n540), .A3(new_n671), .ZN(new_n752));
  INV_X1    g0552(.A(new_n532), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n695), .A2(new_n752), .A3(new_n696), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(KEYINPUT26), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n672), .B(KEYINPUT93), .Z(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n699), .A2(KEYINPUT26), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n748), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n712), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .ZN(new_n761));
  INV_X1    g0561(.A(new_n657), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n483), .A2(new_n547), .A3(new_n489), .A4(new_n490), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(new_n753), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n762), .A2(new_n765), .A3(new_n714), .A4(new_n712), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n527), .A2(new_n530), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n573), .B1(new_n579), .B2(new_n254), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n488), .A2(new_n768), .A3(G179), .A4(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n767), .B1(new_n771), .B2(new_n610), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n543), .A2(new_n311), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n513), .A2(new_n517), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n769), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n773), .A2(new_n775), .A3(KEYINPUT30), .A4(new_n642), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n543), .A2(new_n774), .A3(new_n311), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n610), .A2(KEYINPUT92), .A3(new_n580), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT92), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(new_n642), .B2(new_n594), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n711), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT31), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(KEYINPUT31), .B(new_n711), .C1(new_n777), .C2(new_n782), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n766), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G330), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT90), .B1(new_n754), .B2(new_n698), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n699), .A2(new_n698), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(new_n703), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n672), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n680), .A2(new_n689), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n746), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT29), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n795), .A2(new_n796), .A3(new_n712), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n761), .A2(new_n788), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n742), .B1(new_n799), .B2(G1), .ZN(G364));
  AND2_X1   g0600(.A1(new_n215), .A2(G13), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n248), .B1(new_n801), .B2(G45), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n737), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n727), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G330), .B2(new_n725), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n245), .B1(new_n215), .B2(G169), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT95), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n215), .A2(G179), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(new_n269), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n307), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G190), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G159), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n813), .B1(new_n817), .B2(KEYINPUT32), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n269), .A2(G179), .A3(G200), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n215), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G97), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n215), .A2(new_n311), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G200), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n269), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n818), .B(new_n822), .C1(new_n274), .C2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n811), .A2(G190), .A3(G200), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G87), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n824), .A2(G190), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n817), .B2(KEYINPUT32), .C1(new_n832), .C2(new_n210), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n823), .A2(new_n814), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n823), .A2(G190), .A3(new_n324), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n266), .B1(new_n834), .B2(new_n317), .C1(new_n209), .C2(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n827), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G322), .B1(new_n816), .B2(G329), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n839), .B(new_n264), .C1(new_n840), .C2(new_n834), .ZN(new_n841));
  INV_X1    g0641(.A(G317), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(KEYINPUT33), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n842), .A2(KEYINPUT33), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n831), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n825), .A2(G326), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(new_n459), .C2(new_n828), .ZN(new_n847));
  INV_X1    g0647(.A(G283), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n820), .A2(new_n574), .B1(new_n812), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n841), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n810), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n736), .A2(new_n264), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G355), .B1(new_n463), .B2(new_n736), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n266), .B(new_n736), .C1(new_n213), .C2(new_n445), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT94), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n445), .B2(new_n242), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n854), .A2(KEYINPUT94), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(G13), .A2(G33), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(G20), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n810), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n851), .A2(new_n864), .A3(new_n804), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT97), .Z(new_n866));
  INV_X1    g0666(.A(new_n861), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n725), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n806), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G396));
  INV_X1    g0670(.A(new_n804), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n320), .A2(new_n711), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n321), .A2(new_n325), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT98), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n321), .A2(new_n325), .A3(KEYINPUT98), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n321), .A2(new_n712), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n795), .B2(new_n712), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT99), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n712), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n795), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT99), .B1(new_n704), .B2(new_n882), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n788), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n871), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n877), .A2(new_n878), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n859), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n808), .A2(new_n860), .A3(new_n809), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n804), .B1(new_n893), .B2(G77), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n848), .A2(new_n832), .B1(new_n826), .B2(new_n459), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(G107), .B2(new_n829), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n834), .A2(new_n463), .B1(new_n815), .B2(new_n840), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n266), .B(new_n897), .C1(G294), .C2(new_n838), .ZN(new_n898));
  INV_X1    g0698(.A(new_n812), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G87), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n896), .A2(new_n822), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n834), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n838), .A2(G143), .B1(new_n902), .B2(G159), .ZN(new_n903));
  INV_X1    g0703(.A(G137), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n903), .B1(new_n832), .B2(new_n282), .C1(new_n904), .C2(new_n826), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT34), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n899), .A2(G68), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n264), .B1(new_n816), .B2(G132), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n821), .A2(G58), .B1(new_n829), .B2(G50), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n905), .A2(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n894), .B1(new_n913), .B2(new_n810), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n889), .A2(new_n890), .B1(new_n892), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(G384));
  NOR3_X1   g0716(.A1(new_n328), .A2(new_n382), .A3(new_n442), .ZN(new_n917));
  INV_X1    g0717(.A(new_n797), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n796), .B1(new_n759), .B2(new_n712), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n670), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT102), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n321), .A2(new_n711), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n881), .B1(new_n795), .B2(new_n883), .ZN(new_n925));
  AOI211_X1 g0725(.A(KEYINPUT99), .B(new_n882), .C1(new_n791), .C2(new_n794), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n391), .B1(new_n266), .B2(new_n384), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n928), .A2(G68), .B1(new_n399), .B2(new_n404), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT16), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n333), .B1(new_n929), .B2(KEYINPUT16), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n412), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n932), .A2(new_n709), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n442), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n440), .B1(new_n932), .B2(new_n709), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n420), .A2(new_n421), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT37), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n427), .A2(KEYINPUT100), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n412), .B1(new_n931), .B2(new_n398), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT37), .B1(new_n940), .B2(new_n439), .ZN(new_n941));
  INV_X1    g0741(.A(new_n709), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n414), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT100), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n414), .A2(new_n422), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n939), .A2(new_n941), .A3(new_n943), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n934), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n934), .A2(KEYINPUT38), .A3(new_n947), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(G169), .B1(new_n357), .B2(new_n362), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT14), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n371), .A3(new_n363), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n340), .B(new_n711), .C1(new_n665), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n340), .A2(new_n711), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n375), .A2(new_n381), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n927), .A2(new_n951), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n660), .A2(new_n709), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n949), .A2(KEYINPUT39), .A3(new_n950), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n427), .A2(KEYINPUT101), .A3(new_n440), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n943), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT101), .B1(new_n427), .B2(new_n440), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT37), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n946), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n943), .B1(new_n441), .B2(new_n659), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT38), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT38), .ZN(new_n971));
  AOI221_X4 g0771(.A(new_n971), .B1(new_n938), .B2(new_n946), .C1(new_n442), .C2(new_n933), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n962), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n954), .A2(new_n340), .A3(new_n712), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n961), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n959), .A2(new_n960), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n922), .B(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(KEYINPUT40), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n785), .A2(new_n786), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n891), .B1(new_n980), .B2(new_n766), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n981), .B(new_n958), .C1(new_n972), .C2(new_n948), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n375), .A2(new_n381), .A3(new_n956), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n956), .B1(new_n375), .B2(new_n381), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n787), .A2(new_n879), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n427), .A2(new_n440), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT101), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(new_n943), .A3(new_n963), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n941), .A2(new_n943), .ZN(new_n992));
  AND2_X1   g0792(.A1(new_n939), .A2(new_n945), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n991), .A2(KEYINPUT37), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n971), .B1(new_n994), .B2(new_n968), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n979), .B1(new_n995), .B2(new_n950), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n979), .A2(new_n982), .B1(new_n987), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n917), .A2(new_n787), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  INV_X1    g0800(.A(G330), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n978), .A2(new_n1002), .B1(new_n248), .B2(new_n801), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n978), .B2(new_n1002), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n622), .A2(KEYINPUT35), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n622), .A2(KEYINPUT35), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1005), .A2(G116), .A3(new_n216), .A4(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT36), .Z(new_n1008));
  NAND3_X1  g0808(.A1(new_n213), .A2(G77), .A3(new_n393), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n274), .A2(G68), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n248), .B(G13), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1004), .A2(new_n1008), .A3(new_n1011), .ZN(G367));
  OAI21_X1  g0812(.A(new_n762), .B1(new_n652), .B2(new_n712), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n701), .A2(new_n711), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n728), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n747), .B1(new_n506), .B2(new_n712), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n792), .A2(new_n685), .A3(new_n711), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT43), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n734), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n1015), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT103), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1026), .B2(new_n1015), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1013), .A2(new_n744), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n711), .B1(new_n1031), .B2(new_n644), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1022), .B(new_n1025), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1024), .A3(new_n1023), .A4(new_n1033), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1018), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1025), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1022), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1040), .A2(new_n1017), .A3(new_n1035), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n728), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1015), .B1(new_n734), .B2(new_n729), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT44), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n734), .A2(new_n729), .A3(new_n1015), .ZN(new_n1047));
  XOR2_X1   g0847(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1047), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1043), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n733), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n713), .B(new_n1052), .C1(new_n717), .C2(new_n718), .ZN(new_n1053));
  AND3_X1   g0853(.A1(new_n1053), .A2(new_n726), .A3(new_n734), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n726), .B1(new_n1053), .B2(new_n734), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n798), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1044), .B(KEYINPUT44), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1047), .B(new_n1048), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1058), .A2(new_n1059), .A3(new_n728), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1051), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n799), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n737), .B(KEYINPUT41), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n803), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1021), .A2(new_n867), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n736), .A2(new_n266), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n234), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n862), .B1(new_n206), .B2(new_n314), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n831), .A2(G294), .B1(new_n899), .B2(G97), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n840), .B2(new_n826), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n821), .A2(G107), .B1(new_n902), .B2(G283), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(KEYINPUT105), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT106), .B(G317), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n264), .B1(new_n815), .B2(new_n1073), .C1(new_n835), .C2(new_n459), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n829), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT46), .B1(new_n829), .B2(G116), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1072), .B(new_n1077), .C1(KEYINPUT105), .C2(new_n1071), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n834), .A2(new_n274), .B1(new_n815), .B2(new_n904), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G150), .B2(new_n838), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G143), .A2(new_n825), .B1(new_n831), .B2(G159), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n821), .A2(G68), .B1(new_n829), .B2(G58), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n899), .A2(G77), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n266), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT107), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1078), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT47), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n810), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n804), .B1(new_n1067), .B2(new_n1068), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT108), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1042), .A2(new_n1064), .B1(new_n1065), .B2(new_n1092), .ZN(G387));
  OAI22_X1  g0893(.A1(new_n834), .A2(new_n210), .B1(new_n815), .B2(new_n282), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n264), .B(new_n1094), .C1(G50), .C2(new_n838), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n821), .A2(new_n504), .B1(new_n899), .B2(G97), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n825), .A2(G159), .B1(new_n829), .B2(G77), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n290), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n831), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1073), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n838), .A2(new_n1101), .B1(new_n902), .B2(G303), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT109), .B(G322), .Z(new_n1103));
  OAI221_X1 g0903(.A(new_n1102), .B1(new_n832), .B2(new_n840), .C1(new_n826), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT48), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n820), .A2(new_n848), .B1(new_n828), .B2(new_n574), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n266), .B1(new_n816), .B2(G326), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n463), .C2(new_n812), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT49), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1100), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n810), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n739), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n852), .A2(new_n1115), .B1(new_n307), .B2(new_n736), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n231), .A2(new_n445), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n286), .A2(G50), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT50), .Z(new_n1119));
  OAI211_X1 g0919(.A(new_n739), .B(new_n445), .C1(new_n210), .C2(new_n317), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1066), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1116), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n871), .B1(new_n1122), .B2(new_n863), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1114), .B(new_n1123), .C1(new_n719), .C2(new_n867), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1057), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n737), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1056), .A2(new_n798), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1124), .B1(new_n802), .B2(new_n1056), .C1(new_n1126), .C2(new_n1127), .ZN(G393));
  AND2_X1   g0928(.A1(new_n239), .A2(new_n1066), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n862), .B1(new_n466), .B2(new_n206), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n804), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n820), .A2(new_n317), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n900), .B1(new_n832), .B2(new_n274), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1132), .B(new_n1133), .C1(G68), .C2(new_n829), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n826), .A2(new_n282), .B1(new_n402), .B2(new_n835), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT51), .ZN(new_n1136));
  OR2_X1    g0936(.A1(new_n834), .A2(new_n286), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n264), .B1(new_n816), .B2(G143), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n821), .A2(G116), .B1(new_n902), .B2(G294), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n459), .B2(new_n832), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT110), .Z(new_n1142));
  OAI22_X1  g0942(.A1(new_n826), .A2(new_n842), .B1(new_n840), .B2(new_n835), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT52), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n829), .A2(G283), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n264), .B1(new_n1103), .B2(new_n815), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(new_n813), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1139), .B1(new_n1142), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1131), .B1(new_n1151), .B2(new_n810), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1015), .B2(new_n867), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n1154), .B2(new_n802), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1061), .A2(new_n737), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1057), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT111), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT111), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n737), .A4(new_n1061), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1155), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G390));
  OAI21_X1  g0963(.A(new_n974), .B1(new_n970), .B2(new_n972), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n756), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n701), .A2(new_n698), .A3(new_n541), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n747), .B1(new_n743), .B2(new_n723), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1166), .C1(new_n1167), .C2(new_n679), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n758), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n883), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n924), .B1(new_n957), .B2(new_n955), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n975), .B1(new_n927), .B2(new_n958), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n961), .A2(new_n973), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1173), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n958), .A2(G330), .A3(new_n787), .A4(new_n879), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n923), .B1(new_n885), .B2(new_n884), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n974), .B1(new_n1181), .B2(new_n985), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1175), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1178), .A3(new_n1173), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT115), .B1(new_n1185), .B2(new_n802), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n828), .A2(new_n282), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT53), .ZN(new_n1188));
  INV_X1    g0988(.A(G132), .ZN(new_n1189));
  INV_X1    g0989(.A(G125), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n835), .A2(new_n1189), .B1(new_n815), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n266), .B1(new_n834), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n825), .A2(G128), .B1(new_n899), .B2(G50), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G159), .A2(new_n821), .B1(new_n831), .B2(G137), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1188), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT116), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1132), .B1(G283), .B2(new_n825), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n307), .B2(new_n832), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n835), .A2(new_n463), .B1(new_n815), .B2(new_n574), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n266), .B(new_n1202), .C1(G97), .C2(new_n902), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n830), .A3(new_n908), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1199), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n810), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n804), .C1(new_n1098), .C2(new_n893), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1175), .B2(new_n859), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT117), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT115), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1180), .A2(new_n1211), .A3(new_n1184), .A4(new_n803), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1186), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT114), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n443), .B1(new_n761), .B2(new_n797), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n443), .A2(new_n788), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1215), .A2(new_n669), .A3(new_n1216), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n548), .A2(new_n657), .A3(new_n599), .A4(new_n711), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n785), .A2(new_n786), .ZN(new_n1219));
  OAI211_X1 g1019(.A(G330), .B(new_n879), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n985), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1178), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT112), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n927), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n923), .B1(new_n759), .B2(new_n883), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1178), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1223), .B1(new_n1222), .B2(new_n927), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1217), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT113), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1221), .A2(new_n1178), .A3(new_n1225), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n885), .A2(new_n884), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1233), .A2(new_n924), .B1(new_n1221), .B2(new_n1178), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1223), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1221), .A2(new_n1178), .ZN(new_n1236));
  OAI21_X1  g1036(.A(KEYINPUT112), .B1(new_n1236), .B2(new_n1181), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(KEYINPUT113), .A3(new_n1217), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1185), .A2(new_n1231), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n887), .A2(new_n917), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n920), .A2(new_n670), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n737), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1214), .B1(new_n1240), .B2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1185), .A2(new_n1231), .A3(new_n1239), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1247), .A2(KEYINPUT114), .A3(new_n737), .A4(new_n1244), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1213), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(G378));
  NAND2_X1  g1050(.A1(new_n982), .A2(new_n979), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n987), .A2(new_n996), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(G330), .ZN(new_n1253));
  OR3_X1    g1053(.A1(new_n292), .A2(KEYINPUT55), .A3(new_n709), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT55), .B1(new_n292), .B2(new_n709), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n297), .B2(new_n302), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1259));
  NAND3_X1  g1059(.A1(new_n297), .A2(new_n1256), .A3(new_n302), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1259), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1260), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n1257), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1253), .A2(new_n1261), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1261), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n997), .A2(G330), .A3(new_n1266), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n976), .A2(new_n960), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1265), .A2(new_n1267), .A3(new_n1268), .A4(new_n959), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1266), .B1(new_n997), .B2(G330), .ZN(new_n1270));
  AND4_X1   g1070(.A1(G330), .A2(new_n1251), .A3(new_n1252), .A4(new_n1266), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n977), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n803), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n804), .B1(new_n893), .B2(G50), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n266), .A2(G41), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n829), .B2(G77), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT118), .Z(new_n1278));
  AOI22_X1  g1078(.A1(new_n838), .A2(G107), .B1(new_n816), .B2(G283), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n314), .B2(new_n834), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n821), .A2(G68), .B1(new_n899), .B2(G58), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1281), .B1(new_n466), .B2(new_n832), .C1(new_n463), .C2(new_n826), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1278), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT58), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1276), .B(new_n274), .C1(G33), .C2(G41), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n1190), .A2(new_n826), .B1(new_n832), .B2(new_n1189), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n838), .A2(G128), .B1(new_n902), .B2(G137), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n828), .B2(new_n1192), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1287), .B(new_n1289), .C1(G150), .C2(new_n821), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(KEYINPUT59), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(KEYINPUT59), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n899), .A2(G159), .ZN(new_n1294));
  AOI211_X1 g1094(.A(G33), .B(G41), .C1(new_n816), .C2(G124), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  OAI221_X1 g1096(.A(new_n1286), .B1(KEYINPUT58), .B2(new_n1283), .C1(new_n1292), .C2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1275), .B1(new_n1297), .B2(new_n810), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1266), .B2(new_n860), .ZN(new_n1299));
  XOR2_X1   g1099(.A(new_n1299), .B(KEYINPUT120), .Z(new_n1300));
  AND2_X1   g1100(.A1(new_n1274), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1178), .B1(new_n1183), .B2(new_n1173), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1179), .B(new_n1172), .C1(new_n1182), .C2(new_n1175), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1242), .B1(new_n1304), .B2(new_n1238), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1270), .A2(new_n1271), .A3(new_n977), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1265), .A2(new_n1267), .B1(new_n1268), .B2(new_n959), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT57), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n737), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1244), .A2(new_n1217), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT57), .B1(new_n1310), .B2(new_n1273), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1301), .B1(new_n1309), .B2(new_n1311), .ZN(G375));
  NAND4_X1  g1112(.A1(new_n1237), .A2(new_n1242), .A3(new_n1226), .A4(new_n1224), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT121), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1235), .A2(KEYINPUT121), .A3(new_n1242), .A4(new_n1237), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1318), .A2(new_n1063), .A3(new_n1231), .A4(new_n1239), .ZN(new_n1319));
  XOR2_X1   g1119(.A(new_n1319), .B(KEYINPUT122), .Z(new_n1320));
  NAND2_X1  g1120(.A1(new_n1238), .A2(new_n803), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n804), .B1(new_n893), .B2(G68), .ZN(new_n1322));
  OAI22_X1  g1122(.A1(new_n463), .A2(new_n832), .B1(new_n826), .B2(new_n574), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(G97), .B2(new_n829), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n821), .A2(new_n504), .ZN(new_n1325));
  OAI22_X1  g1125(.A1(new_n835), .A2(new_n848), .B1(new_n834), .B2(new_n307), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n266), .B(new_n1326), .C1(G303), .C2(new_n816), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1324), .A2(new_n1084), .A3(new_n1325), .A4(new_n1327), .ZN(new_n1328));
  AOI22_X1  g1128(.A1(new_n829), .A2(G159), .B1(new_n816), .B2(G128), .ZN(new_n1329));
  XOR2_X1   g1129(.A(new_n1329), .B(KEYINPUT123), .Z(new_n1330));
  OAI22_X1  g1130(.A1(new_n1189), .A2(new_n826), .B1(new_n832), .B2(new_n1192), .ZN(new_n1331));
  OAI221_X1 g1131(.A(new_n266), .B1(new_n834), .B2(new_n282), .C1(new_n904), .C2(new_n835), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n820), .A2(new_n274), .B1(new_n812), .B2(new_n209), .ZN(new_n1333));
  OR3_X1    g1133(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1328), .B1(new_n1330), .B2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1322), .B1(new_n1335), .B2(new_n810), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n958), .B2(new_n860), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1321), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1320), .A2(new_n1339), .ZN(G381));
  INV_X1    g1140(.A(G375), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1186), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1247), .A2(new_n737), .A3(new_n1244), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  OR2_X1    g1144(.A1(G393), .A2(G396), .ZN(new_n1345));
  NOR4_X1   g1145(.A1(G390), .A2(G387), .A3(G384), .A4(new_n1345), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1344), .A2(new_n1339), .A3(new_n1320), .A4(new_n1346), .ZN(G407));
  NAND2_X1  g1147(.A1(new_n1344), .A2(new_n710), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(G407), .A2(G213), .A3(new_n1348), .ZN(G409));
  OR2_X1    g1149(.A1(G387), .A2(new_n1162), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G387), .A2(new_n1162), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(KEYINPUT126), .B1(G387), .B2(new_n1162), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(G393), .B(new_n869), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT61), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1350), .A2(new_n1353), .A3(new_n1351), .A4(new_n1354), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1356), .A2(new_n1357), .A3(new_n1358), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1310), .A2(new_n1063), .A3(new_n1273), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1274), .A2(new_n1299), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1342), .B(new_n1343), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1362), .B1(new_n1249), .B2(G375), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n1364));
  INV_X1    g1164(.A(new_n1364), .ZN(new_n1365));
  OAI211_X1 g1165(.A(new_n1315), .B(new_n1316), .C1(new_n1243), .C2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT125), .ZN(new_n1367));
  NOR3_X1   g1167(.A1(new_n1227), .A2(new_n1217), .A3(new_n1228), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n738), .B1(new_n1368), .B2(KEYINPUT60), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1366), .A2(new_n1367), .A3(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(new_n1367), .B1(new_n1366), .B2(new_n1369), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1339), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1373), .A2(new_n915), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1365), .B1(new_n1238), .B2(new_n1217), .ZN(new_n1375));
  OAI21_X1  g1175(.A(new_n1369), .B1(new_n1317), .B2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1376), .A2(KEYINPUT125), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1377), .A2(new_n1370), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(G384), .A3(new_n1339), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n710), .A2(G213), .ZN(new_n1380));
  NAND4_X1  g1180(.A1(new_n1363), .A2(new_n1374), .A3(new_n1379), .A4(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(new_n1381), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1359), .B1(new_n1382), .B2(KEYINPUT63), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT63), .ZN(new_n1384));
  AOI21_X1  g1184(.A(G384), .B1(new_n1378), .B2(new_n1339), .ZN(new_n1385));
  AOI211_X1 g1185(.A(new_n915), .B(new_n1338), .C1(new_n1377), .C2(new_n1370), .ZN(new_n1386));
  NOR2_X1   g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  NAND3_X1  g1187(.A1(new_n710), .A2(G213), .A3(G2897), .ZN(new_n1388));
  AOI22_X1  g1188(.A1(new_n1387), .A2(new_n1388), .B1(new_n1363), .B2(new_n1380), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1388), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1390), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1391));
  AOI21_X1  g1191(.A(new_n1384), .B1(new_n1389), .B2(new_n1391), .ZN(new_n1392));
  OAI21_X1  g1192(.A(new_n1383), .B1(new_n1392), .B2(new_n1382), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1381), .A2(KEYINPUT62), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1363), .A2(new_n1380), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1374), .A2(new_n1379), .A3(new_n1388), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1395), .A2(new_n1391), .A3(new_n1396), .ZN(new_n1397));
  INV_X1    g1197(.A(KEYINPUT62), .ZN(new_n1398));
  NAND4_X1  g1198(.A1(new_n1387), .A2(new_n1398), .A3(new_n1380), .A4(new_n1363), .ZN(new_n1399));
  NAND4_X1  g1199(.A1(new_n1394), .A2(new_n1397), .A3(new_n1357), .A4(new_n1399), .ZN(new_n1400));
  INV_X1    g1200(.A(KEYINPUT127), .ZN(new_n1401));
  INV_X1    g1201(.A(new_n1358), .ZN(new_n1402));
  AOI22_X1  g1202(.A1(new_n1350), .A2(new_n1351), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1403));
  OAI21_X1  g1203(.A(new_n1401), .B1(new_n1402), .B2(new_n1403), .ZN(new_n1404));
  NAND3_X1  g1204(.A1(new_n1356), .A2(KEYINPUT127), .A3(new_n1358), .ZN(new_n1405));
  AND2_X1   g1205(.A1(new_n1404), .A2(new_n1405), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1400), .A2(new_n1406), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1393), .A2(new_n1407), .ZN(G405));
  NAND2_X1  g1208(.A1(G378), .A2(new_n1341), .ZN(new_n1409));
  NAND3_X1  g1209(.A1(G375), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1409), .A2(new_n1410), .ZN(new_n1411));
  NAND2_X1  g1211(.A1(new_n1411), .A2(new_n1387), .ZN(new_n1412));
  OAI211_X1 g1212(.A(new_n1409), .B(new_n1410), .C1(new_n1385), .C2(new_n1386), .ZN(new_n1413));
  AND4_X1   g1213(.A1(new_n1405), .A2(new_n1404), .A3(new_n1412), .A4(new_n1413), .ZN(new_n1414));
  AOI22_X1  g1214(.A1(new_n1405), .A2(new_n1404), .B1(new_n1412), .B2(new_n1413), .ZN(new_n1415));
  NOR2_X1   g1215(.A1(new_n1414), .A2(new_n1415), .ZN(G402));
endmodule


