//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(G143), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n192), .A2(G143), .ZN(new_n197));
  OAI22_X1  g011(.A1(new_n193), .A2(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(G146), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n200), .A3(new_n191), .A4(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G107), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n203), .A2(G107), .ZN(new_n206));
  OAI21_X1  g020(.A(G101), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT79), .B(G101), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n208), .A2(new_n204), .A3(new_n209), .A4(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n207), .A3(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(KEYINPUT81), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT81), .B1(new_n214), .B2(new_n215), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G134), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G137), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n229), .B2(new_n220), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(G134), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n232), .B1(new_n221), .B2(new_n225), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n220), .B1(new_n229), .B2(new_n222), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n209), .A2(new_n212), .A3(new_n204), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G101), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(KEYINPUT0), .B2(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n199), .A2(new_n200), .B1(new_n246), .B2(KEYINPUT64), .ZN(new_n247));
  INV_X1    g061(.A(new_n244), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n245), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT10), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n241), .A2(new_n253), .B1(new_n214), .B2(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n219), .A2(new_n237), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n237), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n214), .A2(new_n215), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n216), .ZN(new_n261));
  INV_X1    g075(.A(new_n255), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n190), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n213), .A2(new_n207), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n201), .A3(new_n198), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n267), .A2(new_n214), .B1(new_n231), .B2(new_n236), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n214), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT82), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n271), .A2(new_n237), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n265), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n273), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(KEYINPUT83), .C1(new_n268), .C2(new_n269), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n261), .A2(new_n257), .A3(new_n262), .ZN(new_n278));
  INV_X1    g092(.A(new_n190), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n264), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G469), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT72), .B(G902), .Z(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n270), .A2(new_n274), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n190), .B1(new_n256), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n237), .B1(new_n219), .B2(new_n255), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n278), .A3(new_n279), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(G469), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n284), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G125), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n202), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n199), .A2(new_n200), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n246), .A2(KEYINPUT64), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n244), .A3(new_n243), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n249), .A2(new_n248), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(G125), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G224), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(G953), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n295), .B(new_n300), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G119), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT2), .B(G113), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n312), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n240), .A2(new_n315), .A3(new_n252), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n307), .A3(G116), .ZN(new_n319));
  OAI211_X1 g133(.A(G113), .B(new_n319), .C1(new_n311), .C2(new_n318), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n313), .A2(new_n320), .A3(new_n207), .A4(new_n213), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n295), .A2(new_n300), .ZN(new_n323));
  INV_X1    g137(.A(new_n302), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(KEYINPUT7), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n317), .B(new_n326), .ZN(new_n327));
  AND4_X1   g141(.A1(new_n313), .A2(new_n320), .A3(new_n207), .A4(new_n213), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n313), .A2(new_n320), .B1(new_n213), .B2(new_n207), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n322), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n306), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G210), .B1(G237), .B2(G902), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n316), .A2(new_n321), .ZN(new_n334));
  INV_X1    g148(.A(new_n317), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT6), .A3(new_n322), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n323), .B(new_n324), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n334), .A2(new_n339), .A3(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n332), .A2(new_n333), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n333), .B1(new_n332), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G214), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT9), .B(G234), .ZN(new_n348));
  OAI21_X1  g162(.A(G221), .B1(new_n348), .B2(G902), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n349), .B(KEYINPUT78), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n293), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G237), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(G214), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n195), .ZN(new_n356));
  NOR2_X1   g170(.A1(G237), .A2(G953), .ZN(new_n357));
  AOI21_X1  g171(.A(G143), .B1(new_n357), .B2(G214), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT17), .B(G131), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n195), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(G143), .A3(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(KEYINPUT87), .A3(KEYINPUT17), .A4(G131), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n294), .A2(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT73), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(KEYINPUT16), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n192), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n374), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n364), .A2(G131), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n362), .A2(new_n234), .A3(new_n363), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n366), .A2(new_n375), .A3(new_n377), .A4(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G113), .B(G122), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(new_n203), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n369), .A2(G146), .A3(new_n371), .ZN(new_n385));
  XNOR2_X1  g199(.A(G125), .B(G140), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n386), .A2(KEYINPUT75), .A3(new_n192), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT75), .B1(new_n386), .B2(new_n192), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n362), .A2(new_n363), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n364), .A2(KEYINPUT18), .A3(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n382), .A2(new_n384), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n384), .B1(new_n382), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n290), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G475), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n378), .A2(new_n380), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n369), .B2(new_n371), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n386), .A2(KEYINPUT19), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n192), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n377), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n393), .ZN(new_n406));
  INV_X1    g220(.A(new_n384), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n382), .A2(new_n384), .A3(new_n393), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n399), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT20), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT20), .B(new_n399), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n397), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT88), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT88), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n397), .B(new_n416), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G122), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G116), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n309), .A2(G122), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n211), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(G128), .A3(new_n195), .ZN(new_n425));
  XNOR2_X1  g239(.A(G128), .B(G143), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(G134), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n224), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n426), .B(new_n224), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n211), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n433), .A2(new_n420), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n431), .B(new_n432), .C1(new_n435), .C2(new_n211), .ZN(new_n436));
  INV_X1    g250(.A(G217), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n348), .A2(new_n437), .A3(G953), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n430), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n430), .B2(new_n436), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n283), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G952), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(G953), .ZN(new_n448));
  NAND2_X1  g262(.A1(G234), .A2(G237), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n283), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(G953), .A3(new_n449), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT90), .Z(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n352), .A2(new_n418), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n437), .B1(new_n283), .B2(G234), .ZN(new_n459));
  XOR2_X1   g273(.A(G119), .B(G128), .Z(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT24), .B(G110), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n307), .B2(G128), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n464), .B(new_n465), .C1(G119), .C2(new_n194), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n462), .B1(new_n466), .B2(G110), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n377), .B(new_n467), .C1(new_n388), .C2(new_n387), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n377), .A2(new_n375), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n460), .A2(new_n461), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(G110), .B2(new_n466), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT74), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n372), .A2(new_n192), .A3(new_n374), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n192), .B1(new_n372), .B2(new_n374), .ZN(new_n474));
  OAI211_X1 g288(.A(KEYINPUT74), .B(new_n471), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n468), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT22), .B(G137), .Z(new_n478));
  NAND3_X1  g292(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n480), .B(new_n481), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n468), .A3(new_n482), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT25), .B1(new_n490), .B2(new_n283), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n492), .B(new_n451), .C1(new_n484), .C2(new_n489), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n459), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n459), .A2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n226), .A2(new_n230), .A3(G131), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n234), .B1(new_n233), .B2(new_n235), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n250), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT30), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n228), .A2(KEYINPUT66), .A3(G134), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n227), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n202), .A2(new_n236), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n502), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n503), .B1(new_n502), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n315), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n315), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n513), .A3(new_n508), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n357), .A2(G210), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT26), .B(G101), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n499), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n298), .A2(new_n299), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n231), .B2(new_n236), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n202), .A2(new_n236), .A3(new_n507), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n315), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n525), .B2(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n514), .A2(new_n521), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n528), .A2(new_n519), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n534), .C1(KEYINPUT70), .C2(new_n532), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n527), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n519), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n538), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(new_n451), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n531), .B1(new_n526), .B2(new_n529), .ZN(new_n545));
  AOI211_X1 g359(.A(KEYINPUT68), .B(new_n521), .C1(new_n525), .C2(new_n514), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT30), .B1(new_n523), .B2(new_n524), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n509), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n514), .A2(new_n519), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n549), .A2(new_n315), .B1(new_n550), .B2(KEYINPUT67), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n514), .A2(new_n552), .A3(new_n519), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT31), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(KEYINPUT67), .ZN(new_n555));
  AND4_X1   g369(.A1(KEYINPUT31), .A2(new_n512), .A3(new_n555), .A4(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n547), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT69), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n512), .A2(new_n555), .A3(new_n553), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n551), .A2(KEYINPUT31), .A3(new_n553), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT69), .A3(new_n547), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n544), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n567), .ZN(new_n569));
  AOI211_X1 g383(.A(KEYINPUT32), .B(new_n569), .C1(new_n559), .C2(new_n565), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n543), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n458), .A2(new_n498), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n208), .B(KEYINPUT91), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G3));
  AND3_X1   g388(.A1(new_n564), .A2(KEYINPUT69), .A3(new_n547), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT69), .B1(new_n564), .B2(new_n547), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n283), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n577), .A2(G472), .B1(new_n566), .B2(new_n567), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n293), .A2(new_n351), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n497), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT92), .Z(new_n582));
  NAND3_X1  g396(.A1(new_n332), .A2(new_n333), .A3(new_n341), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n345), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n344), .B2(new_n584), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n442), .A2(new_n443), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT94), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n442), .A2(new_n589), .A3(new_n443), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n441), .B(KEYINPUT33), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(G478), .A3(new_n283), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n415), .A3(new_n417), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n455), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n582), .A2(new_n586), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT34), .B(G104), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G6));
  INV_X1    g413(.A(new_n414), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n446), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n455), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT95), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n582), .A2(new_n586), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G107), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G9));
  NOR2_X1   g420(.A1(new_n482), .A2(KEYINPUT36), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n477), .B(new_n607), .Z(new_n608));
  INV_X1    g422(.A(new_n495), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n494), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n456), .A2(new_n418), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n578), .A3(new_n352), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT37), .B(G110), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  XOR2_X1   g430(.A(new_n450), .B(KEYINPUT96), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G900), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n453), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n601), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n585), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n332), .A2(new_n341), .ZN(new_n623));
  INV_X1    g437(.A(new_n333), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n584), .A3(new_n583), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n611), .A2(new_n579), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n571), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n194), .ZN(G30));
  XOR2_X1   g444(.A(new_n620), .B(KEYINPUT39), .Z(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n579), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT40), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n519), .B1(new_n525), .B2(new_n514), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n551), .B2(new_n553), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n636), .B2(G902), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n568), .B2(new_n570), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n344), .B(KEYINPUT38), .Z(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n345), .A3(new_n611), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n415), .A2(new_n446), .A3(new_n417), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n634), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G143), .ZN(G45));
  INV_X1    g458(.A(new_n595), .ZN(new_n645));
  INV_X1    g459(.A(new_n620), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n567), .B1(new_n575), .B2(new_n576), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT32), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n566), .A2(new_n544), .A3(new_n567), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n647), .B1(new_n651), .B2(new_n543), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n628), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G146), .ZN(G48));
  AOI22_X1  g468(.A1(new_n649), .A2(new_n650), .B1(G472), .B2(new_n542), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n349), .A3(new_n284), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n627), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n655), .A2(new_n660), .A3(new_n497), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n596), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT41), .B(G113), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT97), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n662), .B(new_n664), .ZN(G15));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n603), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT98), .B(G116), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G18));
  NAND2_X1  g482(.A1(new_n613), .A2(new_n659), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n655), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n307), .ZN(G21));
  NAND2_X1  g485(.A1(new_n538), .A2(new_n539), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n564), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n567), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(KEYINPUT99), .A3(new_n567), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(G472), .B2(new_n577), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n410), .B(new_n411), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n416), .B1(new_n680), .B2(new_n397), .ZN(new_n681));
  INV_X1    g495(.A(new_n417), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n586), .A4(new_n446), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT100), .B1(new_n641), .B2(new_n627), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n658), .A2(new_n455), .ZN(new_n688));
  AND4_X1   g502(.A1(new_n498), .A2(new_n679), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n419), .ZN(G24));
  INV_X1    g504(.A(new_n611), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n595), .A2(new_n620), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n679), .A2(new_n691), .A3(new_n692), .A4(new_n659), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n695));
  NOR2_X1   g509(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n288), .A2(KEYINPUT101), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n287), .A2(new_n278), .A3(new_n699), .A4(new_n279), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n701), .A2(G469), .A3(new_n286), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n284), .A2(new_n292), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n349), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT102), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n344), .A2(new_n705), .A3(new_n345), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n625), .A2(new_n345), .A3(new_n583), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n704), .A2(new_n709), .A3(new_n497), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n697), .B1(new_n652), .B2(new_n710), .ZN(new_n711));
  AND4_X1   g525(.A1(new_n571), .A2(new_n710), .A3(new_n692), .A4(new_n697), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n695), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n571), .A2(new_n710), .A3(new_n692), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n696), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n652), .A2(new_n697), .A3(new_n710), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  NAND3_X1  g533(.A1(new_n571), .A2(new_n710), .A3(new_n621), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n415), .A2(new_n722), .A3(new_n417), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n722), .B1(new_n415), .B2(new_n417), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n594), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT43), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n418), .A2(new_n727), .A3(new_n594), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n578), .A3(new_n611), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT44), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n286), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n286), .B2(new_n288), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n282), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n291), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n284), .B1(new_n736), .B2(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n349), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(new_n632), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n709), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n732), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT106), .B(G137), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G39));
  AND2_X1   g558(.A1(new_n706), .A2(new_n708), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n655), .A2(new_n497), .A3(new_n692), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT107), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n739), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT47), .B(new_n349), .C1(new_n737), .C2(new_n738), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G140), .ZN(G42));
  NOR4_X1   g567(.A1(new_n611), .A2(new_n414), .A3(new_n446), .A4(new_n620), .ZN(new_n754));
  INV_X1    g568(.A(new_n579), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n571), .A2(new_n754), .A3(new_n755), .A4(new_n745), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n704), .A2(new_n709), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n679), .A2(new_n691), .A3(new_n692), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n758), .A3(new_n720), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n711), .A2(new_n712), .A3(new_n695), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT104), .B1(new_n715), .B2(new_n716), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR3_X1    g577(.A1(new_n344), .A2(new_n455), .A3(new_n346), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n683), .A3(new_n445), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n578), .A2(new_n765), .A3(new_n580), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n766), .B(new_n614), .C1(new_n655), .C2(new_n669), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n689), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n655), .A2(new_n457), .A3(new_n497), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT109), .B1(new_n764), .B2(new_n595), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n344), .A2(new_n455), .A3(new_n346), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n683), .A2(new_n771), .A3(new_n772), .A4(new_n594), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n770), .A2(new_n578), .A3(new_n580), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT110), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n661), .B1(new_n596), .B2(new_n603), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n572), .A2(new_n778), .A3(new_n774), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n768), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT111), .B1(new_n763), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n571), .B(new_n628), .C1(new_n621), .C2(new_n692), .ZN(new_n782));
  INV_X1    g596(.A(new_n704), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n494), .A2(new_n610), .A3(new_n646), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n494), .A2(new_n610), .A3(KEYINPUT112), .A4(new_n646), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n638), .A2(new_n687), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n782), .A2(new_n789), .A3(new_n693), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n782), .A2(new_n789), .A3(new_n693), .A4(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(KEYINPUT113), .A3(new_n791), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n768), .A2(new_n776), .A3(new_n777), .A4(new_n779), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n759), .B1(new_n713), .B2(new_n717), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n781), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n792), .A2(new_n794), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(new_n809), .A3(KEYINPUT54), .A4(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n805), .A2(new_n796), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n796), .B(new_n759), .C1(new_n716), .C2(new_n715), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n799), .A3(new_n797), .A4(new_n795), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n679), .A2(new_n498), .ZN(new_n816));
  INV_X1    g630(.A(new_n594), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT105), .B1(new_n681), .B2(new_n682), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n415), .A2(new_n722), .A3(new_n417), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n618), .B(new_n728), .C1(new_n820), .C2(new_n727), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n726), .A2(KEYINPUT115), .A3(new_n618), .A4(new_n728), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n816), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n659), .ZN(new_n826));
  INV_X1    g640(.A(new_n638), .ZN(new_n827));
  INV_X1    g641(.A(new_n284), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n656), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n349), .A3(new_n706), .A4(new_n708), .ZN(new_n830));
  INV_X1    g644(.A(new_n450), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n497), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n832), .A3(new_n645), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n826), .A2(KEYINPUT119), .A3(new_n448), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n660), .B(new_n816), .C1(new_n823), .C2(new_n824), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n448), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n830), .B1(new_n823), .B2(new_n824), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n655), .A2(new_n497), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT48), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT48), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n843), .A3(new_n840), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n834), .A2(new_n838), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n824), .ZN(new_n846));
  INV_X1    g660(.A(new_n816), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n639), .A2(new_n345), .A3(new_n658), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n418), .A2(new_n827), .A3(new_n832), .A4(new_n817), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n679), .A2(new_n691), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n839), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n816), .B(new_n709), .C1(new_n823), .C2(new_n824), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n829), .A2(new_n350), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n749), .A2(new_n750), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n853), .A2(new_n857), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n845), .A2(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n825), .A2(KEYINPUT50), .A3(new_n848), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT50), .B1(new_n825), .B2(new_n848), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n857), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n853), .A2(new_n869), .A3(new_n857), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n860), .B(KEYINPUT116), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n749), .A2(new_n871), .A3(new_n750), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n825), .A2(new_n872), .A3(new_n745), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n868), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n864), .B1(new_n876), .B2(new_n858), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n808), .A2(new_n810), .A3(new_n815), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n447), .A2(new_n354), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n829), .B(KEYINPUT49), .Z(new_n881));
  INV_X1    g695(.A(KEYINPUT108), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n498), .A2(new_n345), .A3(new_n351), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n639), .B(new_n881), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n638), .A2(new_n725), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n884), .B(new_n885), .C1(new_n882), .C2(new_n883), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n880), .A2(KEYINPUT120), .A3(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n354), .A2(G952), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n283), .B1(new_n811), .B2(new_n814), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(new_n624), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n337), .A2(new_n340), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(new_n338), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT55), .Z(new_n898));
  OAI21_X1  g712(.A(new_n893), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n895), .B2(new_n898), .ZN(G51));
  NAND2_X1  g714(.A1(new_n811), .A2(new_n814), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n902), .A2(new_n815), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n291), .B(KEYINPUT57), .Z(new_n904));
  OAI21_X1  g718(.A(new_n281), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n894), .A2(new_n733), .A3(new_n735), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n892), .B1(new_n905), .B2(new_n906), .ZN(G54));
  AND3_X1   g721(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n408), .A2(new_n409), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n893), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(G60));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT59), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n592), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n902), .B2(new_n815), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n915), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT121), .B1(new_n915), .B2(new_n892), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n808), .A2(new_n810), .A3(new_n815), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n592), .B1(new_n919), .B2(new_n913), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n920), .ZN(G63));
  XNOR2_X1  g735(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n437), .A2(new_n290), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n490), .B1(new_n901), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n892), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n901), .A2(new_n924), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n608), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n928), .A2(KEYINPUT123), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n930), .A3(new_n608), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT61), .B(new_n926), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  NOR3_X1   g750(.A1(new_n454), .A2(new_n301), .A3(new_n354), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n799), .B2(new_n354), .ZN(new_n938));
  INV_X1    g752(.A(G898), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n896), .B1(new_n939), .B2(G953), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n938), .B(new_n940), .Z(G69));
  OAI21_X1  g755(.A(G953), .B1(new_n188), .B2(new_n619), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n782), .A2(new_n693), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n643), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT62), .Z(new_n946));
  OAI21_X1  g760(.A(new_n595), .B1(new_n683), .B2(new_n445), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n840), .A2(new_n633), .A3(new_n745), .A4(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n742), .A3(new_n752), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n354), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n402), .A2(new_n403), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n549), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n953), .B2(KEYINPUT125), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(G900), .B2(G953), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n944), .A2(new_n720), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n840), .A2(new_n687), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n740), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n742), .A2(new_n959), .A3(new_n718), .A4(new_n752), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n960), .B2(G953), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n953), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n954), .B(new_n962), .ZN(G72));
  XOR2_X1   g777(.A(new_n515), .B(KEYINPUT127), .Z(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n949), .B2(new_n780), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n967), .A2(KEYINPUT126), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n966), .C1(new_n949), .C2(new_n780), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n519), .B(new_n964), .C1(new_n968), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n560), .B1(new_n515), .B2(new_n519), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n803), .A2(new_n806), .A3(new_n966), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n960), .B2(new_n780), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n964), .A2(new_n519), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n892), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n972), .A2(new_n974), .A3(new_n977), .ZN(G57));
endmodule


