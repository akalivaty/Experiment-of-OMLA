

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n533), .Z(n899) );
  NOR2_X2 U565 ( .A1(n549), .A2(n548), .ZN(G160) );
  NAND2_X1 U566 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U567 ( .A(n772), .B(n771), .ZN(n773) );
  NAND2_X1 U568 ( .A1(n531), .A2(n1023), .ZN(n775) );
  OR2_X1 U569 ( .A1(n783), .A2(n782), .ZN(n530) );
  OR2_X1 U570 ( .A1(n774), .A2(n783), .ZN(n531) );
  AND2_X1 U571 ( .A1(n784), .A2(n530), .ZN(n532) );
  NOR2_X1 U572 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U573 ( .A1(n713), .A2(n714), .ZN(n712) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n731) );
  XNOR2_X1 U575 ( .A(n732), .B(n731), .ZN(n733) );
  INV_X1 U576 ( .A(KEYINPUT64), .ZN(n771) );
  AND2_X1 U577 ( .A1(n785), .A2(n532), .ZN(n786) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n659) );
  XNOR2_X1 U579 ( .A(n534), .B(KEYINPUT66), .ZN(n891) );
  XOR2_X1 U580 ( .A(KEYINPUT65), .B(n553), .Z(n668) );
  NOR2_X1 U581 ( .A1(n542), .A2(n541), .ZN(G164) );
  NOR2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n899), .A2(G138), .ZN(n536) );
  INV_X1 U584 ( .A(G2105), .ZN(n538) );
  AND2_X1 U585 ( .A1(G2104), .A2(n538), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G102), .A2(n891), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U588 ( .A(n537), .B(KEYINPUT88), .ZN(n542) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U590 ( .A1(G114), .A2(n893), .ZN(n540) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n538), .ZN(n894) );
  NAND2_X1 U592 ( .A1(G126), .A2(n894), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n893), .A2(G113), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n891), .A2(G101), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n543), .Z(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U598 ( .A1(G137), .A2(n899), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G125), .A2(n894), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  INV_X1 U601 ( .A(G651), .ZN(n554) );
  NOR2_X1 U602 ( .A1(G543), .A2(n554), .ZN(n550) );
  XOR2_X1 U603 ( .A(KEYINPUT1), .B(n550), .Z(n672) );
  NAND2_X1 U604 ( .A1(G60), .A2(n672), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G85), .A2(n659), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n558) );
  XOR2_X1 U607 ( .A(KEYINPUT0), .B(G543), .Z(n665) );
  NOR2_X1 U608 ( .A1(G651), .A2(n665), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G47), .A2(n668), .ZN(n556) );
  NOR2_X1 U610 ( .A1(n665), .A2(n554), .ZN(n660) );
  NAND2_X1 U611 ( .A1(G72), .A2(n660), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  OR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(G290) );
  XNOR2_X1 U614 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U615 ( .A(G2446), .B(KEYINPUT106), .Z(n560) );
  XNOR2_X1 U616 ( .A(G2451), .B(G2430), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U618 ( .A(n561), .B(G2427), .Z(n563) );
  XNOR2_X1 U619 ( .A(G1341), .B(G1348), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n563), .B(n562), .ZN(n567) );
  XOR2_X1 U621 ( .A(G2443), .B(G2435), .Z(n565) );
  XNOR2_X1 U622 ( .A(G2438), .B(G2454), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U624 ( .A(n567), .B(n566), .Z(n568) );
  AND2_X1 U625 ( .A1(G14), .A2(n568), .ZN(G401) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U627 ( .A(G57), .ZN(G237) );
  NAND2_X1 U628 ( .A1(n668), .A2(G52), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n672), .A2(G64), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n576) );
  NAND2_X1 U631 ( .A1(G90), .A2(n659), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G77), .A2(n660), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT9), .B(n573), .ZN(n574) );
  XNOR2_X1 U635 ( .A(KEYINPUT67), .B(n574), .ZN(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(G171) );
  NAND2_X1 U637 ( .A1(G89), .A2(n659), .ZN(n577) );
  XNOR2_X1 U638 ( .A(n577), .B(KEYINPUT4), .ZN(n578) );
  XNOR2_X1 U639 ( .A(KEYINPUT72), .B(n578), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n660), .A2(G76), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT73), .B(n579), .Z(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U643 ( .A(n582), .B(KEYINPUT5), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G63), .A2(n672), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G51), .A2(n668), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n585), .Z(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U649 ( .A(n588), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n589) );
  XOR2_X1 U652 ( .A(n589), .B(KEYINPUT10), .Z(n925) );
  NAND2_X1 U653 ( .A1(n925), .A2(G567), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  NAND2_X1 U655 ( .A1(n672), .A2(G56), .ZN(n591) );
  XNOR2_X1 U656 ( .A(KEYINPUT14), .B(n591), .ZN(n597) );
  NAND2_X1 U657 ( .A1(n659), .A2(G81), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G68), .A2(n660), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(n595), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n598), .B(KEYINPUT69), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n668), .A2(G43), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n1028) );
  INV_X1 U666 ( .A(G860), .ZN(n639) );
  OR2_X1 U667 ( .A1(n1028), .A2(n639), .ZN(G153) );
  INV_X1 U668 ( .A(G171), .ZN(G301) );
  AND2_X1 U669 ( .A1(G301), .A2(G868), .ZN(n601) );
  XOR2_X1 U670 ( .A(KEYINPUT70), .B(n601), .Z(n611) );
  NAND2_X1 U671 ( .A1(G66), .A2(n672), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G92), .A2(n659), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U674 ( .A1(G54), .A2(n668), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G79), .A2(n660), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT15), .B(n608), .Z(n1009) );
  NOR2_X1 U679 ( .A1(n1009), .A2(G868), .ZN(n609) );
  XNOR2_X1 U680 ( .A(KEYINPUT71), .B(n609), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(G284) );
  NAND2_X1 U682 ( .A1(G65), .A2(n672), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G78), .A2(n660), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n659), .A2(G91), .ZN(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT68), .B(n614), .Z(n615) );
  NOR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n668), .A2(G53), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(G299) );
  XOR2_X1 U690 ( .A(KEYINPUT74), .B(G868), .Z(n619) );
  NOR2_X1 U691 ( .A1(G286), .A2(n619), .ZN(n621) );
  NOR2_X1 U692 ( .A1(G868), .A2(G299), .ZN(n620) );
  NOR2_X1 U693 ( .A1(n621), .A2(n620), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n639), .A2(G559), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n622), .A2(n1009), .ZN(n623) );
  XNOR2_X1 U696 ( .A(n623), .B(KEYINPUT16), .ZN(n624) );
  XOR2_X1 U697 ( .A(KEYINPUT75), .B(n624), .Z(G148) );
  NAND2_X1 U698 ( .A1(n1009), .A2(G868), .ZN(n625) );
  NOR2_X1 U699 ( .A1(G559), .A2(n625), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n626), .B(KEYINPUT76), .ZN(n628) );
  NOR2_X1 U701 ( .A1(n1028), .A2(G868), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U703 ( .A1(n893), .A2(G111), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G99), .A2(n891), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n894), .A2(G123), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT18), .ZN(n633) );
  NAND2_X1 U708 ( .A1(G135), .A2(n899), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U710 ( .A(KEYINPUT77), .B(n634), .Z(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n943) );
  XNOR2_X1 U712 ( .A(n943), .B(G2096), .ZN(n637) );
  INV_X1 U713 ( .A(G2100), .ZN(n848) );
  NAND2_X1 U714 ( .A1(n637), .A2(n848), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G559), .A2(n1009), .ZN(n638) );
  XOR2_X1 U716 ( .A(n1028), .B(n638), .Z(n681) );
  NAND2_X1 U717 ( .A1(n639), .A2(n681), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G67), .A2(n672), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G55), .A2(n668), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G93), .A2(n659), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G80), .A2(n660), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n684) );
  XOR2_X1 U725 ( .A(n646), .B(n684), .Z(G145) );
  NAND2_X1 U726 ( .A1(G61), .A2(n672), .ZN(n648) );
  NAND2_X1 U727 ( .A1(G86), .A2(n659), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G73), .A2(n660), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT2), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(KEYINPUT81), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n652), .A2(n651), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n668), .A2(G48), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n672), .A2(G62), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n655), .B(KEYINPUT82), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G50), .A2(n668), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U739 ( .A(KEYINPUT83), .B(n658), .ZN(n664) );
  NAND2_X1 U740 ( .A1(G88), .A2(n659), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G75), .A2(n660), .ZN(n661) );
  AND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(G303) );
  INV_X1 U744 ( .A(G303), .ZN(G166) );
  NAND2_X1 U745 ( .A1(n665), .A2(G87), .ZN(n666) );
  XNOR2_X1 U746 ( .A(KEYINPUT80), .B(n666), .ZN(n675) );
  NAND2_X1 U747 ( .A1(G651), .A2(G74), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(KEYINPUT78), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G49), .A2(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U752 ( .A(KEYINPUT79), .B(n673), .Z(n674) );
  NAND2_X1 U753 ( .A1(n675), .A2(n674), .ZN(G288) );
  XNOR2_X1 U754 ( .A(G305), .B(KEYINPUT19), .ZN(n677) );
  XOR2_X1 U755 ( .A(G299), .B(G166), .Z(n676) );
  XNOR2_X1 U756 ( .A(n677), .B(n676), .ZN(n678) );
  XOR2_X1 U757 ( .A(n684), .B(n678), .Z(n679) );
  XNOR2_X1 U758 ( .A(G290), .B(n679), .ZN(n680) );
  XNOR2_X1 U759 ( .A(n680), .B(G288), .ZN(n916) );
  XNOR2_X1 U760 ( .A(n916), .B(n681), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n682), .A2(G868), .ZN(n683) );
  XNOR2_X1 U762 ( .A(n683), .B(KEYINPUT84), .ZN(n686) );
  OR2_X1 U763 ( .A1(G868), .A2(n684), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U765 ( .A1(G2078), .A2(G2084), .ZN(n687) );
  XOR2_X1 U766 ( .A(KEYINPUT20), .B(n687), .Z(n688) );
  NAND2_X1 U767 ( .A1(G2090), .A2(n688), .ZN(n689) );
  XNOR2_X1 U768 ( .A(KEYINPUT21), .B(n689), .ZN(n690) );
  NAND2_X1 U769 ( .A1(n690), .A2(G2072), .ZN(G158) );
  NAND2_X1 U770 ( .A1(G120), .A2(G69), .ZN(n691) );
  NOR2_X1 U771 ( .A1(G237), .A2(n691), .ZN(n692) );
  XNOR2_X1 U772 ( .A(KEYINPUT86), .B(n692), .ZN(n693) );
  NAND2_X1 U773 ( .A1(n693), .A2(G108), .ZN(n846) );
  NAND2_X1 U774 ( .A1(G567), .A2(n846), .ZN(n694) );
  XNOR2_X1 U775 ( .A(n694), .B(KEYINPUT87), .ZN(n700) );
  NAND2_X1 U776 ( .A1(G132), .A2(G82), .ZN(n695) );
  XNOR2_X1 U777 ( .A(n695), .B(KEYINPUT85), .ZN(n696) );
  XNOR2_X1 U778 ( .A(KEYINPUT22), .B(n696), .ZN(n697) );
  NAND2_X1 U779 ( .A1(n697), .A2(G96), .ZN(n698) );
  OR2_X1 U780 ( .A1(G218), .A2(n698), .ZN(n847) );
  AND2_X1 U781 ( .A1(G2106), .A2(n847), .ZN(n699) );
  NOR2_X1 U782 ( .A1(n700), .A2(n699), .ZN(G319) );
  INV_X1 U783 ( .A(G319), .ZN(n702) );
  NAND2_X1 U784 ( .A1(G661), .A2(G483), .ZN(n701) );
  NOR2_X1 U785 ( .A1(n702), .A2(n701), .ZN(n845) );
  NAND2_X1 U786 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U787 ( .A1(G160), .A2(G40), .ZN(n787) );
  INV_X1 U788 ( .A(n787), .ZN(n703) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n788) );
  NAND2_X2 U790 ( .A1(n703), .A2(n788), .ZN(n747) );
  NAND2_X1 U791 ( .A1(G8), .A2(n747), .ZN(n783) );
  NOR2_X1 U792 ( .A1(G1966), .A2(n783), .ZN(n743) );
  INV_X1 U793 ( .A(KEYINPUT98), .ZN(n704) );
  XNOR2_X2 U794 ( .A(n747), .B(n704), .ZN(n719) );
  XNOR2_X1 U795 ( .A(KEYINPUT25), .B(G2078), .ZN(n967) );
  NAND2_X1 U796 ( .A1(n719), .A2(n967), .ZN(n706) );
  INV_X1 U797 ( .A(G1961), .ZN(n864) );
  NAND2_X1 U798 ( .A1(n864), .A2(n747), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n738) );
  AND2_X1 U800 ( .A1(n738), .A2(G171), .ZN(n707) );
  XNOR2_X1 U801 ( .A(KEYINPUT99), .B(n707), .ZN(n734) );
  NAND2_X1 U802 ( .A1(G2072), .A2(n719), .ZN(n708) );
  XNOR2_X1 U803 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  XOR2_X1 U804 ( .A(G1956), .B(KEYINPUT100), .Z(n977) );
  NOR2_X1 U805 ( .A1(n719), .A2(n977), .ZN(n709) );
  INV_X1 U806 ( .A(G299), .ZN(n714) );
  INV_X1 U807 ( .A(KEYINPUT28), .ZN(n711) );
  XNOR2_X1 U808 ( .A(n712), .B(n711), .ZN(n730) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n728) );
  INV_X1 U810 ( .A(G1996), .ZN(n957) );
  OR2_X1 U811 ( .A1(n747), .A2(n957), .ZN(n715) );
  XNOR2_X1 U812 ( .A(n715), .B(KEYINPUT26), .ZN(n718) );
  AND2_X1 U813 ( .A1(n747), .A2(G1341), .ZN(n716) );
  NOR2_X1 U814 ( .A1(n716), .A2(n1028), .ZN(n717) );
  AND2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n1009), .A2(n724), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n719), .A2(G2067), .ZN(n721) );
  NAND2_X1 U818 ( .A1(G1348), .A2(n747), .ZN(n720) );
  NAND2_X1 U819 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n726) );
  OR2_X1 U821 ( .A1(n1009), .A2(n724), .ZN(n725) );
  NAND2_X1 U822 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n756) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n747), .ZN(n744) );
  NOR2_X1 U826 ( .A1(n743), .A2(n744), .ZN(n735) );
  NAND2_X1 U827 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n736), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U830 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U832 ( .A(KEYINPUT31), .B(n741), .Z(n754) );
  AND2_X1 U833 ( .A1(n756), .A2(n754), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U835 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n763) );
  INV_X1 U837 ( .A(G8), .ZN(n753) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n783), .ZN(n749) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U841 ( .A1(n750), .A2(G303), .ZN(n751) );
  XOR2_X1 U842 ( .A(KEYINPUT101), .B(n751), .Z(n752) );
  OR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n757) );
  AND2_X1 U844 ( .A1(n754), .A2(n757), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n760) );
  INV_X1 U846 ( .A(n757), .ZN(n758) );
  OR2_X1 U847 ( .A1(n758), .A2(G286), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U849 ( .A(n761), .B(KEYINPUT32), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n779) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n764) );
  XOR2_X1 U852 ( .A(n764), .B(KEYINPUT102), .Z(n766) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  INV_X1 U854 ( .A(n1011), .ZN(n765) );
  AND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n779), .A2(n767), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n1018) );
  INV_X1 U858 ( .A(n783), .ZN(n768) );
  AND2_X1 U859 ( .A1(n1018), .A2(n768), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n772) );
  NOR2_X1 U861 ( .A1(KEYINPUT33), .A2(n773), .ZN(n776) );
  NAND2_X1 U862 ( .A1(n1011), .A2(KEYINPUT33), .ZN(n774) );
  XOR2_X1 U863 ( .A(G1981), .B(G305), .Z(n1023) );
  OR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n780), .A2(n783), .ZN(n784) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U870 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  XNOR2_X1 U871 ( .A(n786), .B(KEYINPUT103), .ZN(n826) );
  NOR2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n839) );
  INV_X1 U873 ( .A(n839), .ZN(n809) );
  NAND2_X1 U874 ( .A1(n899), .A2(G131), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT92), .B(n789), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G95), .A2(n891), .ZN(n790) );
  XOR2_X1 U877 ( .A(KEYINPUT91), .B(n790), .Z(n791) );
  NAND2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U879 ( .A(KEYINPUT93), .B(n793), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G107), .A2(n893), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G119), .A2(n894), .ZN(n794) );
  AND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n910) );
  XNOR2_X1 U884 ( .A(KEYINPUT94), .B(G1991), .ZN(n961) );
  NAND2_X1 U885 ( .A1(n910), .A2(n961), .ZN(n807) );
  NAND2_X1 U886 ( .A1(n891), .A2(G105), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT38), .ZN(n805) );
  NAND2_X1 U888 ( .A1(G117), .A2(n893), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G141), .A2(n899), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G129), .A2(n894), .ZN(n801) );
  XNOR2_X1 U892 ( .A(KEYINPUT95), .B(n801), .ZN(n802) );
  NOR2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n888) );
  NAND2_X1 U895 ( .A1(G1996), .A2(n888), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U897 ( .A(KEYINPUT96), .B(n808), .Z(n946) );
  NOR2_X1 U898 ( .A1(n809), .A2(n946), .ZN(n830) );
  XNOR2_X1 U899 ( .A(KEYINPUT97), .B(n830), .ZN(n824) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n1015) );
  NAND2_X1 U901 ( .A1(n839), .A2(n1015), .ZN(n810) );
  XNOR2_X1 U902 ( .A(KEYINPUT89), .B(n810), .ZN(n822) );
  NAND2_X1 U903 ( .A1(n899), .A2(G140), .ZN(n812) );
  NAND2_X1 U904 ( .A1(G104), .A2(n891), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT34), .B(n813), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G116), .A2(n893), .ZN(n815) );
  NAND2_X1 U908 ( .A1(G128), .A2(n894), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U910 ( .A(n816), .B(KEYINPUT35), .Z(n817) );
  NOR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U912 ( .A(KEYINPUT36), .B(n819), .Z(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT90), .B(n820), .Z(n904) );
  XNOR2_X1 U914 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NOR2_X1 U915 ( .A1(n904), .A2(n835), .ZN(n939) );
  NAND2_X1 U916 ( .A1(n939), .A2(n839), .ZN(n833) );
  INV_X1 U917 ( .A(n833), .ZN(n821) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n841) );
  NOR2_X1 U921 ( .A1(n888), .A2(G1996), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT104), .ZN(n931) );
  NOR2_X1 U923 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n961), .A2(n910), .ZN(n942) );
  NOR2_X1 U925 ( .A1(n828), .A2(n942), .ZN(n829) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n931), .A2(n831), .ZN(n832) );
  XNOR2_X1 U928 ( .A(KEYINPUT39), .B(n832), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n904), .A2(n835), .ZN(n936) );
  NAND2_X1 U931 ( .A1(n836), .A2(n936), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT105), .B(n837), .Z(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U935 ( .A(KEYINPUT40), .B(n842), .ZN(G329) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n925), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U942 ( .A(G132), .ZN(G219) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G108), .ZN(G238) );
  INV_X1 U945 ( .A(G96), .ZN(G221) );
  INV_X1 U946 ( .A(G82), .ZN(G220) );
  INV_X1 U947 ( .A(G69), .ZN(G235) );
  NOR2_X1 U948 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(n848), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U951 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT42), .B(G2090), .Z(n852) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(G2678), .B(G2096), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U959 ( .A(G2078), .B(G2084), .Z(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U961 ( .A(KEYINPUT110), .B(G1991), .Z(n860) );
  XOR2_X1 U962 ( .A(n957), .B(G1981), .Z(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n861), .B(KEYINPUT41), .Z(n863) );
  XNOR2_X1 U965 ( .A(G1956), .B(G1971), .ZN(n862) );
  XNOR2_X1 U966 ( .A(n863), .B(n862), .ZN(n868) );
  XOR2_X1 U967 ( .A(G1986), .B(G1976), .Z(n866) );
  XOR2_X1 U968 ( .A(G1966), .B(n864), .Z(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U970 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U971 ( .A(KEYINPUT109), .B(G2474), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n894), .ZN(n871) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(n871), .Z(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U976 ( .A1(G112), .A2(n893), .ZN(n873) );
  NAND2_X1 U977 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n899), .A2(G136), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G100), .A2(n891), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U982 ( .A1(G118), .A2(n893), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G130), .A2(n894), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U985 ( .A1(n899), .A2(G142), .ZN(n882) );
  NAND2_X1 U986 ( .A1(G106), .A2(n891), .ZN(n881) );
  NAND2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  XNOR2_X1 U989 ( .A(KEYINPUT112), .B(n884), .ZN(n885) );
  NOR2_X1 U990 ( .A1(n886), .A2(n885), .ZN(n890) );
  XOR2_X1 U991 ( .A(G160), .B(n943), .Z(n887) );
  XNOR2_X1 U992 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U993 ( .A(n890), .B(n889), .Z(n906) );
  NAND2_X1 U994 ( .A1(G103), .A2(n891), .ZN(n892) );
  XNOR2_X1 U995 ( .A(KEYINPUT113), .B(n892), .ZN(n903) );
  NAND2_X1 U996 ( .A1(G115), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G127), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n897), .B(KEYINPUT47), .ZN(n898) );
  XNOR2_X1 U1000 ( .A(n898), .B(KEYINPUT114), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n899), .A2(G139), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n926) );
  XNOR2_X1 U1004 ( .A(n904), .B(n926), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n912) );
  XOR2_X1 U1006 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n908) );
  XNOR2_X1 U1007 ( .A(G164), .B(G162), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1009 ( .A(n910), .B(n909), .Z(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1012 ( .A(n1028), .B(G286), .ZN(n915) );
  XOR2_X1 U1013 ( .A(G301), .B(n1009), .Z(n914) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(G401), .A2(n921), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT115), .B(n922), .Z(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n925), .ZN(G223) );
  XOR2_X1 U1026 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1029 ( .A(KEYINPUT50), .B(n929), .Z(n935) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n932), .Z(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT117), .B(n933), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(G160), .B(G2084), .ZN(n937) );
  NAND2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n948) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1040 ( .A(n944), .B(KEYINPUT116), .ZN(n945) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT52), .B(n949), .ZN(n950) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n975) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n975), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n951), .A2(G29), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n952), .ZN(n1007) );
  XOR2_X1 U1048 ( .A(G2090), .B(G35), .Z(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(G34), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n954), .B(G2084), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n973) );
  XOR2_X1 U1053 ( .A(n957), .B(G32), .Z(n959) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n966) );
  XOR2_X1 U1056 ( .A(G2067), .B(G26), .Z(n960) );
  NAND2_X1 U1057 ( .A1(n960), .A2(G28), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT119), .B(n961), .Z(n962) );
  XNOR2_X1 U1059 ( .A(G25), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1062 ( .A(G27), .B(n967), .Z(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT120), .B(n970), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(G29), .A2(n976), .ZN(n1005) );
  XOR2_X1 U1069 ( .A(G5), .B(G1961), .Z(n992) );
  XNOR2_X1 U1070 ( .A(n977), .B(G20), .ZN(n986) );
  XOR2_X1 U1071 ( .A(G1341), .B(G19), .Z(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G4), .Z(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT125), .B(n978), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n979), .B(G1348), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(G1981), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G6), .B(n982), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT60), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G21), .B(G1966), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT126), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1088 ( .A(G1986), .B(G24), .Z(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT58), .B(n997), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XOR2_X1 U1092 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n1000) );
  XNOR2_X1 U1093 ( .A(n1001), .B(n1000), .ZN(n1002) );
  INV_X1 U1094 ( .A(G16), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1008), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(G11), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1035) );
  XNOR2_X1 U1099 ( .A(n1008), .B(KEYINPUT56), .ZN(n1033) );
  XOR2_X1 U1100 ( .A(G1348), .B(n1009), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(G299), .B(G1956), .Z(n1013) );
  XOR2_X1 U1103 ( .A(G301), .B(G1961), .Z(n1012) );
  NAND2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(G303), .B(G1971), .Z(n1019) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(KEYINPUT122), .B(n1022), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(G1966), .B(G168), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT57), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(G1341), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT123), .B(n1031), .Z(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1120 ( .A(n1036), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

