//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  INV_X1    g004(.A(G15gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G22gat), .ZN(new_n207));
  INV_X1    g006(.A(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G15gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n205), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(G8gat), .B1(new_n203), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n202), .A2(new_n205), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n212), .B(new_n213), .C1(G1gat), .C2(new_n202), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT82), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT82), .B1(new_n211), .B2(new_n214), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT17), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(G43gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G43gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(G43gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(G50gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT15), .ZN(new_n227));
  NOR2_X1   g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT14), .ZN(new_n229));
  INV_X1    g028(.A(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(G29gat), .A2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT14), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n224), .A2(new_n227), .A3(new_n229), .A4(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT15), .ZN(new_n235));
  INV_X1    g034(.A(new_n229), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n228), .B1(KEYINPUT14), .B2(new_n231), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT81), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n218), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n234), .B2(new_n238), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT15), .B1(new_n225), .B2(new_n226), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n237), .A2(new_n236), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT81), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT17), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n217), .B1(new_n243), .B2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT84), .B1(new_n211), .B2(new_n214), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT84), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n252), .B(new_n253), .C1(new_n244), .C2(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(G229gat), .A2(G233gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT83), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT85), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT85), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n250), .A2(new_n261), .A3(new_n254), .A4(new_n257), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT80), .B(G197gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G113gat), .B(G141gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT11), .B(G169gat), .Z(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT12), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n254), .A4(new_n257), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n244), .A2(new_n248), .ZN(new_n271));
  INV_X1    g070(.A(new_n253), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(new_n251), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n256), .B(KEYINPUT13), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n263), .A2(new_n269), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n270), .A2(new_n276), .A3(KEYINPUT87), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT87), .B1(new_n270), .B2(new_n276), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n263), .A2(KEYINPUT86), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n259), .A2(new_n284), .A3(new_n260), .A4(new_n262), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n269), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT89), .B1(G85gat), .B2(G92gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI211_X1 g092(.A(KEYINPUT89), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G85gat), .ZN(new_n296));
  AND2_X1   g095(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT91), .ZN(new_n300));
  INV_X1    g099(.A(G99gat), .ZN(new_n301));
  INV_X1    g100(.A(G106gat), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT8), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n299), .B2(new_n303), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G99gat), .B(G106gat), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT94), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n306), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G57gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G64gat), .ZN(new_n312));
  INV_X1    g111(.A(G64gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G57gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT9), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G71gat), .A2(G78gat), .ZN(new_n316));
  OR2_X1    g115(.A1(G71gat), .A2(G78gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT9), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT88), .B1(new_n313), .B2(G57gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n311), .A3(G64gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(new_n312), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n306), .A2(new_n307), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n295), .B(new_n308), .C1(new_n304), .C2(new_n305), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT93), .B1(new_n331), .B2(new_n326), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n333), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n289), .B(new_n328), .C1(new_n332), .C2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n327), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G230gat), .A2(G233gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n332), .A2(new_n334), .ZN(new_n341));
  INV_X1    g140(.A(new_n328), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G120gat), .B(G148gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G176gat), .ZN(new_n345));
  INV_X1    g144(.A(G204gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n343), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n340), .B1(new_n335), .B2(new_n336), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n352), .A3(KEYINPUT96), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT96), .B1(new_n349), .B2(new_n352), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT40), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(G120gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G113gat), .ZN(new_n365));
  INV_X1    g164(.A(G113gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G120gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT1), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G127gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G134gat), .ZN(new_n370));
  INV_X1    g169(.A(G127gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n368), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n376));
  INV_X1    g175(.A(G141gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(G148gat), .ZN(new_n378));
  INV_X1    g177(.A(G148gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G141gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n376), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382));
  INV_X1    g181(.A(G155gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n385), .B2(KEYINPUT2), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n379), .A2(KEYINPUT70), .A3(G141gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT70), .B1(new_n379), .B2(G141gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT73), .B1(new_n375), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n370), .A4(new_n374), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT75), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n375), .A2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n398), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n393), .A2(new_n396), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT75), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n375), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n408));
  XOR2_X1   g207(.A(KEYINPUT72), .B(KEYINPUT3), .Z(new_n409));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n363), .B1(new_n415), .B2(KEYINPUT39), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n405), .B2(new_n411), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT39), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n397), .B1(new_n392), .B2(new_n407), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n413), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n358), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n400), .B2(KEYINPUT4), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n411), .B(new_n424), .C1(new_n397), .C2(KEYINPUT4), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(KEYINPUT5), .C1(new_n413), .C2(new_n419), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n405), .A2(new_n411), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n363), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G183gat), .ZN(new_n432));
  INV_X1    g231(.A(G190gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(KEYINPUT24), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(KEYINPUT24), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT23), .ZN(new_n440));
  OAI22_X1  g239(.A1(new_n439), .A2(new_n440), .B1(G169gat), .B2(G176gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT25), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT64), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n447), .B2(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n436), .A2(new_n437), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(KEYINPUT64), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n442), .B(new_n440), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT66), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n442), .B2(new_n439), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT26), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT65), .B1(new_n455), .B2(KEYINPUT66), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n454), .A2(new_n455), .B1(new_n442), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n435), .B1(new_n457), .B2(new_n445), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT27), .B(G183gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n433), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT28), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n446), .B(new_n452), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G197gat), .B(G204gat), .ZN(new_n467));
  INV_X1    g266(.A(G211gat), .ZN(new_n468));
  INV_X1    g267(.A(G218gat), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(KEYINPUT22), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G211gat), .B(G218gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OR3_X1    g273(.A1(new_n464), .A2(new_n466), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(new_n313), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n477), .B(G92gat), .Z(new_n478));
  OR2_X1    g277(.A1(new_n464), .A2(KEYINPUT68), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n475), .B(new_n478), .C1(new_n481), .C2(new_n473), .ZN(new_n482));
  INV_X1    g281(.A(new_n478), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  INV_X1    g283(.A(new_n475), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n486), .A3(KEYINPUT30), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n475), .B1(new_n481), .B2(new_n473), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n483), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n415), .A2(KEYINPUT39), .A3(new_n420), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n430), .B1(new_n417), .B2(new_n418), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(KEYINPUT40), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n423), .A2(new_n431), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n465), .A3(new_n392), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n394), .B2(new_n409), .ZN(new_n497));
  OAI221_X1 g296(.A(new_n496), .B1(new_n394), .B2(new_n409), .C1(new_n497), .C2(new_n474), .ZN(new_n498));
  INV_X1    g297(.A(G228gat), .ZN(new_n499));
  INV_X1    g298(.A(G233gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n497), .A2(new_n474), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n499), .A2(new_n500), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n408), .A3(new_n503), .A4(new_n496), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G22gat), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n501), .A2(new_n504), .A3(new_n208), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT78), .ZN(new_n508));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(new_n222), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT76), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n511), .B(KEYINPUT31), .Z(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n501), .A2(new_n504), .A3(new_n208), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n208), .B1(new_n501), .B2(new_n504), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT78), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n506), .A2(new_n514), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(new_n512), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n519), .B(new_n512), .C1(new_n507), .C2(new_n515), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n481), .A2(new_n473), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n474), .B1(new_n464), .B2(new_n466), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT37), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT37), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n483), .B1(new_n488), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(KEYINPUT79), .A3(KEYINPUT37), .A4(new_n526), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT38), .B1(new_n488), .B2(new_n483), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT38), .ZN(new_n535));
  INV_X1    g334(.A(new_n488), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(KEYINPUT37), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n533), .A2(new_n534), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n426), .A2(new_n428), .A3(new_n363), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n431), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n429), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n495), .B(new_n524), .C1(new_n538), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n462), .A2(new_n375), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n462), .A2(new_n375), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G227gat), .A2(G233gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G43gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G71gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(new_n301), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT33), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(KEYINPUT32), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n549), .B1(new_n546), .B2(new_n547), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n554), .B1(new_n557), .B2(KEYINPUT33), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT32), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n556), .B(KEYINPUT67), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n549), .A3(new_n547), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT34), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n551), .A2(KEYINPUT32), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n551), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT67), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .A4(new_n554), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n561), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n563), .B1(new_n561), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n545), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n561), .A2(new_n568), .ZN(new_n573));
  INV_X1    g372(.A(new_n563), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(KEYINPUT36), .A3(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n491), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n543), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n524), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n544), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n570), .A2(new_n571), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(new_n524), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n543), .A4(new_n578), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n524), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT35), .B1(new_n579), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n288), .B(new_n357), .C1(new_n582), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n326), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n371), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n252), .A2(new_n253), .B1(KEYINPUT21), .B2(new_n327), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(G155gat), .B(G183gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n468), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n604), .A2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n331), .A2(new_n271), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n331), .B1(new_n243), .B2(new_n249), .ZN(new_n612));
  NAND3_X1  g411(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n614), .A2(G134gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(G134gat), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  AND3_X1   g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n384), .ZN(new_n621));
  OR3_X1    g420(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n618), .B2(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n591), .B1(new_n610), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(KEYINPUT92), .A3(new_n609), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n590), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n543), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT97), .B(G1gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(G1324gat));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n634));
  INV_X1    g433(.A(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n491), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n636), .B2(KEYINPUT98), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n491), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(G8gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(G1325gat));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n570), .A2(new_n571), .A3(new_n545), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT36), .B1(new_n575), .B2(new_n569), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n572), .A2(new_n576), .A3(KEYINPUT100), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n630), .A2(new_n206), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n583), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n650), .B1(new_n206), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n630), .A2(new_n524), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  NAND3_X1  g454(.A1(new_n544), .A2(new_n649), .A3(new_n581), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n589), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n624), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT102), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n626), .B1(new_n582), .B2(new_n589), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n626), .B1(new_n656), .B2(new_n589), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n658), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n357), .A2(new_n609), .A3(new_n288), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n543), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n661), .A2(new_n667), .ZN(new_n672));
  INV_X1    g471(.A(G29gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n543), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT45), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(G1328gat));
  OAI21_X1  g476(.A(G36gat), .B1(new_n670), .B2(new_n578), .ZN(new_n678));
  INV_X1    g477(.A(G36gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n679), .A3(new_n491), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT46), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(G1329gat));
  INV_X1    g481(.A(new_n649), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n669), .A2(G43gat), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n672), .A2(new_n583), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(G43gat), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n580), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n580), .A2(new_n222), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n688), .A2(G50gat), .B1(new_n672), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g491(.A1(new_n629), .A2(new_n657), .A3(new_n288), .A4(new_n357), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n674), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G57gat), .ZN(G1332gat));
  INV_X1    g494(.A(KEYINPUT49), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n693), .B(new_n491), .C1(new_n696), .C2(new_n313), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT103), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n313), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1333gat));
  AOI21_X1  g499(.A(G71gat), .B1(new_n693), .B2(new_n583), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n683), .A2(G71gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g503(.A1(new_n693), .A2(new_n580), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g505(.A1(new_n286), .A2(new_n287), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n278), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n609), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n666), .A2(new_n357), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710), .B2(new_n543), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n663), .A2(KEYINPUT51), .A3(new_n709), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT51), .B1(new_n663), .B2(new_n709), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n296), .A3(new_n357), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n717), .B2(new_n543), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1336gat));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n710), .A2(new_n578), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n297), .A2(new_n298), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n712), .A2(new_n713), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n578), .A2(G92gat), .A3(new_n356), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n722), .A2(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n725), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  OAI22_X1  g528(.A1(new_n721), .A2(new_n726), .B1(new_n727), .B2(new_n729), .ZN(G1337gat));
  OAI21_X1  g529(.A(G99gat), .B1(new_n710), .B2(new_n649), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n301), .A3(new_n583), .A4(new_n357), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1338gat));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n524), .A2(new_n356), .A3(G106gat), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT53), .B1(new_n716), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n666), .A2(new_n580), .A3(new_n357), .A4(new_n709), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G106gat), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n735), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n738), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n737), .A2(G106gat), .B1(new_n724), .B2(new_n735), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n744), .B(KEYINPUT106), .C1(new_n745), .C2(new_n740), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1339gat));
  NAND4_X1  g546(.A1(new_n625), .A2(new_n627), .A3(new_n288), .A4(new_n356), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT54), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n337), .A2(new_n749), .A3(new_n338), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n335), .A2(new_n340), .A3(new_n336), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT54), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n347), .B(new_n750), .C1(new_n752), .C2(new_n351), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n349), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n339), .A2(KEYINPUT54), .A3(new_n751), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n348), .B1(new_n351), .B2(new_n749), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT55), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n288), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n274), .A2(new_n275), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n257), .B1(new_n250), .B2(new_n254), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n268), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n278), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n355), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(new_n353), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT107), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n756), .A2(KEYINPUT55), .A3(new_n757), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n349), .ZN(new_n768));
  INV_X1    g567(.A(new_n758), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n708), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n278), .B(new_n762), .C1(new_n354), .C2(new_n355), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n766), .A2(new_n626), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n758), .A2(new_n763), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n624), .A2(new_n776), .A3(new_n768), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n610), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n775), .B1(new_n774), .B2(new_n777), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n748), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n584), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n674), .A3(new_n578), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n288), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n674), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n782), .A2(new_n787), .A3(new_n674), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n578), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n708), .A2(new_n366), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(G1340gat));
  OAI21_X1  g590(.A(G120gat), .B1(new_n783), .B2(new_n356), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n357), .A2(new_n364), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n789), .B2(new_n793), .ZN(G1341gat));
  OAI21_X1  g593(.A(G127gat), .B1(new_n783), .B2(new_n610), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n609), .A2(new_n371), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1342gat));
  NOR2_X1   g598(.A1(new_n626), .A2(G134gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n786), .A2(new_n578), .A3(new_n788), .A4(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n801), .A2(KEYINPUT56), .ZN(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n783), .B2(new_n626), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(KEYINPUT56), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n781), .A2(new_n580), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n649), .A2(new_n674), .A3(new_n578), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n288), .A2(G141gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(KEYINPUT115), .B2(new_n810), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(KEYINPUT58), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n807), .B(KEYINPUT111), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT57), .B1(new_n781), .B2(new_n580), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n580), .A2(KEYINPUT57), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n624), .B1(new_n770), .B2(new_n772), .ZN(new_n819));
  INV_X1    g618(.A(new_n777), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT112), .B(new_n610), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n748), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n626), .B1(new_n759), .B2(new_n765), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n777), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT112), .B1(new_n824), .B2(new_n610), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n818), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n828), .B(new_n818), .C1(new_n822), .C2(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n708), .B(new_n815), .C1(new_n816), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT116), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n814), .B1(new_n832), .B2(new_n377), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n815), .B1(new_n816), .B2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT114), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n815), .C1(new_n816), .C2(new_n830), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n708), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n813), .B1(new_n839), .B2(G141gat), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(G1344gat));
  NAND3_X1  g641(.A1(new_n808), .A2(new_n379), .A3(new_n357), .ZN(new_n843));
  AOI211_X1 g642(.A(KEYINPUT59), .B(new_n379), .C1(new_n838), .C2(new_n357), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n610), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n748), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n847), .B2(new_n580), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT118), .Z(new_n849));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n806), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n781), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n580), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n357), .A3(new_n815), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n845), .B1(new_n855), .B2(G148gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n843), .B1(new_n844), .B2(new_n856), .ZN(G1345gat));
  NAND3_X1  g656(.A1(new_n808), .A2(new_n383), .A3(new_n609), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n610), .B1(new_n835), .B2(new_n837), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n383), .ZN(G1346gat));
  AOI21_X1  g659(.A(new_n384), .B1(new_n838), .B2(new_n624), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n808), .A2(new_n384), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n626), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT119), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n626), .B1(new_n835), .B2(new_n837), .ZN(new_n866));
  OAI221_X1 g665(.A(new_n865), .B1(new_n626), .B2(new_n862), .C1(new_n866), .C2(new_n384), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(G1347gat));
  NOR2_X1   g667(.A1(new_n674), .A2(new_n578), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n782), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n708), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(G169gat), .ZN(G1348gat));
  NOR2_X1   g672(.A1(new_n870), .A2(new_n356), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT120), .B(G176gat), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n874), .B(new_n875), .ZN(G1349gat));
  OAI22_X1  g675(.A1(new_n870), .A2(new_n610), .B1(KEYINPUT121), .B2(new_n432), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n459), .B1(KEYINPUT121), .B2(G183gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n871), .A2(new_n609), .A3(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n877), .B(new_n879), .C1(KEYINPUT122), .C2(KEYINPUT60), .ZN(new_n880));
  NAND2_X1  g679(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1350gat));
  NAND4_X1  g681(.A1(new_n781), .A2(new_n624), .A3(new_n584), .A4(new_n869), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G190gat), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n884), .A2(KEYINPUT124), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(KEYINPUT124), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(KEYINPUT61), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n883), .A2(G190gat), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n884), .A2(KEYINPUT124), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT125), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1351gat));
  NAND3_X1  g696(.A1(new_n649), .A2(new_n491), .A3(new_n580), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT126), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n781), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(G197gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n674), .B1(new_n898), .B2(KEYINPUT126), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n900), .A2(new_n901), .A3(new_n708), .A4(new_n902), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n649), .A2(new_n869), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n854), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n708), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n901), .ZN(G1352gat));
  NAND4_X1  g706(.A1(new_n900), .A2(new_n346), .A3(new_n357), .A4(new_n902), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n854), .A2(new_n357), .A3(new_n904), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n912), .B(new_n913), .C1(new_n914), .C2(new_n346), .ZN(G1353gat));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n468), .A3(new_n609), .A4(new_n902), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n854), .A2(new_n609), .A3(new_n904), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n917), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n918));
  AOI21_X1  g717(.A(KEYINPUT63), .B1(new_n917), .B2(G211gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1354gat));
  NOR2_X1   g719(.A1(new_n626), .A2(new_n469), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n900), .A2(new_n624), .A3(new_n902), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n905), .A2(new_n921), .B1(new_n922), .B2(new_n469), .ZN(G1355gat));
endmodule


