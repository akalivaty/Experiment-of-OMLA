//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n229));
  OR2_X1    g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n214), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT66), .B(G50), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n256), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n255), .A2(KEYINPUT69), .A3(new_n257), .A4(new_n258), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G226), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G222), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G223), .A3(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n271), .B(new_n273), .C1(new_n274), .C2(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n253), .A2(new_n254), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n258), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n255), .A2(new_n278), .A3(G274), .A4(new_n257), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n265), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G190), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n254), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n208), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G50), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(G50), .B2(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n209), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT8), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G58), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n209), .A2(new_n267), .ZN(new_n295));
  INV_X1    g0095(.A(G150), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n209), .B1(new_n201), .B2(new_n202), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n294), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(new_n254), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n289), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n289), .B(KEYINPUT73), .C1(new_n301), .C2(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(KEYINPUT9), .A3(new_n305), .ZN(new_n309));
  INV_X1    g0109(.A(new_n279), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n310), .B1(new_n275), .B2(new_n276), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n263), .B2(new_n264), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n282), .A2(new_n308), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n309), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n282), .A4(new_n308), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n281), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n302), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n283), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n216), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G20), .A2(G33), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n274), .B2(new_n290), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT11), .A3(new_n300), .ZN(new_n332));
  INV_X1    g0132(.A(new_n285), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G68), .A3(new_n286), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT11), .B1(new_n331), .B2(new_n300), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n217), .B1(new_n261), .B2(new_n262), .ZN(new_n340));
  MUX2_X1   g0140(.A(G226), .B(G232), .S(G1698), .Z(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n272), .B1(G33), .B2(G97), .ZN(new_n342));
  INV_X1    g0142(.A(new_n276), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n279), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n340), .A2(KEYINPUT13), .A3(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n339), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n340), .A2(new_n344), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(G179), .A3(new_n345), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n345), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n339), .B1(new_n354), .B2(G169), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n338), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n346), .A2(new_n347), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n338), .B1(new_n357), .B2(G190), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT74), .B1(new_n354), .B2(G200), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT74), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  AOI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n351), .C2(new_n345), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n358), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT16), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n247), .A2(new_n216), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n366), .B2(new_n201), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n329), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n268), .A2(new_n209), .A3(new_n269), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT7), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n269), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n216), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI211_X1 g0177(.A(KEYINPUT75), .B(new_n216), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n375), .A2(new_n369), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n301), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n255), .A2(G274), .A3(new_n257), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n267), .A2(new_n218), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n264), .A2(G1698), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G223), .B2(G1698), .ZN(new_n387));
  AND2_X1   g0187(.A1(KEYINPUT3), .A2(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT3), .A2(G33), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n383), .A2(new_n278), .B1(new_n391), .B2(new_n276), .ZN(new_n392));
  INV_X1    g0192(.A(G190), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n255), .A2(G232), .A3(new_n257), .A4(new_n258), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n392), .A2(KEYINPUT78), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT78), .ZN(new_n396));
  NOR2_X1   g0196(.A1(G223), .A2(G1698), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n264), .B2(G1698), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n384), .B1(new_n398), .B2(new_n272), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n279), .B(new_n394), .C1(new_n399), .C2(new_n343), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(new_n361), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(G190), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n395), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n291), .A2(new_n293), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n286), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n405), .A2(new_n285), .B1(new_n283), .B2(new_n404), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT76), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n382), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n400), .A2(G169), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n391), .A2(new_n276), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(G179), .A3(new_n279), .A4(new_n394), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT77), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n413), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n408), .B1(new_n379), .B2(new_n381), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT18), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT7), .B1(new_n390), .B2(new_n209), .ZN(new_n423));
  INV_X1    g0223(.A(new_n374), .ZN(new_n424));
  OAI21_X1  g0224(.A(G68), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n369), .B1(new_n425), .B2(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n375), .A2(new_n376), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(new_n370), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n300), .B1(new_n429), .B2(new_n365), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n409), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n417), .A4(new_n419), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n412), .A2(new_n422), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n270), .A2(G232), .B1(new_n390), .B2(G107), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n310), .B1(new_n438), .B2(new_n276), .ZN(new_n439));
  INV_X1    g0239(.A(G244), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n320), .C1(new_n440), .C2(new_n263), .ZN(new_n441));
  INV_X1    g0241(.A(new_n439), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n263), .A2(new_n440), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n444), .B2(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n333), .A2(G77), .A3(new_n286), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT72), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G77), .B2(new_n283), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT70), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n404), .B(new_n449), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n450), .A2(new_n295), .B1(new_n209), .B2(new_n274), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT71), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n290), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI221_X1 g0257(.A(KEYINPUT71), .B1(new_n209), .B2(new_n274), .C1(new_n450), .C2(new_n295), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n448), .B1(new_n459), .B2(new_n300), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n445), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n444), .A2(G190), .ZN(new_n462));
  OAI21_X1  g0262(.A(G200), .B1(new_n442), .B2(new_n443), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n325), .A2(new_n364), .A3(new_n435), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(KEYINPUT83), .A3(new_n208), .A4(G45), .ZN(new_n470));
  INV_X1    g0270(.A(G41), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n208), .B(G45), .C1(new_n471), .C2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n472), .A2(new_n473), .B1(KEYINPUT5), .B2(new_n471), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n383), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n471), .A2(KEYINPUT5), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n255), .A2(new_n257), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(G264), .ZN(new_n480));
  OAI211_X1 g0280(.A(G257), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n481));
  INV_X1    g0281(.A(G1698), .ZN(new_n482));
  OAI211_X1 g0282(.A(G250), .B(new_n482), .C1(new_n388), .C2(new_n389), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G294), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n276), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n475), .A2(new_n480), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G169), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n475), .A2(new_n480), .A3(G179), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT86), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n209), .B2(G107), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n267), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n493), .A2(new_n495), .B1(new_n497), .B2(new_n209), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n209), .B(G87), .C1(new_n388), .C2(new_n389), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n499), .B(KEYINPUT22), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n506), .B2(new_n498), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n300), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT25), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n283), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n283), .A2(new_n509), .A3(G107), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n208), .A2(G33), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n283), .A2(new_n513), .A3(new_n254), .A4(new_n284), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n511), .A2(new_n512), .B1(new_n494), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n488), .A2(new_n518), .A3(new_n489), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n491), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT88), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n480), .A2(new_n486), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(KEYINPUT87), .A3(new_n393), .A4(new_n475), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT87), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n487), .B2(new_n361), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n487), .A2(G190), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n502), .A2(new_n503), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n506), .A2(new_n498), .A3(new_n505), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n515), .B1(new_n530), .B2(new_n300), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n520), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n521), .B1(new_n520), .B2(new_n532), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(G107), .B1(new_n423), .B2(new_n424), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  AND2_X1   g0337(.A1(G97), .A2(G107), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n205), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n494), .A2(KEYINPUT6), .A3(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT79), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n295), .B2(new_n274), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n329), .A2(KEYINPUT79), .A3(G77), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n541), .A2(G20), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n301), .B1(new_n536), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n544), .ZN(new_n548));
  INV_X1    g0348(.A(new_n540), .ZN(new_n549));
  XNOR2_X1  g0349(.A(G97), .B(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n537), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n551), .B2(new_n209), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n494), .B1(new_n373), .B2(new_n374), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT80), .B(new_n300), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n514), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(G97), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n283), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n555), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT4), .B1(new_n270), .B2(G244), .ZN(new_n564));
  AND2_X1   g0364(.A1(KEYINPUT4), .A2(G244), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n482), .B(new_n565), .C1(new_n388), .C2(new_n389), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G250), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n272), .A2(new_n572), .A3(G250), .A4(G1698), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n343), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n478), .A2(new_n479), .A3(G257), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n475), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n575), .A2(new_n577), .A3(G190), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n255), .A2(new_n257), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n470), .B2(new_n474), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n476), .A2(new_n470), .A3(new_n477), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(G257), .B1(new_n383), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(new_n482), .C1(new_n388), .C2(new_n389), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n567), .B(new_n566), .C1(new_n584), .C2(KEYINPUT4), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n571), .A2(new_n573), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n276), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(G200), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n547), .B(new_n563), .C1(new_n578), .C2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n322), .B1(new_n575), .B2(new_n577), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n582), .A2(new_n587), .A3(new_n320), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n554), .A2(new_n562), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n590), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G45), .ZN(new_n595));
  OR3_X1    g0395(.A1(new_n595), .A2(G1), .A3(G274), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n219), .B1(new_n595), .B2(G1), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n255), .A2(new_n596), .A3(new_n257), .A4(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G238), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n440), .B2(G1698), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n497), .B1(new_n600), .B2(new_n272), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(new_n343), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G200), .ZN(new_n603));
  NAND3_X1  g0403(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n209), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n206), .B2(G87), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n209), .B(G68), .C1(new_n388), .C2(new_n389), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n290), .B2(new_n556), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n300), .B1(new_n326), .B2(new_n454), .ZN(new_n611));
  INV_X1    g0411(.A(new_n514), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G87), .ZN(new_n613));
  OAI211_X1 g0413(.A(G190), .B(new_n598), .C1(new_n601), .C2(new_n343), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n603), .A2(new_n611), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n300), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n612), .A2(new_n455), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n454), .A2(new_n326), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n602), .A2(new_n322), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n320), .B(new_n598), .C1(new_n601), .C2(new_n343), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n589), .A2(new_n594), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(G264), .B(G1698), .C1(new_n388), .C2(new_n389), .ZN(new_n627));
  OAI211_X1 g0427(.A(G257), .B(new_n482), .C1(new_n388), .C2(new_n389), .ZN(new_n628));
  INV_X1    g0428(.A(G303), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n272), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n276), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n478), .A2(new_n479), .A3(G270), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n475), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n567), .B(new_n209), .C1(G33), .C2(new_n556), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n496), .A2(G20), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(new_n300), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n300), .A4(new_n635), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n283), .A2(new_n496), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n612), .B2(new_n496), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n322), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT21), .B1(new_n633), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n475), .A2(new_n632), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n642), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n646), .A2(G179), .A3(new_n631), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n633), .A2(new_n643), .A3(KEYINPUT21), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n633), .A2(G200), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n633), .A2(new_n393), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n589), .A2(new_n594), .A3(KEYINPUT84), .A4(new_n623), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n626), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n467), .A2(new_n535), .A3(new_n656), .ZN(G372));
  INV_X1    g0457(.A(new_n416), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT18), .B1(new_n421), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n431), .A2(new_n432), .A3(new_n416), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n337), .B1(new_n354), .B2(new_n393), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n360), .B1(new_n357), .B2(new_n361), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n354), .A2(KEYINPUT74), .A3(G200), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n356), .B1(new_n666), .B2(new_n461), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n412), .A2(new_n434), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n319), .B1(new_n669), .B2(KEYINPUT90), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n671), .B(new_n662), .C1(new_n667), .C2(new_n668), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n324), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n615), .A2(new_n622), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n594), .B2(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n575), .A2(new_n577), .A3(G179), .ZN(new_n678));
  AOI21_X1  g0478(.A(G169), .B1(new_n582), .B2(new_n587), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n563), .A2(new_n547), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n623), .A4(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n508), .A2(new_n516), .B1(new_n488), .B2(new_n489), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n648), .A2(new_n649), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT89), .B1(new_n685), .B2(new_n644), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n645), .A2(new_n687), .A3(new_n648), .A4(new_n649), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n532), .A2(new_n594), .A3(new_n589), .A4(new_n623), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n683), .B(new_n622), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n674), .B1(new_n467), .B2(new_n692), .ZN(G369));
  OR2_X1    g0493(.A1(new_n533), .A2(new_n534), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(G213), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n531), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n520), .B2(new_n701), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n647), .A2(new_n700), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n686), .A2(new_n688), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n654), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n685), .A2(new_n644), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n700), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n694), .A2(new_n703), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n684), .A2(new_n701), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0519(.A(new_n212), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G1), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n228), .B2(new_n722), .ZN(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n726));
  XNOR2_X1  g0526(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n691), .A2(new_n728), .A3(new_n701), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n683), .A2(KEYINPUT95), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n682), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n622), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n532), .A2(new_n594), .A3(new_n589), .A4(new_n623), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n520), .A2(new_n713), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n700), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  XOR2_X1   g0540(.A(KEYINPUT94), .B(KEYINPUT30), .Z(new_n741));
  INV_X1    g0541(.A(new_n602), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n522), .A2(new_n582), .A3(new_n587), .A4(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n475), .A2(new_n631), .A3(new_n632), .A4(G179), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n575), .A2(new_n577), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n742), .A2(new_n480), .A3(new_n486), .ZN(new_n747));
  INV_X1    g0547(.A(new_n744), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n582), .A2(new_n587), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n742), .A2(G179), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n750), .A2(new_n487), .A3(new_n633), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n745), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n753), .B2(new_n700), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n650), .A2(new_n653), .A3(new_n700), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n626), .A2(new_n655), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n756), .B1(new_n535), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n740), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n727), .B1(new_n762), .B2(G1), .ZN(G364));
  AND2_X1   g0563(.A1(new_n209), .A2(G13), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n208), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n721), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n710), .B2(G330), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n710), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT96), .Z(new_n770));
  NOR3_X1   g0570(.A1(new_n393), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n209), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G97), .ZN(new_n774));
  NAND2_X1  g0574(.A1(G20), .A2(G179), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n361), .A3(G190), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n774), .B1(new_n216), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT98), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n209), .A2(G179), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT32), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n780), .A2(new_n393), .A3(G200), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n272), .C1(new_n494), .C2(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n393), .A2(new_n361), .ZN(new_n789));
  INV_X1    g0589(.A(new_n775), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n788), .A2(new_n274), .B1(new_n791), .B2(new_n202), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n775), .A2(new_n393), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n789), .A2(new_n780), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n794), .A2(new_n247), .B1(new_n795), .B2(new_n218), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n782), .A2(KEYINPUT32), .A3(new_n783), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n786), .A2(new_n792), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n777), .A2(new_n799), .B1(new_n785), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n794), .A2(new_n802), .B1(new_n795), .B2(new_n629), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n791), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n272), .B1(new_n805), .B2(G326), .ZN(new_n806));
  INV_X1    g0606(.A(new_n782), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G329), .B1(G311), .B2(new_n787), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(G294), .B2(new_n773), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n779), .A2(new_n798), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n254), .B1(G20), .B2(new_n322), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n767), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G13), .A2(G33), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n710), .A2(G20), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n812), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n720), .A2(new_n390), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n820), .A2(G355), .B1(new_n496), .B2(new_n720), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n250), .A2(G45), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT97), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n720), .A2(new_n272), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n228), .B2(G45), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n814), .B(new_n817), .C1(new_n819), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n770), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n691), .A2(new_n701), .ZN(new_n830));
  AND3_X1   g0630(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n460), .A2(new_n701), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n461), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n445), .A2(new_n460), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n701), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n831), .A2(new_n834), .A3(new_n700), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n691), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n840), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n759), .A2(G330), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n830), .A2(KEYINPUT100), .A3(new_n836), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n839), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n767), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n848), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n839), .A2(new_n845), .A3(new_n847), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n760), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n812), .A2(new_n815), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n849), .B1(new_n274), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n805), .A2(G137), .B1(G150), .B2(new_n776), .ZN(new_n859));
  XOR2_X1   g0659(.A(KEYINPUT99), .B(G143), .Z(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n783), .B2(new_n788), .C1(new_n794), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  INV_X1    g0664(.A(G132), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n272), .B1(new_n782), .B2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n216), .A2(new_n785), .B1(new_n795), .B2(new_n202), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n866), .B(new_n867), .C1(G58), .C2(new_n773), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n777), .A2(new_n800), .B1(new_n785), .B2(new_n218), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n272), .B(new_n870), .C1(G294), .C2(new_n793), .ZN(new_n871));
  INV_X1    g0671(.A(new_n795), .ZN(new_n872));
  AOI22_X1  g0672(.A1(G303), .A2(new_n805), .B1(new_n872), .B2(G107), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n807), .A2(G311), .B1(G116), .B2(new_n787), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n774), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n836), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n858), .B1(new_n813), .B2(new_n876), .C1(new_n877), .C2(new_n816), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n856), .A2(new_n878), .ZN(G384));
  NAND2_X1  g0679(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n229), .A2(new_n496), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n541), .B2(KEYINPUT35), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT103), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n227), .B(G77), .C1(new_n247), .C2(new_n216), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n202), .A2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n208), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n589), .A2(new_n594), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n736), .A2(new_n892), .A3(new_n532), .A4(new_n623), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n731), .B1(new_n677), .B2(new_n682), .ZN(new_n894));
  INV_X1    g0694(.A(new_n732), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n622), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n728), .B1(new_n896), .B2(new_n701), .ZN(new_n897));
  INV_X1    g0697(.A(new_n729), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n466), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT106), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT106), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n466), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n673), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT107), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n662), .A2(new_n698), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n840), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT101), .B1(new_n691), .B2(new_n840), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n835), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT14), .B1(new_n357), .B2(new_n322), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n352), .A3(new_n348), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n338), .B(new_n700), .C1(new_n666), .C2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n356), .B(new_n363), .C1(new_n337), .C2(new_n701), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n380), .A2(KEYINPUT16), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n430), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n408), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n698), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n435), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n417), .A2(new_n419), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n431), .ZN(new_n921));
  INV_X1    g0721(.A(new_n698), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n431), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n410), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n916), .A2(new_n408), .B1(new_n416), .B2(new_n922), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n410), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n919), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n435), .A2(new_n918), .B1(new_n925), .B2(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n905), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n910), .A2(new_n338), .A3(new_n701), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n919), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n939), .A2(new_n930), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT105), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n431), .A2(new_n416), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n923), .A3(new_n410), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT37), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n412), .A2(new_n659), .A3(new_n660), .A4(new_n434), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n698), .B1(new_n382), .B2(new_n409), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n945), .A2(new_n925), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n942), .B1(new_n948), .B2(KEYINPUT38), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT38), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n923), .B1(new_n668), .B2(new_n661), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n382), .A2(new_n403), .A3(new_n409), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n947), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT37), .B1(new_n920), .B2(new_n431), .ZN(new_n954));
  AOI22_X1  g0754(.A1(KEYINPUT37), .A2(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(KEYINPUT105), .B(new_n950), .C1(new_n951), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n949), .A2(new_n956), .A3(new_n933), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n941), .B1(new_n940), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n936), .B1(new_n938), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n904), .B(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(G330), .ZN(new_n962));
  INV_X1    g0762(.A(new_n957), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n759), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n756), .B(KEYINPUT108), .C1(new_n535), .C2(new_n758), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n836), .B1(new_n912), .B2(new_n911), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT40), .B1(new_n963), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT40), .B1(new_n931), .B2(new_n933), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n965), .A2(new_n466), .A3(new_n966), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n962), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n974), .B2(new_n973), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n961), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n208), .B2(new_n764), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n961), .A2(new_n976), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n891), .B1(new_n978), .B2(new_n979), .ZN(G367));
  NAND2_X1  g0780(.A1(new_n681), .A2(new_n700), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n892), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n594), .B1(new_n982), .B2(new_n520), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT109), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n701), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n984), .B2(new_n983), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n694), .A2(new_n703), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT110), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n680), .A2(new_n681), .A3(new_n700), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n714), .A4(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT110), .B1(new_n715), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n986), .B1(new_n994), .B2(KEYINPUT42), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT42), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n611), .A2(new_n613), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n700), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n623), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n622), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n998), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n712), .A2(new_n990), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n995), .A2(new_n1005), .A3(new_n1004), .A4(new_n997), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1010), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n721), .B(new_n1015), .Z(new_n1016));
  NAND3_X1  g0816(.A1(new_n715), .A2(new_n716), .A3(new_n990), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT112), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n715), .A2(new_n1019), .A3(new_n716), .A4(new_n990), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT45), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n717), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n990), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n717), .A2(KEYINPUT44), .A3(new_n992), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1018), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1023), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n712), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n714), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n704), .B(new_n1032), .C1(new_n520), .C2(new_n701), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1033), .A2(new_n711), .A3(new_n715), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n711), .B1(new_n1033), .B2(new_n715), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1036), .A2(new_n761), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n712), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1023), .A2(new_n1028), .A3(new_n1038), .A4(new_n1029), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1031), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1016), .B1(new_n1040), .B2(new_n762), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1014), .B1(new_n1041), .B2(new_n766), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1004), .A2(new_n818), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n824), .A2(new_n240), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n818), .B(new_n812), .C1(new_n720), .C2(new_n455), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n849), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n785), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(G77), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n247), .B2(new_n795), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n390), .B(new_n1049), .C1(G159), .C2(new_n776), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G50), .A2(new_n787), .B1(new_n793), .B2(G150), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n860), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1052), .A2(new_n805), .B1(new_n807), .B2(G137), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n772), .A2(new_n216), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT114), .B1(new_n795), .B2(new_n496), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT46), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(KEYINPUT113), .B(G311), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n556), .A2(new_n785), .B1(new_n791), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n272), .B(new_n1060), .C1(G294), .C2(new_n776), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n794), .A2(new_n629), .B1(new_n788), .B2(new_n800), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G317), .B2(new_n807), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1061), .B(new_n1063), .C1(new_n494), .C2(new_n772), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT47), .Z(new_n1066));
  OAI211_X1 g0866(.A(new_n1043), .B(new_n1046), .C1(new_n1066), .C2(new_n813), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1042), .A2(new_n1067), .ZN(G387));
  OAI22_X1  g0868(.A1(new_n795), .A2(new_n274), .B1(new_n782), .B2(new_n296), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n390), .B(new_n1069), .C1(G97), .C2(new_n1047), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n773), .A2(new_n455), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n791), .A2(new_n783), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT116), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n794), .A2(new_n202), .B1(new_n788), .B2(new_n216), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n404), .B2(new_n776), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G303), .A2(new_n787), .B1(new_n793), .B2(G317), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n802), .B2(new_n791), .C1(new_n777), .C2(new_n1059), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(G294), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n772), .A2(new_n800), .B1(new_n795), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(KEYINPUT49), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n272), .B1(new_n807), .B2(G326), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n496), .C2(new_n785), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT49), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n812), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n824), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n237), .B2(G45), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n450), .A2(G50), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT50), .Z(new_n1093));
  OAI211_X1 g0893(.A(new_n723), .B(new_n595), .C1(new_n216), .C2(new_n274), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n820), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1095), .B1(G107), .B2(new_n212), .C1(new_n723), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n849), .B1(new_n1097), .B2(new_n819), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1089), .B1(new_n1098), .B2(KEYINPUT115), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(KEYINPUT115), .B2(new_n1098), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT117), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n706), .B2(new_n818), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1036), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n766), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1037), .A2(new_n722), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n762), .B2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(G393));
  AND2_X1   g0907(.A1(new_n1040), .A2(new_n721), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1031), .A2(new_n1039), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1037), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n992), .A2(new_n818), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n819), .B1(new_n556), .B2(new_n212), .C1(new_n1090), .C2(new_n244), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n767), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n772), .A2(new_n274), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n390), .B(new_n1114), .C1(G87), .C2(new_n1047), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n777), .A2(new_n202), .B1(new_n795), .B2(new_n216), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n807), .B2(new_n1052), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(new_n450), .C2(new_n788), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n805), .A2(G150), .B1(G159), .B2(new_n793), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n390), .B1(new_n785), .B2(new_n494), .C1(new_n772), .C2(new_n496), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n788), .A2(new_n1081), .B1(new_n795), .B2(new_n800), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n777), .A2(new_n629), .B1(new_n782), .B2(new_n802), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n805), .A2(G317), .B1(G311), .B2(new_n793), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1118), .A2(new_n1120), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1113), .B1(new_n1127), .B2(new_n812), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1109), .A2(new_n766), .B1(new_n1111), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1110), .A2(new_n1129), .ZN(G390));
  NAND4_X1  g0930(.A1(new_n965), .A2(new_n466), .A3(G330), .A4(new_n966), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n902), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n901), .B1(new_n739), .B2(new_n466), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n674), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n913), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n760), .B2(new_n836), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n965), .A2(G330), .A3(new_n967), .A4(new_n966), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n908), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n965), .A2(G330), .A3(new_n877), .A4(new_n966), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1136), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n759), .A2(new_n913), .A3(new_n877), .A4(G330), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n896), .A2(new_n701), .A3(new_n833), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1143), .A2(new_n835), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n835), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n738), .B2(new_n833), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n937), .B(new_n957), .C1(new_n1150), .C2(new_n1136), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n938), .B1(new_n908), .B2(new_n913), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1143), .C1(new_n958), .C2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n957), .A2(new_n940), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n941), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1149), .B1(new_n843), .B2(new_n844), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n937), .B1(new_n1157), .B2(new_n1136), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1144), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n913), .B1(new_n1159), .B2(new_n1149), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n945), .A2(new_n925), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n946), .A2(new_n947), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT38), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(KEYINPUT105), .B1(KEYINPUT38), .B2(new_n932), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n938), .B1(new_n1164), .B2(new_n949), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1156), .A2(new_n1158), .B1(new_n1160), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1153), .B1(new_n1166), .B2(new_n1138), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1148), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1151), .B1(new_n958), .B2(new_n1152), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n965), .A2(G330), .A3(new_n966), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n967), .A3(new_n1170), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1171), .A2(new_n1135), .A3(new_n1153), .A4(new_n1147), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1168), .A2(new_n721), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1171), .A2(new_n766), .A3(new_n1153), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n857), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n767), .B1(new_n404), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n872), .A2(G150), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT53), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G159), .B2(new_n773), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT54), .B(G143), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n787), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n807), .A2(G125), .B1(new_n776), .B2(G137), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n794), .A2(new_n865), .B1(new_n791), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n390), .B(new_n1185), .C1(G50), .C2(new_n1047), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n390), .B1(new_n795), .B2(new_n218), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT118), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n777), .A2(new_n494), .B1(new_n785), .B2(new_n216), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1190), .A2(new_n1114), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G97), .A2(new_n787), .B1(new_n793), .B2(G116), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n805), .A2(G283), .B1(new_n807), .B2(G294), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1187), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1176), .B1(new_n1195), .B2(new_n812), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n958), .B2(new_n816), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1174), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1173), .A2(new_n1198), .ZN(G378));
  NAND4_X1  g0999(.A1(new_n957), .A2(new_n965), .A3(new_n966), .A4(new_n967), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1200), .A2(KEYINPUT40), .B1(new_n970), .B2(new_n971), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n698), .B1(new_n304), .B2(new_n305), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n325), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n325), .A2(new_n1202), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1201), .A2(new_n962), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1208), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n973), .B2(G330), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n960), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1208), .B1(new_n1201), .B2(new_n962), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n973), .A2(G330), .A3(new_n1210), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n959), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1208), .A2(new_n815), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n767), .B1(G50), .B2(new_n1175), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1184), .A2(new_n794), .B1(new_n777), .B2(new_n865), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n805), .A2(G125), .B1(G137), .B2(new_n787), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n795), .B2(new_n1180), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G150), .C2(new_n773), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT59), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n267), .B(new_n471), .C1(new_n785), .C2(new_n783), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G124), .B2(new_n807), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n785), .A2(new_n247), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT119), .Z(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n390), .A2(new_n471), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n805), .B2(G116), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n274), .B2(new_n795), .C1(new_n494), .C2(new_n794), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n807), .A2(G283), .B1(new_n455), .B2(new_n787), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n556), .B2(new_n777), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1231), .A2(new_n1234), .A3(new_n1054), .A4(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1232), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1228), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1218), .B1(new_n1241), .B2(new_n812), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1216), .A2(new_n766), .B1(new_n1217), .B2(new_n1242), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1212), .A2(new_n1215), .B1(new_n1172), .B2(new_n1135), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n721), .B1(new_n1244), .B2(KEYINPUT57), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n908), .A2(new_n1139), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1135), .B1(new_n1167), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT57), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1213), .A2(new_n1214), .A3(new_n959), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n959), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT120), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT120), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1212), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1248), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1243), .B1(new_n1245), .B2(new_n1254), .ZN(G375));
  INV_X1    g1055(.A(new_n1016), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1246), .A2(new_n1134), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1148), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1147), .A2(new_n766), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n767), .B1(G68), .B2(new_n1175), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n805), .A2(G132), .B1(new_n807), .B2(G128), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1230), .B(new_n1261), .C1(new_n783), .C2(new_n795), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n390), .B1(new_n1181), .B2(new_n776), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G137), .A2(new_n793), .B1(new_n787), .B2(G150), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1263), .B(new_n1264), .C1(new_n202), .C2(new_n772), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G107), .A2(new_n787), .B1(new_n776), .B2(G116), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1266), .B1(new_n556), .B2(new_n795), .C1(new_n800), .C2(new_n794), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n805), .A2(G294), .B1(new_n807), .B2(G303), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(new_n390), .A3(new_n1071), .A4(new_n1048), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1262), .A2(new_n1265), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1260), .B1(new_n1270), .B2(new_n812), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n913), .B2(new_n816), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1259), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1258), .A2(new_n1274), .ZN(G381));
  NAND3_X1  g1075(.A1(new_n1104), .A2(new_n1106), .A3(new_n828), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n856), .A2(new_n878), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT121), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G378), .A2(KEYINPUT122), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT122), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1173), .A2(new_n1198), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G375), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G387), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G390), .A2(G381), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1280), .A2(new_n1285), .A3(new_n1286), .A4(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(KEYINPUT123), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT124), .B1(new_n856), .B2(new_n878), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n856), .A2(KEYINPUT124), .A3(new_n878), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1246), .A2(new_n1134), .A3(KEYINPUT60), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n721), .B1(new_n1246), .B2(new_n1134), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT60), .B1(new_n1246), .B2(new_n1134), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1297), .B(new_n1299), .C1(new_n1303), .C2(new_n1273), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n722), .B1(new_n1135), .B2(new_n1147), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1257), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1246), .A2(new_n1134), .A3(KEYINPUT60), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1309), .A2(new_n1274), .A3(KEYINPUT124), .A4(new_n1278), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(G2897), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1304), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1304), .B2(new_n1310), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1295), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1296), .B(new_n1298), .C1(new_n1309), .C2(new_n1274), .ZN(new_n1316));
  AND4_X1   g1116(.A1(KEYINPUT124), .A2(new_n1309), .A3(new_n1274), .A4(new_n1278), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1311), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1304), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT125), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G378), .B(new_n1243), .C1(new_n1245), .C2(new_n1254), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n765), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1247), .B(new_n1256), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1217), .A2(new_n1242), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1281), .B(new_n1283), .C1(new_n1323), .C2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1290), .B1(new_n1322), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1294), .B1(new_n1321), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1322), .A2(new_n1327), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1290), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1304), .A2(new_n1310), .ZN(new_n1333));
  AND4_X1   g1133(.A1(new_n1330), .A2(new_n1331), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1330), .B1(new_n1328), .B2(new_n1333), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1329), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(G390), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(new_n1042), .B2(new_n1067), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n828), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1277), .A2(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1339), .A2(new_n1341), .ZN(new_n1342));
  AOI211_X1 g1142(.A(new_n1340), .B(new_n1277), .C1(new_n1042), .C2(new_n1067), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1337), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(G387), .A2(new_n1341), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1345), .B(G390), .C1(new_n1341), .C2(new_n1339), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT63), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n1315), .A3(new_n1320), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1350), .A2(new_n1352), .A3(new_n1347), .A4(new_n1294), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1331), .A2(KEYINPUT63), .A3(new_n1332), .A4(new_n1333), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT127), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1328), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1333), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  OAI22_X1  g1158(.A1(new_n1336), .A2(new_n1347), .B1(new_n1353), .B2(new_n1358), .ZN(G405));
  NAND3_X1  g1159(.A1(G375), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1360));
  AND2_X1   g1160(.A1(new_n1360), .A2(new_n1322), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1333), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1361), .A2(new_n1333), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1347), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  OR2_X1    g1165(.A1(new_n1361), .A2(new_n1333), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1347), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1366), .A2(new_n1367), .A3(new_n1362), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(G402));
endmodule


