

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G2105), .A2(n524), .ZN(n980) );
  XOR2_X1 U551 ( .A(KEYINPUT17), .B(n521), .Z(n981) );
  NOR2_X1 U552 ( .A1(n517), .A2(n802), .ZN(n516) );
  AND2_X1 U553 ( .A1(n899), .A2(n815), .ZN(n517) );
  OR2_X1 U554 ( .A1(n768), .A2(n767), .ZN(n518) );
  XNOR2_X1 U555 ( .A(KEYINPUT107), .B(n763), .ZN(n519) );
  XOR2_X1 U556 ( .A(n719), .B(n718), .Z(n520) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n714) );
  XNOR2_X1 U558 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n736) );
  XNOR2_X1 U559 ( .A(n737), .B(n736), .ZN(n745) );
  INV_X1 U560 ( .A(n886), .ZN(n757) );
  OR2_X1 U561 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U562 ( .A1(n683), .A2(n769), .ZN(n727) );
  NAND2_X1 U563 ( .A1(G8), .A2(n727), .ZN(n768) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n769) );
  XNOR2_X1 U565 ( .A(n525), .B(KEYINPUT66), .ZN(n978) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NAND2_X1 U567 ( .A1(G138), .A2(n981), .ZN(n523) );
  INV_X1 U568 ( .A(G2104), .ZN(n524) );
  NAND2_X1 U569 ( .A1(G102), .A2(n980), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n529) );
  AND2_X1 U571 ( .A1(G2105), .A2(n524), .ZN(n525) );
  NAND2_X1 U572 ( .A1(G126), .A2(n978), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n977) );
  NAND2_X1 U574 ( .A1(G114), .A2(n977), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U576 ( .A1(n529), .A2(n528), .ZN(G164) );
  NAND2_X1 U577 ( .A1(n977), .A2(G113), .ZN(n532) );
  NAND2_X1 U578 ( .A1(G101), .A2(n980), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U580 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U581 ( .A1(G137), .A2(n981), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G125), .A2(n978), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U584 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U585 ( .A(G651), .ZN(n541) );
  NOR2_X1 U586 ( .A1(G543), .A2(n541), .ZN(n537) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n537), .Z(n643) );
  NAND2_X1 U588 ( .A1(G64), .A2(n643), .ZN(n540) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n620) );
  NOR2_X1 U590 ( .A1(G651), .A2(n620), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT65), .B(n538), .Z(n649) );
  NAND2_X1 U592 ( .A1(G52), .A2(n649), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n547) );
  NOR2_X1 U594 ( .A1(n620), .A2(n541), .ZN(n638) );
  NAND2_X1 U595 ( .A1(n638), .A2(G77), .ZN(n544) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT64), .ZN(n641) );
  NAND2_X1 U598 ( .A1(G90), .A2(n641), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n545), .Z(n546) );
  NOR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U603 ( .A1(G99), .A2(n980), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G111), .A2(n977), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n978), .A2(G123), .ZN(n550) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(n550), .Z(n551) );
  NOR2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n981), .A2(G135), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n998) );
  XNOR2_X1 U611 ( .A(G2096), .B(n998), .ZN(n555) );
  OR2_X1 U612 ( .A1(G2100), .A2(n555), .ZN(G156) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  NAND2_X1 U614 ( .A1(n641), .A2(G89), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT73), .B(n556), .Z(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G76), .A2(n638), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n649), .A2(G51), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT74), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G63), .A2(n643), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U627 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n820) );
  NAND2_X1 U631 ( .A1(n820), .A2(G567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U633 ( .A1(G56), .A2(n643), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT14), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT69), .B(n571), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G81), .A2(n641), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT12), .B(n572), .Z(n575) );
  NAND2_X1 U638 ( .A1(n638), .A2(G68), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(n573), .Z(n574) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n649), .A2(G43), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n1007) );
  INV_X1 U645 ( .A(G860), .ZN(n600) );
  OR2_X1 U646 ( .A1(n1007), .A2(n600), .ZN(G153) );
  XNOR2_X1 U647 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U648 ( .A1(n649), .A2(G54), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G92), .A2(n641), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G66), .A2(n643), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G79), .A2(n638), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT15), .ZN(n1004) );
  INV_X1 U656 ( .A(G868), .ZN(n662) );
  NAND2_X1 U657 ( .A1(n1004), .A2(n662), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U660 ( .A(n590), .B(KEYINPUT72), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G65), .A2(n643), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G53), .A2(n649), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n638), .A2(G78), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G91), .A2(n641), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n893) );
  XOR2_X1 U668 ( .A(n893), .B(KEYINPUT68), .Z(G299) );
  XNOR2_X1 U669 ( .A(KEYINPUT75), .B(G868), .ZN(n597) );
  NOR2_X1 U670 ( .A1(G286), .A2(n597), .ZN(n599) );
  NOR2_X1 U671 ( .A1(G299), .A2(G868), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U673 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U674 ( .A(n1004), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n601), .A2(n608), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(n1004), .A2(n662), .ZN(n603) );
  XOR2_X1 U678 ( .A(KEYINPUT76), .B(n603), .Z(n604) );
  NOR2_X1 U679 ( .A1(G559), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G868), .A2(n1007), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U682 ( .A(KEYINPUT77), .B(n607), .Z(G282) );
  NAND2_X1 U683 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(n1007), .ZN(n659) );
  NOR2_X1 U685 ( .A1(n659), .A2(G860), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G67), .A2(n643), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G55), .A2(n649), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n638), .A2(G80), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G93), .A2(n641), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  OR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n663) );
  XOR2_X1 U693 ( .A(n616), .B(n663), .Z(G145) );
  NAND2_X1 U694 ( .A1(G49), .A2(n649), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT78), .B(n619), .Z(n624) );
  NAND2_X1 U698 ( .A1(G87), .A2(n620), .ZN(n621) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(n621), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n643), .A2(n622), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U702 ( .A1(G72), .A2(n638), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G47), .A2(n649), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G85), .A2(n641), .ZN(n627) );
  XNOR2_X1 U706 ( .A(KEYINPUT67), .B(n627), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n643), .A2(G60), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U710 ( .A1(n638), .A2(G75), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G88), .A2(n641), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U713 ( .A1(G62), .A2(n643), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G50), .A2(n649), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(G166) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n640) );
  NAND2_X1 U718 ( .A1(G73), .A2(n638), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n640), .B(n639), .ZN(n648) );
  NAND2_X1 U720 ( .A1(G86), .A2(n641), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G61), .A2(n643), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n646), .Z(n647) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n649), .A2(G48), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(G305) );
  XOR2_X1 U728 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n653) );
  XNOR2_X1 U729 ( .A(G299), .B(KEYINPUT83), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n654) );
  XOR2_X1 U731 ( .A(n663), .B(n654), .Z(n656) );
  XNOR2_X1 U732 ( .A(G290), .B(G166), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U734 ( .A(n657), .B(G305), .Z(n658) );
  XNOR2_X1 U735 ( .A(G288), .B(n658), .ZN(n1005) );
  XNOR2_X1 U736 ( .A(n1005), .B(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n660), .A2(G868), .ZN(n661) );
  XOR2_X1 U738 ( .A(KEYINPUT85), .B(n661), .Z(n665) );
  NAND2_X1 U739 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G108), .A2(n671), .ZN(n945) );
  NAND2_X1 U750 ( .A1(G567), .A2(n945), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G132), .A2(G82), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(KEYINPUT86), .ZN(n673) );
  XNOR2_X1 U753 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  NOR2_X1 U754 ( .A1(G218), .A2(n674), .ZN(n675) );
  XOR2_X1 U755 ( .A(KEYINPUT87), .B(n675), .Z(n676) );
  NAND2_X1 U756 ( .A1(G96), .A2(n676), .ZN(n944) );
  NAND2_X1 U757 ( .A1(G2106), .A2(n944), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U759 ( .A(KEYINPUT88), .B(n679), .Z(G319) );
  INV_X1 U760 ( .A(G319), .ZN(n681) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n822) );
  NAND2_X1 U763 ( .A1(n822), .A2(G36), .ZN(G176) );
  XNOR2_X1 U764 ( .A(G166), .B(KEYINPUT89), .ZN(G303) );
  NOR2_X1 U765 ( .A1(G2090), .A2(G303), .ZN(n682) );
  NAND2_X1 U766 ( .A1(G8), .A2(n682), .ZN(n746) );
  XOR2_X1 U767 ( .A(G2078), .B(KEYINPUT25), .Z(n867) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n770) );
  INV_X1 U769 ( .A(n770), .ZN(n683) );
  NOR2_X1 U770 ( .A1(n867), .A2(n727), .ZN(n685) );
  INV_X1 U771 ( .A(n727), .ZN(n700) );
  NOR2_X1 U772 ( .A1(n700), .A2(G1961), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U774 ( .A(KEYINPUT97), .B(n686), .ZN(n720) );
  NAND2_X1 U775 ( .A1(G171), .A2(n720), .ZN(n687) );
  XNOR2_X1 U776 ( .A(n687), .B(KEYINPUT98), .ZN(n712) );
  INV_X1 U777 ( .A(G1996), .ZN(n688) );
  NOR2_X1 U778 ( .A1(n727), .A2(n688), .ZN(n689) );
  XOR2_X1 U779 ( .A(n689), .B(KEYINPUT26), .Z(n691) );
  NAND2_X1 U780 ( .A1(n727), .A2(G1341), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U782 ( .A1(n1007), .A2(n692), .ZN(n696) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n727), .ZN(n694) );
  NAND2_X1 U784 ( .A1(G2067), .A2(n700), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U786 ( .A1(n1004), .A2(n697), .ZN(n695) );
  OR2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n1004), .A2(n697), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n700), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U791 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  AND2_X1 U792 ( .A1(G1956), .A2(n727), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n893), .A2(n706), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n893), .A2(n706), .ZN(n707) );
  XOR2_X1 U797 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U799 ( .A(KEYINPUT29), .B(n710), .Z(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n725) );
  XNOR2_X1 U801 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(KEYINPUT30), .ZN(n719) );
  NOR2_X1 U803 ( .A1(n768), .A2(G1966), .ZN(n715) );
  XNOR2_X1 U804 ( .A(n715), .B(n714), .ZN(n739) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n727), .ZN(n741) );
  INV_X1 U806 ( .A(G8), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n741), .A2(n716), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n739), .A2(n717), .ZN(n718) );
  NOR2_X1 U809 ( .A1(G168), .A2(n520), .ZN(n722) );
  NOR2_X1 U810 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U812 ( .A(KEYINPUT31), .B(n723), .Z(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n738) );
  AND2_X1 U814 ( .A1(G286), .A2(G8), .ZN(n726) );
  NAND2_X1 U815 ( .A1(n738), .A2(n726), .ZN(n735) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n727), .ZN(n728) );
  XOR2_X1 U817 ( .A(KEYINPUT103), .B(n728), .Z(n731) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n768), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(KEYINPUT102), .ZN(n730) );
  NOR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G303), .ZN(n733) );
  OR2_X1 U822 ( .A1(n716), .A2(n733), .ZN(n734) );
  AND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U825 ( .A(n740), .B(KEYINPUT101), .ZN(n743) );
  NAND2_X1 U826 ( .A1(n741), .A2(G8), .ZN(n742) );
  NAND2_X1 U827 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U828 ( .A1(n745), .A2(n744), .ZN(n750) );
  NAND2_X1 U829 ( .A1(n746), .A2(n750), .ZN(n747) );
  NAND2_X1 U830 ( .A1(n747), .A2(n768), .ZN(n762) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n889) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n895) );
  XOR2_X1 U833 ( .A(n895), .B(KEYINPUT105), .Z(n748) );
  NOR2_X1 U834 ( .A1(n889), .A2(n748), .ZN(n749) );
  XNOR2_X1 U835 ( .A(n749), .B(KEYINPUT106), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n891) );
  INV_X1 U838 ( .A(n891), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n768), .A2(n752), .ZN(n753) );
  AND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U841 ( .A1(KEYINPUT33), .A2(n755), .ZN(n760) );
  NAND2_X1 U842 ( .A1(n889), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n768), .A2(n756), .ZN(n758) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n886) );
  OR2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U847 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n764) );
  XNOR2_X1 U848 ( .A(n764), .B(KEYINPUT94), .ZN(n766) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XNOR2_X1 U850 ( .A(n766), .B(n765), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n519), .A2(n518), .ZN(n803) );
  XNOR2_X1 U852 ( .A(G1986), .B(G290), .ZN(n899) );
  NOR2_X1 U853 ( .A1(n770), .A2(n769), .ZN(n815) );
  NAND2_X1 U854 ( .A1(G104), .A2(n980), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G140), .A2(n981), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n773), .ZN(n778) );
  NAND2_X1 U858 ( .A1(G116), .A2(n977), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G128), .A2(n978), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U861 ( .A(KEYINPUT35), .B(n776), .Z(n777) );
  NOR2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U863 ( .A(KEYINPUT36), .B(n779), .ZN(n974) );
  XNOR2_X1 U864 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NOR2_X1 U865 ( .A1(n974), .A2(n812), .ZN(n835) );
  NAND2_X1 U866 ( .A1(n815), .A2(n835), .ZN(n810) );
  NAND2_X1 U867 ( .A1(G117), .A2(n977), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G129), .A2(n978), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U870 ( .A(KEYINPUT92), .B(n782), .ZN(n786) );
  NAND2_X1 U871 ( .A1(G105), .A2(n980), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT38), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(KEYINPUT93), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n981), .A2(G141), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n990) );
  AND2_X1 U877 ( .A1(n990), .A2(G1996), .ZN(n799) );
  NAND2_X1 U878 ( .A1(n981), .A2(G131), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G107), .A2(n977), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G119), .A2(n978), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n980), .A2(G95), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT90), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U886 ( .A(KEYINPUT91), .B(n796), .Z(n804) );
  INV_X1 U887 ( .A(n804), .ZN(n994) );
  INV_X1 U888 ( .A(G1991), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n994), .A2(n797), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n842) );
  INV_X1 U891 ( .A(n815), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n842), .A2(n800), .ZN(n807) );
  INV_X1 U893 ( .A(n807), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n810), .A2(n801), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n516), .ZN(n818) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n990), .ZN(n856) );
  NOR2_X1 U897 ( .A1(G1991), .A2(n804), .ZN(n840) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n840), .A2(n805), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n856), .A2(n808), .ZN(n809) );
  XNOR2_X1 U902 ( .A(n809), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n974), .A2(n812), .ZN(n837) );
  NAND2_X1 U905 ( .A1(n813), .A2(n837), .ZN(n814) );
  XNOR2_X1 U906 ( .A(KEYINPUT108), .B(n814), .ZN(n816) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U909 ( .A(n819), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U915 ( .A(KEYINPUT111), .B(n824), .Z(G188) );
  NAND2_X1 U917 ( .A1(G124), .A2(n978), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n825), .B(KEYINPUT44), .ZN(n827) );
  NAND2_X1 U919 ( .A1(G136), .A2(n981), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(KEYINPUT112), .B(n828), .ZN(n833) );
  NAND2_X1 U922 ( .A1(G100), .A2(n980), .ZN(n830) );
  NAND2_X1 U923 ( .A1(G112), .A2(n977), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  XOR2_X1 U925 ( .A(KEYINPUT113), .B(n831), .Z(n832) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U927 ( .A(KEYINPUT114), .B(n834), .ZN(G162) );
  INV_X1 U928 ( .A(n835), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(n844) );
  XNOR2_X1 U930 ( .A(G160), .B(G2084), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n838), .A2(n998), .ZN(n839) );
  NOR2_X1 U932 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U934 ( .A1(n844), .A2(n843), .ZN(n861) );
  NAND2_X1 U935 ( .A1(G103), .A2(n980), .ZN(n846) );
  NAND2_X1 U936 ( .A1(G139), .A2(n981), .ZN(n845) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(n851) );
  NAND2_X1 U938 ( .A1(G115), .A2(n977), .ZN(n848) );
  NAND2_X1 U939 ( .A1(G127), .A2(n978), .ZN(n847) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U941 ( .A(KEYINPUT47), .B(n849), .Z(n850) );
  NOR2_X1 U942 ( .A1(n851), .A2(n850), .ZN(n999) );
  XOR2_X1 U943 ( .A(G2072), .B(n999), .Z(n853) );
  XOR2_X1 U944 ( .A(G164), .B(G2078), .Z(n852) );
  NOR2_X1 U945 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U946 ( .A(KEYINPUT50), .B(n854), .Z(n859) );
  XOR2_X1 U947 ( .A(G2090), .B(G162), .Z(n855) );
  NOR2_X1 U948 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U949 ( .A(KEYINPUT51), .B(n857), .ZN(n858) );
  NOR2_X1 U950 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U951 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U952 ( .A(KEYINPUT52), .B(n862), .ZN(n863) );
  NAND2_X1 U953 ( .A1(n863), .A2(G29), .ZN(n942) );
  XNOR2_X1 U954 ( .A(G1996), .B(G32), .ZN(n865) );
  XNOR2_X1 U955 ( .A(G33), .B(G2072), .ZN(n864) );
  NOR2_X1 U956 ( .A1(n865), .A2(n864), .ZN(n872) );
  XOR2_X1 U957 ( .A(G2067), .B(G26), .Z(n866) );
  NAND2_X1 U958 ( .A1(n866), .A2(G28), .ZN(n870) );
  XNOR2_X1 U959 ( .A(G27), .B(n867), .ZN(n868) );
  XNOR2_X1 U960 ( .A(KEYINPUT120), .B(n868), .ZN(n869) );
  NOR2_X1 U961 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U962 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U963 ( .A(G25), .B(G1991), .ZN(n873) );
  NOR2_X1 U964 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U965 ( .A(n875), .B(KEYINPUT121), .ZN(n876) );
  XNOR2_X1 U966 ( .A(n876), .B(KEYINPUT53), .ZN(n879) );
  XOR2_X1 U967 ( .A(G2084), .B(G34), .Z(n877) );
  XNOR2_X1 U968 ( .A(KEYINPUT54), .B(n877), .ZN(n878) );
  NAND2_X1 U969 ( .A1(n879), .A2(n878), .ZN(n881) );
  XNOR2_X1 U970 ( .A(G35), .B(G2090), .ZN(n880) );
  NOR2_X1 U971 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U972 ( .A(n882), .B(KEYINPUT122), .ZN(n883) );
  NOR2_X1 U973 ( .A1(G29), .A2(n883), .ZN(n884) );
  XNOR2_X1 U974 ( .A(KEYINPUT55), .B(n884), .ZN(n885) );
  NAND2_X1 U975 ( .A1(n885), .A2(G11), .ZN(n940) );
  XNOR2_X1 U976 ( .A(G16), .B(KEYINPUT56), .ZN(n913) );
  XNOR2_X1 U977 ( .A(G168), .B(G1966), .ZN(n887) );
  NAND2_X1 U978 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U979 ( .A(KEYINPUT57), .B(n888), .ZN(n911) );
  NAND2_X1 U980 ( .A1(G303), .A2(G1971), .ZN(n901) );
  INV_X1 U981 ( .A(n889), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U983 ( .A(n892), .B(KEYINPUT123), .ZN(n897) );
  XOR2_X1 U984 ( .A(n893), .B(G1956), .Z(n894) );
  NOR2_X1 U985 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U986 ( .A1(n897), .A2(n896), .ZN(n898) );
  NOR2_X1 U987 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U988 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U989 ( .A(n902), .B(KEYINPUT124), .ZN(n904) );
  XOR2_X1 U990 ( .A(G1961), .B(G171), .Z(n903) );
  NOR2_X1 U991 ( .A1(n904), .A2(n903), .ZN(n908) );
  XNOR2_X1 U992 ( .A(n1007), .B(G1341), .ZN(n906) );
  XNOR2_X1 U993 ( .A(n1004), .B(G1348), .ZN(n905) );
  NOR2_X1 U994 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U995 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U996 ( .A(KEYINPUT125), .B(n909), .ZN(n910) );
  NAND2_X1 U997 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U998 ( .A1(n913), .A2(n912), .ZN(n938) );
  INV_X1 U999 ( .A(G16), .ZN(n936) );
  XOR2_X1 U1000 ( .A(G20), .B(G1956), .Z(n917) );
  XNOR2_X1 U1001 ( .A(G1981), .B(G6), .ZN(n915) );
  XNOR2_X1 U1002 ( .A(G19), .B(G1341), .ZN(n914) );
  NOR2_X1 U1003 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1004 ( .A1(n917), .A2(n916), .ZN(n920) );
  XOR2_X1 U1005 ( .A(KEYINPUT59), .B(G1348), .Z(n918) );
  XNOR2_X1 U1006 ( .A(G4), .B(n918), .ZN(n919) );
  NOR2_X1 U1007 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1008 ( .A(KEYINPUT60), .B(n921), .ZN(n931) );
  XNOR2_X1 U1009 ( .A(G1966), .B(KEYINPUT126), .ZN(n922) );
  XNOR2_X1 U1010 ( .A(n922), .B(G21), .ZN(n929) );
  XNOR2_X1 U1011 ( .A(G1971), .B(G22), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(G23), .B(G1976), .ZN(n923) );
  NOR2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G1986), .B(G24), .Z(n925) );
  NAND2_X1 U1015 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1016 ( .A(KEYINPUT58), .B(n927), .ZN(n928) );
  NOR2_X1 U1017 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1018 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1019 ( .A(G5), .B(G1961), .ZN(n932) );
  NOR2_X1 U1020 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1021 ( .A(KEYINPUT61), .B(n934), .ZN(n935) );
  NAND2_X1 U1022 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1023 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1024 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1025 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1026 ( .A(KEYINPUT62), .B(n943), .Z(G311) );
  XNOR2_X1 U1027 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1028 ( .A(G132), .ZN(G219) );
  INV_X1 U1029 ( .A(G120), .ZN(G236) );
  INV_X1 U1030 ( .A(G96), .ZN(G221) );
  INV_X1 U1031 ( .A(G82), .ZN(G220) );
  INV_X1 U1032 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1033 ( .A1(n945), .A2(n944), .ZN(G325) );
  INV_X1 U1034 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1035 ( .A(G2443), .B(G2430), .Z(n947) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G2451), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(n947), .B(n946), .ZN(n954) );
  XOR2_X1 U1038 ( .A(G2438), .B(KEYINPUT109), .Z(n949) );
  XNOR2_X1 U1039 ( .A(G1348), .B(G2454), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(n949), .B(n948), .ZN(n950) );
  XOR2_X1 U1041 ( .A(n950), .B(G2435), .Z(n952) );
  XNOR2_X1 U1042 ( .A(G2446), .B(G2427), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n952), .B(n951), .ZN(n953) );
  XNOR2_X1 U1044 ( .A(n954), .B(n953), .ZN(n955) );
  NAND2_X1 U1045 ( .A1(n955), .A2(G14), .ZN(n956) );
  XOR2_X1 U1046 ( .A(KEYINPUT110), .B(n956), .Z(G401) );
  XOR2_X1 U1047 ( .A(G2100), .B(G2096), .Z(n958) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G2072), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(n958), .B(n957), .ZN(n962) );
  XOR2_X1 U1050 ( .A(G2678), .B(KEYINPUT42), .Z(n960) );
  XNOR2_X1 U1051 ( .A(G2067), .B(KEYINPUT43), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n960), .B(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(n962), .B(n961), .Z(n964) );
  XNOR2_X1 U1054 ( .A(G2078), .B(G2084), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(G227) );
  XOR2_X1 U1056 ( .A(G1966), .B(G1971), .Z(n966) );
  XNOR2_X1 U1057 ( .A(G1996), .B(G1986), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n966), .B(n965), .ZN(n967) );
  XOR2_X1 U1059 ( .A(n967), .B(G2474), .Z(n969) );
  XNOR2_X1 U1060 ( .A(G1991), .B(G1956), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n973) );
  XOR2_X1 U1062 ( .A(KEYINPUT41), .B(G1976), .Z(n971) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G1961), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n971), .B(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n973), .B(n972), .ZN(G229) );
  XNOR2_X1 U1066 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n974), .B(KEYINPUT46), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n993) );
  NAND2_X1 U1069 ( .A1(G118), .A2(n977), .ZN(n989) );
  NAND2_X1 U1070 ( .A1(G130), .A2(n978), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(KEYINPUT115), .B(n979), .ZN(n987) );
  NAND2_X1 U1072 ( .A1(G106), .A2(n980), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(G142), .A2(n981), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT45), .B(n984), .Z(n985) );
  XNOR2_X1 U1076 ( .A(KEYINPUT116), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n991) );
  XOR2_X1 U1079 ( .A(n991), .B(n990), .Z(n992) );
  XOR2_X1 U1080 ( .A(n993), .B(n992), .Z(n996) );
  XNOR2_X1 U1081 ( .A(G164), .B(n994), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n996), .B(n995), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1084 ( .A(G160), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(n1002), .B(G162), .ZN(n1003) );
  NOR2_X1 U1087 ( .A1(G37), .A2(n1003), .ZN(G395) );
  XNOR2_X1 U1088 ( .A(G171), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(n1006), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1090 ( .A(n1007), .B(G286), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1010), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(KEYINPUT118), .B(n1011), .ZN(G397) );
  NOR2_X1 U1094 ( .A1(G227), .A2(G229), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT119), .B(n1012), .Z(n1013) );
  XNOR2_X1 U1096 ( .A(n1013), .B(KEYINPUT49), .ZN(n1014) );
  NOR2_X1 U1097 ( .A1(G401), .A2(n1014), .ZN(n1015) );
  AND2_X1 U1098 ( .A1(n1015), .A2(G319), .ZN(n1017) );
  NOR2_X1 U1099 ( .A1(G395), .A2(G397), .ZN(n1016) );
  NAND2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(G225) );
  INV_X1 U1101 ( .A(G225), .ZN(G308) );
  INV_X1 U1102 ( .A(G108), .ZN(G238) );
endmodule

