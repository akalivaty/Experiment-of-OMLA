

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782;

  INV_X1 U380 ( .A(n710), .ZN(n362) );
  INV_X1 U381 ( .A(n619), .ZN(n367) );
  XNOR2_X1 U382 ( .A(n602), .B(KEYINPUT19), .ZN(n610) );
  OR2_X1 U383 ( .A1(n674), .A2(n429), .ZN(n385) );
  XNOR2_X1 U384 ( .A(n394), .B(n393), .ZN(n537) );
  XNOR2_X1 U385 ( .A(n471), .B(KEYINPUT3), .ZN(n394) );
  NAND2_X1 U386 ( .A1(n770), .A2(G224), .ZN(n540) );
  XNOR2_X1 U387 ( .A(n526), .B(KEYINPUT4), .ZN(n546) );
  INV_X1 U388 ( .A(n361), .ZN(n685) );
  NAND2_X1 U389 ( .A1(n363), .A2(n362), .ZN(n361) );
  XNOR2_X1 U390 ( .A(n682), .B(n364), .ZN(n363) );
  INV_X1 U391 ( .A(n681), .ZN(n364) );
  NOR2_X2 U392 ( .A1(n367), .A2(n365), .ZN(n630) );
  NAND2_X1 U393 ( .A1(n366), .A2(n618), .ZN(n365) );
  INV_X1 U394 ( .A(n627), .ZN(n366) );
  NAND2_X1 U395 ( .A1(n655), .A2(KEYINPUT44), .ZN(n653) );
  NAND2_X1 U396 ( .A1(n372), .A2(n410), .ZN(n655) );
  AND2_X2 U397 ( .A1(n580), .A2(n452), .ZN(n567) );
  AND2_X2 U398 ( .A1(n369), .A2(n419), .ZN(n371) );
  NAND2_X1 U399 ( .A1(n426), .A2(n431), .ZN(n602) );
  INV_X4 U400 ( .A(G953), .ZN(n770) );
  XNOR2_X1 U401 ( .A(n567), .B(n566), .ZN(n425) );
  INV_X1 U402 ( .A(n598), .ZN(n368) );
  NAND2_X2 U403 ( .A1(n659), .A2(n712), .ZN(n432) );
  NOR2_X2 U404 ( .A1(n665), .A2(n664), .ZN(n698) );
  XNOR2_X2 U405 ( .A(G113), .B(KEYINPUT87), .ZN(n471) );
  XNOR2_X2 U406 ( .A(n546), .B(n466), .ZN(n767) );
  AND2_X1 U407 ( .A1(n445), .A2(n443), .ZN(n651) );
  NOR2_X1 U408 ( .A1(n581), .A2(n622), .ZN(n582) );
  NAND2_X1 U409 ( .A1(n432), .A2(n660), .ZN(n665) );
  NAND2_X1 U410 ( .A1(n434), .A2(n373), .ZN(n395) );
  OR2_X1 U411 ( .A1(n777), .A2(n436), .ZN(n435) );
  XNOR2_X1 U412 ( .A(n448), .B(n447), .ZN(n627) );
  INV_X2 U413 ( .A(n590), .ZN(n718) );
  NAND2_X1 U414 ( .A1(n610), .A2(n561), .ZN(n563) );
  INV_X1 U415 ( .A(n640), .ZN(n369) );
  NAND2_X1 U416 ( .A1(n570), .A2(n454), .ZN(n639) );
  XNOR2_X2 U417 ( .A(n631), .B(KEYINPUT111), .ZN(n383) );
  XNOR2_X2 U418 ( .A(n767), .B(n488), .ZN(n486) );
  XNOR2_X1 U419 ( .A(n384), .B(n503), .ZN(n721) );
  NAND2_X1 U420 ( .A1(n699), .A2(n532), .ZN(n384) );
  AND2_X1 U421 ( .A1(G234), .A2(n770), .ZN(n495) );
  OR2_X1 U422 ( .A1(n573), .A2(n577), .ZN(n574) );
  INV_X1 U423 ( .A(KEYINPUT36), .ZN(n381) );
  XNOR2_X1 U424 ( .A(G146), .B(G125), .ZN(n490) );
  AND2_X1 U425 ( .A1(n439), .A2(n437), .ZN(n617) );
  INV_X1 U426 ( .A(G143), .ZN(n462) );
  XNOR2_X1 U427 ( .A(n389), .B(KEYINPUT78), .ZN(n436) );
  NAND2_X1 U428 ( .A1(n765), .A2(KEYINPUT2), .ZN(n389) );
  NOR2_X1 U429 ( .A1(n721), .A2(n722), .ZN(n454) );
  OR2_X2 U430 ( .A1(n402), .A2(n400), .ZN(n609) );
  NAND2_X1 U431 ( .A1(n404), .A2(n403), .ZN(n402) );
  NAND2_X1 U432 ( .A1(n450), .A2(G902), .ZN(n403) );
  XNOR2_X1 U433 ( .A(G119), .B(G116), .ZN(n393) );
  XNOR2_X1 U434 ( .A(G134), .B(G116), .ZN(n523) );
  INV_X1 U435 ( .A(KEYINPUT100), .ZN(n522) );
  XNOR2_X1 U436 ( .A(G107), .B(G122), .ZN(n520) );
  XOR2_X1 U437 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n521) );
  XNOR2_X1 U438 ( .A(G107), .B(G104), .ZN(n481) );
  INV_X1 U439 ( .A(n765), .ZN(n433) );
  INV_X1 U440 ( .A(KEYINPUT109), .ZN(n421) );
  NAND2_X1 U441 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U442 ( .A(n718), .ZN(n423) );
  XNOR2_X1 U443 ( .A(n632), .B(KEYINPUT108), .ZN(n424) );
  XNOR2_X1 U444 ( .A(n620), .B(KEYINPUT41), .ZN(n749) );
  XNOR2_X1 U445 ( .A(n624), .B(KEYINPUT39), .ZN(n637) );
  NAND2_X1 U446 ( .A1(n391), .A2(n390), .ZN(n624) );
  NOR2_X1 U447 ( .A1(n733), .A2(n622), .ZN(n390) );
  INV_X1 U448 ( .A(n623), .ZN(n391) );
  OR2_X1 U449 ( .A1(n382), .A2(n381), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n388), .B(n642), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n416), .B(KEYINPUT103), .ZN(n415) );
  NAND2_X1 U452 ( .A1(n718), .A2(n408), .ZN(n416) );
  AND2_X1 U453 ( .A1(n431), .A2(n430), .ZN(n397) );
  NAND2_X1 U454 ( .A1(n454), .A2(n609), .ZN(n622) );
  XNOR2_X1 U455 ( .A(n519), .B(n518), .ZN(n573) );
  BUF_X1 U456 ( .A(n721), .Z(n408) );
  XNOR2_X1 U457 ( .A(n499), .B(n498), .ZN(n699) );
  BUF_X1 U458 ( .A(n698), .Z(n704) );
  NOR2_X1 U459 ( .A1(n770), .A2(G952), .ZN(n710) );
  NOR2_X1 U460 ( .A1(n444), .A2(n649), .ZN(n443) );
  NOR2_X1 U461 ( .A1(n648), .A2(n725), .ZN(n444) );
  NOR2_X1 U462 ( .A1(n616), .A2(n370), .ZN(n439) );
  INV_X1 U463 ( .A(KEYINPUT83), .ZN(n604) );
  XNOR2_X1 U464 ( .A(KEYINPUT46), .B(KEYINPUT64), .ZN(n447) );
  XNOR2_X1 U465 ( .A(n487), .B(n451), .ZN(n450) );
  INV_X1 U466 ( .A(G469), .ZN(n451) );
  OR2_X1 U467 ( .A1(n450), .A2(G902), .ZN(n401) );
  NAND2_X1 U468 ( .A1(n413), .A2(n450), .ZN(n404) );
  XNOR2_X1 U469 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n467) );
  XOR2_X1 U470 ( .A(G101), .B(G137), .Z(n468) );
  XNOR2_X1 U471 ( .A(G143), .B(G113), .ZN(n510) );
  XNOR2_X1 U472 ( .A(G122), .B(KEYINPUT98), .ZN(n514) );
  XOR2_X1 U473 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n515) );
  NAND2_X1 U474 ( .A1(n442), .A2(n441), .ZN(n375) );
  NAND2_X1 U475 ( .A1(n490), .A2(KEYINPUT10), .ZN(n442) );
  INV_X1 U476 ( .A(KEYINPUT10), .ZN(n489) );
  XNOR2_X1 U477 ( .A(n464), .B(KEYINPUT69), .ZN(n465) );
  INV_X1 U478 ( .A(G134), .ZN(n464) );
  INV_X1 U479 ( .A(n548), .ZN(n660) );
  XNOR2_X1 U480 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n541) );
  NAND2_X1 U481 ( .A1(G237), .A2(G234), .ZN(n456) );
  XNOR2_X1 U482 ( .A(n633), .B(n396), .ZN(n733) );
  INV_X1 U483 ( .A(KEYINPUT38), .ZN(n396) );
  NAND2_X1 U484 ( .A1(n552), .A2(n660), .ZN(n430) );
  AND2_X1 U485 ( .A1(n385), .A2(n427), .ZN(n426) );
  NOR2_X1 U486 ( .A1(n428), .A2(n732), .ZN(n427) );
  INV_X1 U487 ( .A(n430), .ZN(n428) );
  XNOR2_X1 U488 ( .A(G128), .B(G119), .ZN(n492) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(G110), .Z(n493) );
  XNOR2_X1 U490 ( .A(n375), .B(n440), .ZN(n766) );
  INV_X1 U491 ( .A(n491), .ZN(n440) );
  INV_X1 U492 ( .A(G146), .ZN(n488) );
  XOR2_X1 U493 ( .A(G137), .B(G140), .Z(n491) );
  NAND2_X1 U494 ( .A1(n412), .A2(n369), .ZN(n411) );
  XNOR2_X1 U495 ( .A(n639), .B(KEYINPUT105), .ZN(n412) );
  NAND2_X1 U496 ( .A1(n392), .A2(n449), .ZN(n623) );
  INV_X1 U497 ( .A(n599), .ZN(n449) );
  XNOR2_X1 U498 ( .A(n479), .B(KEYINPUT30), .ZN(n392) );
  XNOR2_X1 U499 ( .A(n625), .B(n575), .ZN(n598) );
  XNOR2_X1 U500 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n535) );
  XNOR2_X1 U501 ( .A(n525), .B(n524), .ZN(n531) );
  XNOR2_X1 U502 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U503 ( .A(n680), .B(KEYINPUT59), .Z(n681) );
  XNOR2_X1 U504 ( .A(n422), .B(n420), .ZN(n634) );
  XNOR2_X1 U505 ( .A(n421), .B(KEYINPUT43), .ZN(n420) );
  XNOR2_X1 U506 ( .A(n398), .B(KEYINPUT42), .ZN(n781) );
  NAND2_X1 U507 ( .A1(n637), .A2(n758), .ZN(n765) );
  XNOR2_X1 U508 ( .A(n626), .B(KEYINPUT40), .ZN(n782) );
  OR2_X2 U509 ( .A1(n377), .A2(n376), .ZN(n603) );
  NAND2_X1 U510 ( .A1(n379), .A2(n374), .ZN(n377) );
  XNOR2_X1 U511 ( .A(n386), .B(n399), .ZN(n410) );
  INV_X1 U512 ( .A(KEYINPUT35), .ZN(n399) );
  XNOR2_X1 U513 ( .A(n594), .B(n593), .ZN(n646) );
  XNOR2_X1 U514 ( .A(n569), .B(KEYINPUT104), .ZN(n645) );
  AND2_X1 U515 ( .A1(n446), .A2(n725), .ZN(n647) );
  INV_X1 U516 ( .A(n699), .ZN(n406) );
  AND2_X1 U517 ( .A1(n615), .A2(KEYINPUT79), .ZN(n370) );
  AND2_X1 U518 ( .A1(n646), .A2(n645), .ZN(n372) );
  NOR2_X1 U519 ( .A1(n777), .A2(n433), .ZN(n373) );
  AND2_X1 U520 ( .A1(n718), .A2(n378), .ZN(n374) );
  XNOR2_X1 U521 ( .A(n375), .B(n508), .ZN(n516) );
  NOR2_X1 U522 ( .A1(n383), .A2(n381), .ZN(n376) );
  NAND2_X1 U523 ( .A1(n383), .A2(n380), .ZN(n379) );
  AND2_X1 U524 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U525 ( .A(n602), .ZN(n382) );
  NAND2_X1 U526 ( .A1(n721), .A2(n600), .ZN(n601) );
  INV_X1 U527 ( .A(n490), .ZN(n544) );
  NAND2_X1 U528 ( .A1(n397), .A2(n385), .ZN(n633) );
  NAND2_X1 U529 ( .A1(n387), .A2(n644), .ZN(n386) );
  NAND2_X1 U530 ( .A1(n750), .A2(n641), .ZN(n388) );
  NAND2_X1 U531 ( .A1(n395), .A2(n714), .ZN(n715) );
  NOR2_X1 U532 ( .A1(n662), .A2(n395), .ZN(n663) );
  XNOR2_X1 U533 ( .A(n395), .B(KEYINPUT125), .ZN(n769) );
  NAND2_X1 U534 ( .A1(n782), .A2(n781), .ZN(n448) );
  NAND2_X1 U535 ( .A1(n749), .A2(n621), .ZN(n398) );
  INV_X1 U536 ( .A(n410), .ZN(n686) );
  XNOR2_X2 U537 ( .A(n609), .B(KEYINPUT1), .ZN(n570) );
  NOR2_X1 U538 ( .A1(n413), .A2(n401), .ZN(n400) );
  XNOR2_X2 U539 ( .A(n486), .B(n485), .ZN(n413) );
  OR2_X2 U540 ( .A1(n636), .A2(n435), .ZN(n638) );
  XNOR2_X1 U541 ( .A(n701), .B(n405), .ZN(n703) );
  INV_X1 U542 ( .A(n702), .ZN(n405) );
  XNOR2_X1 U543 ( .A(n407), .B(n406), .ZN(n700) );
  NAND2_X1 U544 ( .A1(n704), .A2(G217), .ZN(n407) );
  NOR2_X2 U545 ( .A1(n677), .A2(n710), .ZN(n679) );
  NAND2_X2 U546 ( .A1(n371), .A2(n368), .ZN(n631) );
  NAND2_X1 U547 ( .A1(n409), .A2(n425), .ZN(n594) );
  XNOR2_X1 U548 ( .A(n414), .B(KEYINPUT77), .ZN(n409) );
  XNOR2_X2 U549 ( .A(n411), .B(KEYINPUT33), .ZN(n750) );
  XNOR2_X1 U550 ( .A(n413), .B(n707), .ZN(n708) );
  NAND2_X1 U551 ( .A1(n415), .A2(n640), .ZN(n414) );
  NOR2_X1 U552 ( .A1(n680), .A2(G902), .ZN(n519) );
  XNOR2_X1 U553 ( .A(n516), .B(n417), .ZN(n680) );
  XNOR2_X1 U554 ( .A(n418), .B(n453), .ZN(n417) );
  XNOR2_X1 U555 ( .A(n513), .B(n512), .ZN(n418) );
  INV_X1 U556 ( .A(n606), .ZN(n419) );
  NAND2_X1 U557 ( .A1(n425), .A2(n568), .ZN(n569) );
  NAND2_X1 U558 ( .A1(n425), .A2(n640), .ZN(n588) );
  OR2_X1 U559 ( .A1(n552), .A2(n660), .ZN(n429) );
  NAND2_X1 U560 ( .A1(n674), .A2(n552), .ZN(n431) );
  NAND2_X1 U561 ( .A1(n432), .A2(n715), .ZN(n716) );
  INV_X1 U562 ( .A(n636), .ZN(n434) );
  NAND2_X1 U563 ( .A1(n438), .A2(n614), .ZN(n437) );
  XNOR2_X1 U564 ( .A(n613), .B(KEYINPUT47), .ZN(n438) );
  XNOR2_X1 U565 ( .A(n766), .B(KEYINPUT93), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n544), .A2(n489), .ZN(n441) );
  XNOR2_X2 U567 ( .A(n587), .B(n586), .ZN(n640) );
  XNOR2_X2 U568 ( .A(n574), .B(KEYINPUT101), .ZN(n625) );
  AND2_X2 U569 ( .A1(n609), .A2(n608), .ZN(n621) );
  OR2_X2 U570 ( .A1(n446), .A2(n648), .ZN(n445) );
  XNOR2_X1 U571 ( .A(n582), .B(KEYINPUT94), .ZN(n446) );
  AND2_X1 U572 ( .A1(n734), .A2(n565), .ZN(n452) );
  XOR2_X1 U573 ( .A(n515), .B(n514), .Z(n453) );
  INV_X1 U574 ( .A(KEYINPUT48), .ZN(n629) );
  XNOR2_X1 U575 ( .A(n517), .B(G475), .ZN(n518) );
  XNOR2_X1 U576 ( .A(n658), .B(KEYINPUT45), .ZN(n661) );
  INV_X1 U577 ( .A(KEYINPUT14), .ZN(n455) );
  XNOR2_X1 U578 ( .A(n456), .B(n455), .ZN(n559) );
  NAND2_X1 U579 ( .A1(G953), .A2(G902), .ZN(n457) );
  NOR2_X1 U580 ( .A1(n559), .A2(n457), .ZN(n458) );
  XNOR2_X1 U581 ( .A(n458), .B(KEYINPUT107), .ZN(n459) );
  NOR2_X1 U582 ( .A1(G900), .A2(n459), .ZN(n461) );
  NAND2_X1 U583 ( .A1(n770), .A2(G952), .ZN(n557) );
  NOR2_X1 U584 ( .A1(n559), .A2(n557), .ZN(n460) );
  NOR2_X1 U585 ( .A1(n461), .A2(n460), .ZN(n599) );
  XNOR2_X2 U586 ( .A(G128), .B(KEYINPUT65), .ZN(n463) );
  XNOR2_X2 U587 ( .A(n463), .B(n462), .ZN(n526) );
  XOR2_X2 U588 ( .A(KEYINPUT68), .B(G131), .Z(n509) );
  XNOR2_X1 U589 ( .A(n509), .B(n465), .ZN(n466) );
  XNOR2_X1 U590 ( .A(n468), .B(n467), .ZN(n470) );
  NOR2_X1 U591 ( .A1(G953), .A2(G237), .ZN(n507) );
  NAND2_X1 U592 ( .A1(n507), .A2(G210), .ZN(n469) );
  XNOR2_X1 U593 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U594 ( .A(n472), .B(n537), .ZN(n473) );
  XNOR2_X1 U595 ( .A(n486), .B(n473), .ZN(n666) );
  INV_X1 U596 ( .A(G902), .ZN(n532) );
  NAND2_X1 U597 ( .A1(n666), .A2(n532), .ZN(n475) );
  INV_X1 U598 ( .A(G472), .ZN(n474) );
  XNOR2_X2 U599 ( .A(n475), .B(n474), .ZN(n587) );
  INV_X1 U600 ( .A(G237), .ZN(n476) );
  NAND2_X1 U601 ( .A1(n532), .A2(n476), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n549), .A2(G214), .ZN(n478) );
  INV_X1 U603 ( .A(KEYINPUT90), .ZN(n477) );
  XNOR2_X1 U604 ( .A(n478), .B(n477), .ZN(n732) );
  NOR2_X1 U605 ( .A1(n587), .A2(n732), .ZN(n479) );
  NAND2_X1 U606 ( .A1(G227), .A2(n770), .ZN(n480) );
  XNOR2_X1 U607 ( .A(n491), .B(n480), .ZN(n484) );
  XNOR2_X1 U608 ( .A(n481), .B(G110), .ZN(n483) );
  XNOR2_X1 U609 ( .A(G101), .B(KEYINPUT75), .ZN(n482) );
  XNOR2_X1 U610 ( .A(n483), .B(n482), .ZN(n538) );
  XOR2_X1 U611 ( .A(n484), .B(n538), .Z(n485) );
  XNOR2_X1 U612 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n487) );
  XNOR2_X1 U613 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U614 ( .A(n494), .B(KEYINPUT23), .Z(n497) );
  XNOR2_X1 U615 ( .A(KEYINPUT8), .B(n495), .ZN(n527) );
  NAND2_X1 U616 ( .A1(n527), .A2(G221), .ZN(n496) );
  XNOR2_X1 U617 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U618 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n502) );
  XNOR2_X1 U619 ( .A(G902), .B(KEYINPUT15), .ZN(n548) );
  NAND2_X1 U620 ( .A1(G234), .A2(n548), .ZN(n500) );
  XNOR2_X1 U621 ( .A(KEYINPUT20), .B(n500), .ZN(n504) );
  AND2_X1 U622 ( .A1(G217), .A2(n504), .ZN(n501) );
  XNOR2_X1 U623 ( .A(n502), .B(n501), .ZN(n503) );
  AND2_X1 U624 ( .A1(n504), .A2(G221), .ZN(n506) );
  INV_X1 U625 ( .A(KEYINPUT21), .ZN(n505) );
  XNOR2_X1 U626 ( .A(n506), .B(n505), .ZN(n722) );
  INV_X1 U627 ( .A(n622), .ZN(n554) );
  NAND2_X1 U628 ( .A1(G214), .A2(n507), .ZN(n508) );
  XNOR2_X1 U629 ( .A(n509), .B(KEYINPUT97), .ZN(n513) );
  XOR2_X1 U630 ( .A(G140), .B(G104), .Z(n511) );
  XNOR2_X1 U631 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U632 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n517) );
  INV_X1 U633 ( .A(n573), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n521), .B(n520), .ZN(n525) );
  INV_X1 U635 ( .A(n526), .ZN(n529) );
  NAND2_X1 U636 ( .A1(n527), .A2(G217), .ZN(n528) );
  XNOR2_X1 U637 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U638 ( .A(n531), .B(n530), .ZN(n702) );
  NAND2_X1 U639 ( .A1(n702), .A2(n532), .ZN(n533) );
  XNOR2_X1 U640 ( .A(n533), .B(G478), .ZN(n577) );
  INV_X1 U641 ( .A(n577), .ZN(n534) );
  OR2_X1 U642 ( .A1(n573), .A2(n534), .ZN(n643) );
  XNOR2_X1 U643 ( .A(n535), .B(G122), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n537), .B(n536), .ZN(n539) );
  XNOR2_X1 U645 ( .A(n539), .B(n538), .ZN(n693) );
  XNOR2_X1 U646 ( .A(n540), .B(KEYINPUT88), .ZN(n542) );
  XNOR2_X1 U647 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U648 ( .A(n543), .B(n544), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U650 ( .A(n693), .B(n547), .ZN(n674) );
  NAND2_X1 U651 ( .A1(n549), .A2(G210), .ZN(n551) );
  INV_X1 U652 ( .A(KEYINPUT89), .ZN(n550) );
  XNOR2_X1 U653 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U654 ( .A1(n643), .A2(n633), .ZN(n553) );
  NAND2_X1 U655 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U656 ( .A1(n623), .A2(n555), .ZN(n605) );
  XOR2_X1 U657 ( .A(n605), .B(G143), .Z(G45) );
  INV_X1 U658 ( .A(n570), .ZN(n590) );
  BUF_X2 U659 ( .A(n587), .Z(n725) );
  NAND2_X1 U660 ( .A1(n725), .A2(n408), .ZN(n556) );
  NOR2_X1 U661 ( .A1(n718), .A2(n556), .ZN(n568) );
  XOR2_X1 U662 ( .A(G898), .B(KEYINPUT91), .Z(n689) );
  NOR2_X1 U663 ( .A1(n689), .A2(n770), .ZN(n694) );
  NAND2_X1 U664 ( .A1(n694), .A2(G902), .ZN(n558) );
  NAND2_X1 U665 ( .A1(n558), .A2(n557), .ZN(n560) );
  INV_X1 U666 ( .A(n559), .ZN(n746) );
  AND2_X1 U667 ( .A1(n560), .A2(n746), .ZN(n561) );
  INV_X1 U668 ( .A(KEYINPUT0), .ZN(n562) );
  XNOR2_X2 U669 ( .A(n563), .B(n562), .ZN(n580) );
  NOR2_X1 U670 ( .A1(n564), .A2(n577), .ZN(n734) );
  INV_X1 U671 ( .A(n722), .ZN(n565) );
  XOR2_X1 U672 ( .A(KEYINPUT67), .B(KEYINPUT22), .Z(n566) );
  XNOR2_X1 U673 ( .A(n645), .B(G110), .ZN(G12) );
  NOR2_X1 U674 ( .A1(n639), .A2(n725), .ZN(n729) );
  NAND2_X1 U675 ( .A1(n729), .A2(n580), .ZN(n572) );
  XNOR2_X1 U676 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n571) );
  XNOR2_X1 U677 ( .A(n572), .B(n571), .ZN(n648) );
  INV_X1 U678 ( .A(KEYINPUT106), .ZN(n575) );
  NAND2_X1 U679 ( .A1(n648), .A2(n368), .ZN(n576) );
  XNOR2_X1 U680 ( .A(n576), .B(G113), .ZN(G15) );
  AND2_X1 U681 ( .A1(n573), .A2(n577), .ZN(n758) );
  NAND2_X1 U682 ( .A1(n648), .A2(n758), .ZN(n579) );
  XNOR2_X1 U683 ( .A(G116), .B(KEYINPUT116), .ZN(n578) );
  XNOR2_X1 U684 ( .A(n579), .B(n578), .ZN(G18) );
  XNOR2_X1 U685 ( .A(n580), .B(KEYINPUT92), .ZN(n641) );
  INV_X1 U686 ( .A(n641), .ZN(n581) );
  NAND2_X1 U687 ( .A1(n647), .A2(n758), .ZN(n585) );
  XOR2_X1 U688 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n583) );
  XNOR2_X1 U689 ( .A(n583), .B(G107), .ZN(n584) );
  XNOR2_X1 U690 ( .A(n585), .B(n584), .ZN(G9) );
  XOR2_X1 U691 ( .A(KEYINPUT102), .B(KEYINPUT6), .Z(n586) );
  XNOR2_X1 U692 ( .A(n588), .B(KEYINPUT84), .ZN(n592) );
  INV_X1 U693 ( .A(n408), .ZN(n589) );
  NAND2_X1 U694 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U695 ( .A1(n592), .A2(n591), .ZN(n650) );
  XOR2_X1 U696 ( .A(G101), .B(n650), .Z(G3) );
  XNOR2_X1 U697 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n593) );
  XOR2_X1 U698 ( .A(G119), .B(KEYINPUT127), .Z(n595) );
  XNOR2_X1 U699 ( .A(n646), .B(n595), .ZN(G21) );
  XNOR2_X1 U700 ( .A(G104), .B(KEYINPUT113), .ZN(n597) );
  NAND2_X1 U701 ( .A1(n647), .A2(n368), .ZN(n596) );
  XOR2_X1 U702 ( .A(n597), .B(n596), .Z(G6) );
  NOR2_X1 U703 ( .A1(n722), .A2(n599), .ZN(n600) );
  XNOR2_X1 U704 ( .A(KEYINPUT70), .B(n601), .ZN(n606) );
  XNOR2_X2 U705 ( .A(n603), .B(KEYINPUT112), .ZN(n778) );
  XNOR2_X1 U706 ( .A(n778), .B(n604), .ZN(n619) );
  INV_X1 U707 ( .A(n605), .ZN(n612) );
  NOR2_X2 U708 ( .A1(n606), .A2(n725), .ZN(n607) );
  XNOR2_X1 U709 ( .A(n607), .B(KEYINPUT28), .ZN(n608) );
  AND2_X2 U710 ( .A1(n621), .A2(n610), .ZN(n762) );
  NAND2_X1 U711 ( .A1(n762), .A2(KEYINPUT79), .ZN(n611) );
  NAND2_X1 U712 ( .A1(n612), .A2(n611), .ZN(n616) );
  OR2_X1 U713 ( .A1(n625), .A2(n758), .ZN(n736) );
  NAND2_X1 U714 ( .A1(n762), .A2(n736), .ZN(n613) );
  INV_X1 U715 ( .A(KEYINPUT79), .ZN(n614) );
  NAND2_X1 U716 ( .A1(KEYINPUT47), .A2(n736), .ZN(n615) );
  XNOR2_X1 U717 ( .A(KEYINPUT74), .B(n617), .ZN(n618) );
  NOR2_X1 U718 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U719 ( .A1(n734), .A2(n737), .ZN(n620) );
  NAND2_X1 U720 ( .A1(n637), .A2(n625), .ZN(n626) );
  XNOR2_X1 U721 ( .A(n630), .B(n629), .ZN(n636) );
  NOR2_X1 U722 ( .A1(n732), .A2(n631), .ZN(n632) );
  AND2_X1 U723 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U724 ( .A(n635), .B(KEYINPUT110), .ZN(n777) );
  XNOR2_X1 U725 ( .A(n638), .B(KEYINPUT81), .ZN(n659) );
  INV_X1 U726 ( .A(KEYINPUT34), .ZN(n642) );
  INV_X1 U727 ( .A(n643), .ZN(n644) );
  INV_X1 U728 ( .A(n736), .ZN(n649) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(KEYINPUT85), .ZN(n657) );
  OR2_X1 U732 ( .A1(n655), .A2(KEYINPUT44), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n658) );
  BUF_X2 U734 ( .A(n661), .Z(n712) );
  INV_X1 U735 ( .A(n661), .ZN(n662) );
  NOR2_X1 U736 ( .A1(n663), .A2(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U737 ( .A1(n698), .A2(G472), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT62), .ZN(n667) );
  XNOR2_X1 U739 ( .A(n668), .B(n667), .ZN(n670) );
  INV_X1 U740 ( .A(n710), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n672), .B(n671), .ZN(G57) );
  NAND2_X1 U744 ( .A1(n698), .A2(G210), .ZN(n676) );
  XOR2_X1 U745 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U747 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U748 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n679), .B(n678), .ZN(G51) );
  NAND2_X1 U750 ( .A1(n698), .A2(G475), .ZN(n682) );
  XNOR2_X1 U751 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(G60) );
  XOR2_X1 U753 ( .A(G122), .B(KEYINPUT126), .Z(n687) );
  XNOR2_X1 U754 ( .A(n686), .B(n687), .ZN(G24) );
  NAND2_X1 U755 ( .A1(n712), .A2(n770), .ZN(n692) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n688) );
  XNOR2_X1 U757 ( .A(KEYINPUT61), .B(n688), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n697) );
  INV_X1 U760 ( .A(n693), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n697), .B(n696), .ZN(G69) );
  NOR2_X1 U763 ( .A1(n700), .A2(n710), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n704), .A2(G478), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n703), .A2(n710), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n704), .A2(G469), .ZN(n709) );
  XNOR2_X1 U767 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n706) );
  XNOR2_X1 U768 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U770 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(G54) );
  NOR2_X1 U772 ( .A1(n712), .A2(KEYINPUT2), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n713), .B(KEYINPUT80), .ZN(n717) );
  INV_X1 U774 ( .A(KEYINPUT2), .ZN(n714) );
  OR2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n755) );
  XNOR2_X1 U776 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n454), .A2(n718), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n720), .B(n719), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n722), .A2(n408), .ZN(n723) );
  XOR2_X1 U780 ( .A(KEYINPUT49), .B(n723), .Z(n724) );
  NAND2_X1 U781 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U782 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U783 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U784 ( .A(n730), .B(KEYINPUT51), .ZN(n731) );
  NAND2_X1 U785 ( .A1(n731), .A2(n749), .ZN(n744) );
  NAND2_X1 U786 ( .A1(n733), .A2(n732), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U789 ( .A(KEYINPUT119), .B(n738), .Z(n739) );
  NAND2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U791 ( .A(KEYINPUT120), .B(n741), .ZN(n742) );
  NAND2_X1 U792 ( .A1(n742), .A2(n750), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U794 ( .A(KEYINPUT52), .B(n745), .Z(n748) );
  NAND2_X1 U795 ( .A1(n746), .A2(G952), .ZN(n747) );
  NOR2_X1 U796 ( .A1(n748), .A2(n747), .ZN(n753) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(n770), .ZN(n752) );
  NOR2_X1 U799 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U801 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n756) );
  XNOR2_X1 U802 ( .A(n757), .B(n756), .ZN(G75) );
  XOR2_X1 U803 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n760) );
  NAND2_X1 U804 ( .A1(n762), .A2(n758), .ZN(n759) );
  XNOR2_X1 U805 ( .A(n760), .B(n759), .ZN(n761) );
  XNOR2_X1 U806 ( .A(G128), .B(n761), .ZN(G30) );
  AND2_X1 U807 ( .A1(n762), .A2(n368), .ZN(n764) );
  XNOR2_X1 U808 ( .A(G146), .B(KEYINPUT115), .ZN(n763) );
  XNOR2_X1 U809 ( .A(n764), .B(n763), .ZN(G48) );
  XNOR2_X1 U810 ( .A(G134), .B(n765), .ZN(G36) );
  XNOR2_X1 U811 ( .A(n767), .B(n766), .ZN(n772) );
  INV_X1 U812 ( .A(n772), .ZN(n768) );
  XNOR2_X1 U813 ( .A(n769), .B(n768), .ZN(n771) );
  NAND2_X1 U814 ( .A1(n771), .A2(n770), .ZN(n776) );
  XNOR2_X1 U815 ( .A(G227), .B(n772), .ZN(n773) );
  NAND2_X1 U816 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U817 ( .A1(n774), .A2(G953), .ZN(n775) );
  NAND2_X1 U818 ( .A1(n776), .A2(n775), .ZN(G72) );
  XOR2_X1 U819 ( .A(G140), .B(n777), .Z(G42) );
  XNOR2_X1 U820 ( .A(n778), .B(KEYINPUT117), .ZN(n779) );
  XNOR2_X1 U821 ( .A(n779), .B(KEYINPUT37), .ZN(n780) );
  XNOR2_X1 U822 ( .A(G125), .B(n780), .ZN(G27) );
  XNOR2_X1 U823 ( .A(G137), .B(n781), .ZN(G39) );
  XNOR2_X1 U824 ( .A(n782), .B(G131), .ZN(G33) );
endmodule

