//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141, new_n1143,
    new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n449), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n462));
  AOI211_X1 g037(.A(new_n461), .B(new_n462), .C1(new_n455), .C2(G2106), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT68), .B(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AOI21_X1  g050(.A(G2105), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n465), .A2(new_n480), .A3(G125), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n477), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n476), .A2(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n472), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n472), .A2(new_n477), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n485), .B1(new_n486), .B2(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND2_X1  g066(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .A4(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n472), .B2(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT4), .B1(new_n498), .B2(new_n477), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n465), .A2(new_n480), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(G138), .A3(new_n477), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(KEYINPUT69), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT70), .Z(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G88), .B1(new_n516), .B2(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  AND2_X1   g094(.A1(new_n514), .A2(G89), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n521), .B(new_n523), .C1(new_n524), .C2(new_n515), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n520), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n509), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n513), .A2(new_n530), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G171));
  AOI22_X1  g108(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n509), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n514), .A2(G81), .B1(new_n516), .B2(G43), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n537), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n535), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  AOI22_X1  g122(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n509), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n516), .A2(KEYINPUT9), .A3(G53), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n515), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n507), .A2(KEYINPUT72), .A3(new_n512), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT72), .B1(new_n507), .B2(new_n512), .ZN(new_n557));
  OAI21_X1  g132(.A(G91), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n558), .A2(KEYINPUT73), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(new_n555), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n560), .B1(new_n562), .B2(G91), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n549), .B(new_n554), .C1(new_n559), .C2(new_n563), .ZN(G299));
  XOR2_X1   g139(.A(G171), .B(KEYINPUT74), .Z(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G301));
  NAND2_X1  g141(.A1(new_n562), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n516), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(new_n562), .A2(G86), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n505), .B2(new_n506), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT76), .B(G651), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n571), .A2(new_n572), .A3(new_n578), .A4(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n509), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n513), .A2(new_n585), .B1(new_n515), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(new_n562), .A2(G92), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n507), .A2(G66), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n509), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(G54), .B2(new_n516), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT77), .B1(new_n598), .B2(G868), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n565), .A2(new_n600), .ZN(new_n601));
  MUX2_X1   g176(.A(new_n599), .B(KEYINPUT77), .S(new_n601), .Z(G284));
  MUX2_X1   g177(.A(new_n599), .B(KEYINPUT77), .S(new_n601), .Z(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n608), .B2(G860), .ZN(G148));
  INV_X1    g184(.A(new_n540), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n610), .A2(new_n538), .B1(new_n509), .B2(new_n534), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n600), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n597), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(new_n489), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G135), .ZN(new_n617));
  INV_X1    g192(.A(new_n486), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(new_n477), .B2(G111), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n617), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND3_X1  g198(.A1(new_n500), .A2(new_n477), .A3(new_n474), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT13), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2443), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2446), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n643), .A2(G14), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n645), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2100), .Z(new_n652));
  AND2_X1   g227(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n647), .A2(new_n648), .ZN(new_n654));
  AOI21_X1  g229(.A(KEYINPUT18), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT81), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  AOI22_X1  g240(.A1(new_n663), .A2(new_n664), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OR3_X1    g241(.A1(new_n660), .A2(new_n665), .A3(new_n662), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n666), .B(new_n667), .C1(new_n664), .C2(new_n663), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT22), .B(G1981), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(G1971), .Z(new_n679));
  NOR2_X1   g254(.A1(G16), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(G16), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT33), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n676), .A2(G6), .ZN(new_n685));
  INV_X1    g260(.A(G305), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n676), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT32), .B(G1981), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n679), .A2(new_n684), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n676), .A2(G24), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n588), .B2(new_n676), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT82), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT36), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n618), .A2(G119), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n616), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(new_n477), .B2(G107), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G25), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT35), .B(G1991), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n697), .B2(KEYINPUT36), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G35), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G162), .B2(new_n710), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT29), .Z(new_n713));
  INV_X1    g288(.A(G2090), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT94), .Z(new_n716));
  NOR2_X1   g291(.A1(G16), .A2(G19), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n541), .B2(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G1341), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(G1341), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n676), .A2(KEYINPUT23), .A3(G20), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n723));
  INV_X1    g298(.A(G20), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n725), .C1(new_n605), .C2(new_n676), .ZN(new_n726));
  INV_X1    g301(.A(G1956), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(KEYINPUT24), .A2(G34), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n710), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n710), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2084), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n720), .A2(new_n721), .A3(new_n728), .A4(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G5), .A2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G171), .B2(G16), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n710), .A2(G33), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n616), .A2(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n500), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(new_n477), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n743));
  NAND3_X1  g318(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n740), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n710), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT86), .B(G2072), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT90), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n710), .B1(new_n753), .B2(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT91), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(G28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(KEYINPUT91), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n755), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n750), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n710), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n763), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n764));
  INV_X1    g339(.A(G128), .ZN(new_n765));
  INV_X1    g340(.A(G140), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n764), .B1(new_n486), .B2(new_n765), .C1(new_n766), .C2(new_n489), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n710), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT84), .B(G2067), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n616), .A2(G141), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT87), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n474), .A2(G105), .A3(new_n477), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT26), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n774), .B(new_n776), .C1(new_n618), .C2(G129), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G32), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n771), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n713), .A2(new_n714), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n759), .B(new_n782), .C1(KEYINPUT93), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n785));
  NOR2_X1   g360(.A1(G27), .A2(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G164), .B2(G29), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT92), .B(G2078), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n784), .B(new_n790), .C1(new_n710), .C2(new_n622), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n735), .A2(new_n738), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n780), .A2(new_n781), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT88), .Z(new_n794));
  NOR2_X1   g369(.A1(new_n697), .A2(KEYINPUT36), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n699), .B2(new_n707), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n709), .A2(new_n792), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n676), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n676), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT89), .B(G1966), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NOR2_X1   g376(.A1(new_n598), .A2(new_n676), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G4), .B2(new_n676), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1348), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n797), .A2(new_n801), .A3(new_n805), .ZN(G311));
  AND3_X1   g381(.A1(new_n709), .A2(new_n792), .A3(new_n796), .ZN(new_n807));
  INV_X1    g382(.A(new_n801), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n807), .A2(new_n808), .A3(new_n804), .A4(new_n794), .ZN(G150));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n513), .A2(new_n810), .B1(new_n515), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(new_n509), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n541), .B(new_n816), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n598), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT96), .Z(new_n824));
  INV_X1    g399(.A(G860), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n818), .B1(new_n824), .B2(new_n826), .ZN(G145));
  OAI211_X1 g402(.A(G126), .B(new_n465), .C1(new_n474), .C2(new_n464), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n477), .B1(new_n828), .B2(new_n496), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT4), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n501), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n493), .A2(new_n494), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n477), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n767), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n778), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n746), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n618), .A2(G130), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n616), .A2(G142), .ZN(new_n841));
  NOR2_X1   g416(.A1(G106), .A2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n704), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n626), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n836), .A2(new_n747), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n836), .A2(new_n747), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT98), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n839), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n846), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n837), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n490), .B(KEYINPUT97), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n732), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n622), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n839), .A2(new_n849), .A3(KEYINPUT99), .A4(new_n846), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n852), .A2(new_n854), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n837), .B(new_n853), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n857), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(G303), .B(G288), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(G290), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(G290), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G305), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n686), .A3(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n819), .B(new_n613), .Z(new_n874));
  AOI21_X1  g449(.A(new_n597), .B1(new_n605), .B2(KEYINPUT100), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(KEYINPUT100), .B2(new_n605), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n597), .A2(new_n877), .A3(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(KEYINPUT41), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n874), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n873), .A2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(G868), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n816), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(G868), .B2(new_n886), .ZN(G295));
  OAI21_X1  g462(.A(new_n885), .B1(G868), .B2(new_n886), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  AND2_X1   g464(.A1(G286), .A2(G171), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(G301), .B2(G168), .ZN(new_n891));
  XOR2_X1   g466(.A(new_n819), .B(new_n891), .Z(new_n892));
  NOR2_X1   g467(.A1(new_n879), .A2(KEYINPUT41), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n876), .B2(new_n878), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n892), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n819), .B(new_n891), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n878), .A3(new_n876), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n870), .A2(new_n871), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n861), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n904));
  OR3_X1    g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n895), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n892), .B(new_n907), .C1(new_n881), .C2(new_n906), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n872), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n909), .B2(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n889), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n909), .A2(new_n903), .A3(new_n904), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n904), .B1(new_n902), .B2(new_n903), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT103), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n916), .B2(new_n912), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n917), .B2(new_n889), .ZN(G397));
  NOR2_X1   g493(.A1(new_n611), .A2(KEYINPUT120), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n921));
  AOI21_X1  g496(.A(G1384), .B1(new_n831), .B2(new_n833), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT45), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n479), .A2(new_n481), .ZN(new_n925));
  OAI21_X1  g500(.A(G40), .B1(new_n925), .B2(new_n477), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n476), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G40), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n482), .A2(new_n928), .ZN(new_n929));
  AOI22_X1  g504(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n929), .B(KEYINPUT104), .C1(G2105), .C2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G1996), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n921), .A2(new_n923), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n922), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT118), .B(G1341), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT58), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT119), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n933), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n933), .B2(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n919), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT59), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT59), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(new_n919), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n550), .A2(KEYINPUT115), .A3(new_n553), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT57), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(G299), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n558), .B(KEYINPUT73), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(new_n549), .A3(new_n554), .A4(new_n949), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT56), .B(G2072), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n921), .A2(new_n934), .A3(new_n923), .A4(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n927), .A2(new_n931), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n954), .B(new_n956), .C1(new_n961), .C2(G1956), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT116), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n956), .B1(new_n961), .B2(G1956), .ZN(new_n965));
  INV_X1    g540(.A(new_n954), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n958), .B(G1384), .C1(new_n831), .C2(new_n833), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n934), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n727), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(KEYINPUT116), .A3(new_n954), .A4(new_n956), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n967), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n962), .A2(KEYINPUT61), .ZN(new_n976));
  AOI211_X1 g551(.A(KEYINPUT117), .B(new_n954), .C1(new_n971), .C2(new_n956), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n965), .B2(new_n966), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n946), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT121), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n946), .A2(new_n975), .A3(KEYINPUT121), .A4(new_n980), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n935), .A2(G2067), .ZN(new_n985));
  INV_X1    g560(.A(G1348), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(new_n970), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(new_n598), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(KEYINPUT60), .B2(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n983), .A2(new_n984), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n977), .A2(new_n979), .B1(new_n597), .B2(new_n987), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n964), .A3(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n921), .A2(new_n934), .A3(new_n923), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G2078), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n921), .A2(KEYINPUT108), .A3(new_n923), .A4(new_n934), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1961), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n970), .A2(KEYINPUT123), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT123), .B1(new_n970), .B2(new_n1003), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n476), .B(KEYINPUT124), .Z(new_n1007));
  NAND3_X1  g582(.A1(new_n921), .A2(new_n929), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT125), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n923), .B1(KEYINPUT126), .B2(new_n998), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n1001), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT125), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n921), .A2(new_n1013), .A3(new_n1007), .A4(new_n929), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1002), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G171), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT127), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n961), .A2(G1961), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n995), .A2(new_n1001), .A3(G2078), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n1021), .B(new_n1022), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(G301), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1016), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1002), .A2(new_n1006), .A3(G301), .A4(new_n1015), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1023), .B2(G301), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G286), .A2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  INV_X1    g607(.A(G1966), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1032), .A2(new_n961), .B1(new_n995), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  OAI221_X1 g610(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n995), .A2(new_n1033), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G2084), .B2(new_n970), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(new_n1038), .C1(new_n1040), .C2(G286), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(G8), .A3(G286), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1028), .A2(new_n1020), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n997), .B2(new_n999), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n961), .A2(new_n714), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G303), .A2(G8), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1051), .B(G8), .C1(new_n1045), .C2(new_n1047), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1035), .B1(new_n934), .B2(new_n922), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n681), .A2(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1056), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n581), .A2(new_n578), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT110), .B(G1981), .Z(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1062), .A2(new_n571), .A3(new_n572), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n507), .A2(G86), .A3(new_n512), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n572), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT111), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1069), .A3(new_n572), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n581), .A3(new_n578), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(G1981), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1065), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1065), .A2(new_n1072), .A3(new_n1073), .A4(KEYINPUT49), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n1056), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(KEYINPUT113), .A3(new_n1056), .A4(new_n1078), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1058), .B(new_n1061), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1053), .A2(new_n1054), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1026), .A2(new_n1044), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n994), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1087), .A2(KEYINPUT62), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1023), .A2(G301), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(KEYINPUT62), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1088), .A2(new_n1084), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1083), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1093));
  NOR2_X1   g668(.A1(G288), .A2(G1976), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n686), .B2(new_n1064), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1056), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1092), .A2(new_n1054), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1034), .A2(new_n1035), .A3(G286), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1053), .A2(new_n1083), .A3(new_n1054), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1098), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1086), .A2(new_n1091), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n778), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n921), .A2(new_n957), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(G1996), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT105), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n767), .B(G2067), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT106), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1110), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT107), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(G1996), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1112), .B(new_n1117), .C1(new_n778), .C2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n704), .B(new_n706), .Z(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n588), .B(new_n694), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1108), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1110), .A2(new_n694), .A3(new_n588), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n1125), .B(KEYINPUT48), .Z(new_n1126));
  NOR2_X1   g701(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n704), .A2(new_n706), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1119), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n767), .A2(G2067), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1115), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1118), .A2(KEYINPUT46), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1115), .B1(new_n1114), .B2(new_n778), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1118), .A2(KEYINPUT46), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT47), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1127), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1124), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g713(.A1(G401), .A2(G227), .ZN(new_n1140));
  NAND3_X1  g714(.A1(new_n864), .A2(G319), .A3(new_n1140), .ZN(new_n1141));
  NOR3_X1   g715(.A1(new_n917), .A2(new_n1141), .A3(G229), .ZN(G308));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1143));
  INV_X1    g717(.A(new_n912), .ZN(new_n1144));
  NAND3_X1  g718(.A1(new_n1144), .A2(KEYINPUT103), .A3(new_n915), .ZN(new_n1145));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n674), .A3(new_n1145), .A4(new_n914), .ZN(G225));
endmodule


