//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(G125), .B(G140), .ZN(new_n194));
  MUX2_X1   g008(.A(new_n193), .B(new_n194), .S(KEYINPUT16), .Z(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n194), .A2(new_n196), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G128), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G110), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n201), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n209), .A2(KEYINPUT76), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT76), .B1(new_n209), .B2(new_n212), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n199), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT77), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n199), .B(KEYINPUT77), .C1(new_n213), .C2(new_n214), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(new_n208), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT75), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n195), .B(G146), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n210), .A2(new_n211), .ZN(new_n223));
  OR3_X1    g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(KEYINPUT70), .A2(G953), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT70), .A2(G953), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n219), .B2(new_n224), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n191), .B1(new_n233), .B2(new_n188), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n219), .A2(new_n224), .ZN(new_n235));
  INV_X1    g049(.A(new_n230), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n219), .A2(new_n224), .A3(new_n230), .ZN(new_n238));
  AND4_X1   g052(.A1(new_n188), .A2(new_n237), .A3(new_n238), .A4(new_n191), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n189), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n189), .A2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n227), .A2(G210), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n246));
  XNOR2_X1  g060(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G137), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT11), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n254), .B2(G137), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n258), .A2(new_n253), .A3(new_n261), .A4(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n262), .A2(new_n263), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n260), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT0), .B(G128), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT65), .A3(G146), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(new_n269), .B2(G146), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT64), .B1(new_n269), .B2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT64), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n196), .A3(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n268), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G143), .B(G146), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT0), .A3(G128), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT66), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n272), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n277), .A2(new_n283), .A3(new_n270), .ZN(new_n284));
  INV_X1    g098(.A(new_n268), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n280), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n267), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n196), .A2(G143), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n200), .B1(new_n290), .B2(KEYINPUT1), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(G146), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n252), .A2(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n255), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n293), .A2(new_n296), .B1(G131), .B2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n261), .A4(new_n258), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n264), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g117(.A(G116), .B(G119), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n306), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n304), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n278), .A2(new_n281), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n299), .A2(new_n301), .B1(new_n267), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n310), .B(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n251), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n298), .A2(G131), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n291), .B1(new_n273), .B2(new_n277), .ZN(new_n320));
  INV_X1    g134(.A(new_n296), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n301), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n300), .A2(new_n264), .B1(new_n259), .B2(G131), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n286), .A2(new_n280), .ZN(new_n325));
  OAI22_X1  g139(.A1(new_n322), .A2(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT28), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n250), .B1(new_n318), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n333), .B(new_n250), .C1(new_n318), .C2(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT30), .B1(new_n289), .B2(new_n302), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n336), .A2(KEYINPUT68), .B1(KEYINPUT30), .B2(new_n313), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n303), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n341), .A3(new_n310), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(new_n317), .A3(new_n249), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(KEYINPUT31), .A3(new_n317), .A4(new_n249), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n335), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT32), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n335), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n346), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT32), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n348), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n326), .B(new_n316), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n359), .A2(new_n330), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n249), .A2(KEYINPUT29), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n188), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n342), .A2(new_n317), .A3(new_n250), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n249), .B1(new_n318), .B2(new_n330), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G472), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n243), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n227), .A2(G227), .ZN(new_n368));
  XOR2_X1   g182(.A(G110), .B(G140), .Z(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G107), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n372), .B2(G104), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT80), .B1(new_n374), .B2(G107), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n374), .A3(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n372), .A3(G104), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n375), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G101), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n372), .A2(G104), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(G107), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT3), .B1(new_n384), .B2(KEYINPUT79), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n372), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(G104), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n383), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n296), .B1(new_n291), .B2(new_n279), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT82), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n381), .A2(new_n388), .A3(new_n392), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n388), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT83), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n381), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n293), .A2(new_n296), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n267), .ZN(new_n402));
  XOR2_X1   g216(.A(new_n402), .B(KEYINPUT12), .Z(new_n403));
  INV_X1    g217(.A(KEYINPUT10), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n293), .B2(new_n296), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n381), .A2(new_n388), .A3(new_n397), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(new_n381), .B2(new_n388), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT84), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n405), .B(new_n410), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n372), .A2(KEYINPUT79), .A3(G104), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT3), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n382), .B1(new_n416), .B2(new_n386), .ZN(new_n417));
  INV_X1    g231(.A(G101), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n386), .ZN(new_n420));
  INV_X1    g234(.A(new_n382), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n422), .A2(G101), .B1(new_n420), .B2(new_n383), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n419), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n394), .A2(new_n404), .B1(new_n424), .B2(new_n312), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n324), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n412), .A2(new_n425), .A3(KEYINPUT85), .A4(new_n324), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n371), .B1(new_n403), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n371), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n324), .B1(new_n412), .B2(new_n425), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n370), .B1(new_n428), .B2(new_n429), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n435), .B1(new_n436), .B2(KEYINPUT86), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n431), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G469), .B1(new_n438), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT87), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT87), .B(G469), .C1(new_n438), .C2(G902), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n436), .A2(new_n403), .ZN(new_n444));
  INV_X1    g258(.A(new_n435), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n371), .B1(new_n430), .B2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n443), .B(new_n188), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT9), .B(G234), .ZN(new_n449));
  OAI21_X1  g263(.A(G221), .B1(new_n449), .B2(G902), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT88), .B(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n205), .A2(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G113), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n454), .A2(KEYINPUT90), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n454), .A2(KEYINPUT90), .B1(KEYINPUT5), .B2(new_n304), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n455), .A2(new_n456), .B1(new_n304), .B2(new_n308), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n453), .B(G113), .C1(new_n305), .C2(new_n451), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n309), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n457), .A2(new_n399), .B1(new_n395), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(KEYINPUT89), .B(KEYINPUT8), .Z(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G224), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT7), .B1(new_n465), .B2(G953), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n325), .A2(G125), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n293), .A2(new_n192), .A3(new_n296), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n469), .A3(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT91), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n459), .B1(new_n396), .B2(new_n398), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n424), .A2(new_n310), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n462), .A3(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n468), .A2(new_n469), .A3(new_n467), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(new_n470), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(new_n481), .C1(new_n460), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n462), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n424), .A2(new_n310), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n478), .A3(KEYINPUT6), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(new_n484), .C1(new_n485), .C2(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n469), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n465), .A2(G953), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n487), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n483), .A2(new_n493), .A3(new_n188), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT92), .Z(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n483), .A2(new_n493), .A3(new_n188), .A4(new_n496), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G475), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n227), .A2(G143), .A3(G214), .A4(new_n244), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n225), .A2(G214), .A3(new_n244), .A4(new_n226), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n269), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT18), .A3(G131), .ZN(new_n507));
  NAND2_X1  g321(.A1(KEYINPUT18), .A2(G131), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n194), .A2(new_n196), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n507), .B(new_n509), .C1(new_n198), .C2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n261), .B1(new_n503), .B2(new_n505), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n222), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n261), .A3(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n516), .A2(KEYINPUT17), .A3(new_n512), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n511), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(G113), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n374), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n520), .B(new_n511), .C1(new_n514), .C2(new_n517), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n502), .B1(new_n524), .B2(new_n188), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n527));
  INV_X1    g341(.A(new_n523), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n516), .B2(new_n512), .ZN(new_n530));
  INV_X1    g344(.A(new_n512), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT94), .A3(new_n515), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n194), .B(KEYINPUT19), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n197), .B1(new_n196), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n520), .B1(new_n535), .B2(new_n511), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n527), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n528), .A2(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(KEYINPUT95), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n543), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n540), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n526), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G952), .ZN(new_n549));
  AOI211_X1 g363(.A(G953), .B(new_n549), .C1(G234), .C2(G237), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n188), .B(new_n227), .C1(G234), .C2(G237), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT21), .B(G898), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT101), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G478), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n449), .A2(new_n187), .A3(G953), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n200), .A2(G143), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n200), .B2(G143), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n269), .A2(KEYINPUT97), .A3(G128), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(KEYINPUT13), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT13), .B1(new_n565), .B2(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(G134), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n563), .A2(new_n254), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G116), .B(G122), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT96), .B(G107), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT99), .ZN(new_n577));
  INV_X1    g391(.A(G122), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G116), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n372), .B1(new_n579), .B2(KEYINPUT14), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(new_n573), .ZN(new_n581));
  INV_X1    g395(.A(new_n572), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n254), .B1(new_n563), .B2(new_n571), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n577), .B1(new_n576), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n560), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n584), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT99), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n559), .A3(new_n585), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n558), .B1(new_n592), .B2(new_n188), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n188), .A3(new_n558), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(KEYINPUT100), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n597));
  AOI211_X1 g411(.A(G902), .B(new_n557), .C1(new_n588), .C2(new_n591), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n597), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n555), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n501), .A2(new_n548), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n367), .A2(new_n448), .A3(new_n450), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND3_X1  g417(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n604), .A2(new_n555), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n592), .A2(new_n188), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(new_n556), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n592), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n588), .A2(new_n591), .A3(KEYINPUT33), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n556), .A2(G902), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n610), .A2(new_n606), .A3(new_n611), .A4(new_n612), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n547), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n605), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G472), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n353), .B2(new_n188), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n347), .A2(new_n349), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n621), .A2(new_n622), .A3(new_n243), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n448), .A2(new_n450), .A3(new_n619), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT103), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n624), .B(new_n626), .ZN(G6));
  NAND2_X1  g441(.A1(new_n442), .A2(new_n447), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n403), .A2(new_n430), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n370), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n430), .A2(KEYINPUT86), .A3(new_n371), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n445), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n188), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT87), .B1(new_n635), .B2(G469), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n450), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n527), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n540), .B2(new_n541), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n538), .B(new_n527), .C1(new_n528), .C2(new_n536), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n525), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n596), .A3(new_n599), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n605), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n638), .A2(new_n623), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  NOR2_X1   g461(.A1(new_n236), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n235), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n241), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n237), .A2(new_n238), .ZN(new_n652));
  OAI211_X1 g466(.A(KEYINPUT78), .B(new_n190), .C1(new_n652), .C2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n233), .A2(new_n188), .A3(new_n191), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n651), .B1(new_n655), .B2(new_n189), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n621), .A2(new_n622), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n448), .A2(new_n450), .A3(new_n601), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  INV_X1    g475(.A(new_n551), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(G900), .ZN(new_n663));
  INV_X1    g477(.A(new_n550), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n551), .A2(KEYINPUT104), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n596), .A2(new_n642), .A3(new_n599), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n240), .A2(new_n650), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n501), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n356), .B2(new_n366), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n448), .A3(new_n450), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  AOI21_X1  g488(.A(new_n250), .B1(new_n342), .B2(new_n317), .ZN(new_n675));
  AOI21_X1  g489(.A(G902), .B1(new_n357), .B2(new_n250), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n356), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n498), .A2(new_n500), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n499), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n547), .A2(new_n596), .A3(new_n599), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n681), .A2(new_n682), .A3(new_n670), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n667), .B(KEYINPUT39), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n638), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n679), .B(new_n684), .C1(new_n688), .C2(KEYINPUT40), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n269), .ZN(G45));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n354), .B1(new_n353), .B2(new_n348), .ZN(new_n694));
  AOI211_X1 g508(.A(KEYINPUT32), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n366), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n547), .A2(new_n614), .A3(new_n615), .A4(new_n668), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n656), .A2(new_n697), .A3(new_n604), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n693), .B1(new_n637), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n697), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n501), .A3(new_n670), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n356), .B2(new_n366), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n448), .A4(new_n450), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n430), .A2(new_n445), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n707), .A2(new_n370), .B1(new_n436), .B2(new_n403), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n450), .A3(new_n447), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n712), .A3(new_n447), .A4(new_n450), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n367), .A3(new_n619), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT108), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n367), .A2(new_n644), .A3(new_n713), .A4(new_n711), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NAND3_X1  g534(.A1(new_n670), .A2(new_n548), .A3(new_n600), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n356), .B2(new_n366), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n501), .A3(new_n713), .A4(new_n711), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n605), .A2(new_n683), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n360), .A2(new_n250), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n349), .B1(new_n352), .B2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n621), .A2(new_n243), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n725), .A2(new_n728), .A3(new_n713), .A4(new_n711), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  NOR4_X1   g544(.A1(new_n621), .A2(new_n656), .A3(new_n697), .A4(new_n727), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n501), .A3(new_n713), .A4(new_n711), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  INV_X1    g547(.A(new_n450), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n632), .A2(KEYINPUT109), .A3(new_n633), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n434), .B2(new_n437), .ZN(new_n737));
  OAI211_X1 g551(.A(G469), .B(new_n630), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n443), .A2(new_n188), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n447), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n734), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n680), .A2(new_n499), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n367), .A2(new_n742), .A3(new_n701), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n734), .B(new_n743), .C1(new_n738), .C2(new_n741), .ZN(new_n748));
  OR2_X1    g562(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n367), .A3(new_n701), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT111), .B(G131), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G33));
  AND4_X1   g567(.A1(new_n367), .A2(new_n742), .A3(new_n669), .A4(new_n744), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n254), .ZN(G36));
  OAI211_X1 g569(.A(KEYINPUT45), .B(new_n630), .C1(new_n735), .C2(new_n737), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n443), .B1(new_n634), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n739), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n447), .B1(new_n759), .B2(KEYINPUT46), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n450), .B(new_n685), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n617), .A2(new_n548), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT43), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n616), .A2(KEYINPUT43), .A3(new_n547), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n768), .B(new_n670), .C1(new_n622), .C2(new_n621), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n743), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n763), .B(new_n771), .C1(new_n770), .C2(new_n769), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  OAI21_X1  g587(.A(new_n450), .B1(new_n760), .B2(new_n761), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(KEYINPUT47), .B(new_n450), .C1(new_n760), .C2(new_n761), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n696), .ZN(new_n779));
  INV_X1    g593(.A(new_n243), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n697), .A3(new_n743), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(new_n681), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(new_n450), .A3(new_n499), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n785), .A3(new_n764), .ZN(new_n786));
  INV_X1    g600(.A(new_n679), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n709), .A2(new_n447), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n700), .A2(new_n704), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n670), .A2(new_n683), .A3(new_n604), .A4(new_n667), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n742), .A2(new_n679), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n673), .A2(new_n732), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n792), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n673), .A2(new_n732), .A3(new_n795), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n705), .A3(KEYINPUT52), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n754), .B1(new_n747), .B2(new_n750), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n715), .A2(new_n719), .A3(new_n723), .A4(new_n729), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n593), .A2(new_n598), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT112), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT112), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n548), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n605), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n448), .A2(new_n450), .A3(new_n623), .A4(new_n807), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n602), .A2(new_n624), .A3(new_n658), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n731), .A2(new_n742), .A3(new_n744), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n748), .A2(new_n812), .A3(new_n731), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n804), .A2(new_n805), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n642), .A2(new_n668), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n744), .A2(new_n670), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n779), .A2(new_n816), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n811), .A2(new_n813), .B1(new_n638), .B2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n801), .A2(new_n802), .A3(new_n809), .A4(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n798), .A2(new_n705), .A3(KEYINPUT52), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n800), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n798), .B2(new_n705), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n819), .B(KEYINPUT53), .C1(new_n820), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT54), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n714), .A2(new_n744), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n767), .A2(new_n664), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n367), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT48), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n831), .A2(new_n728), .ZN(new_n834));
  INV_X1    g648(.A(new_n714), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n604), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n549), .B(G953), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n679), .A2(new_n243), .A3(new_n664), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n830), .A2(KEYINPUT116), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n787), .A2(new_n780), .A3(new_n550), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n714), .A2(new_n744), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n833), .B(new_n837), .C1(new_n618), .C2(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n776), .B(new_n777), .C1(new_n450), .C2(new_n788), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n834), .A2(new_n744), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n621), .A2(new_n656), .A3(new_n727), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n830), .A2(new_n850), .A3(new_n831), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n617), .A2(new_n547), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n839), .A2(new_n843), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT115), .B1(new_n835), .B2(new_n499), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n714), .A2(new_n855), .A3(new_n682), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n831), .A2(new_n681), .A3(new_n728), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT50), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  AOI211_X1 g675(.A(new_n861), .B(new_n858), .C1(new_n854), .C2(new_n856), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n851), .B(new_n853), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT51), .B1(new_n849), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n853), .A2(new_n851), .ZN(new_n865));
  INV_X1    g679(.A(new_n860), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n857), .A2(KEYINPUT50), .A3(new_n859), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n848), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n845), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n800), .A2(new_n819), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n820), .A2(new_n826), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n715), .A2(new_n719), .A3(new_n723), .A4(new_n729), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n602), .A2(new_n624), .A3(new_n658), .A4(new_n808), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n801), .A3(new_n818), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n824), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n829), .A2(new_n871), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n882));
  INV_X1    g696(.A(G953), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n549), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n881), .A2(KEYINPUT117), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n791), .B1(new_n885), .B2(new_n886), .ZN(G75));
  NOR2_X1   g701(.A1(new_n227), .A2(G952), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT120), .Z(new_n889));
  AOI21_X1  g703(.A(new_n188), .B1(new_n872), .B2(new_n878), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(new_n496), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n487), .A2(new_n489), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n492), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n889), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(new_n188), .C1(new_n872), .C2(new_n878), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n898), .A2(new_n900), .A3(new_n497), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n872), .A2(new_n878), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G902), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n899), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n496), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT119), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n895), .B1(new_n903), .B2(new_n909), .ZN(G51));
  XNOR2_X1  g724(.A(new_n904), .B(new_n879), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n739), .B(KEYINPUT57), .Z(new_n912));
  OAI22_X1  g726(.A1(new_n911), .A2(new_n912), .B1(new_n446), .B2(new_n444), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n756), .A3(new_n758), .A4(new_n907), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n888), .B1(new_n913), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n907), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n540), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n540), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n888), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n879), .B1(new_n825), .B2(new_n827), .ZN(new_n924));
  INV_X1    g738(.A(new_n880), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n610), .A2(new_n611), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT121), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n610), .A2(new_n611), .A3(new_n923), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n889), .B1(new_n911), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(G63));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT60), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n872), .B2(new_n878), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n889), .B1(new_n936), .B2(new_n233), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n904), .A2(new_n649), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n933), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n904), .A2(new_n649), .A3(new_n938), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n943), .B(new_n889), .C1(new_n233), .C2(new_n936), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(KEYINPUT122), .A3(new_n933), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n944), .B2(new_n933), .ZN(new_n948));
  INV_X1    g762(.A(new_n937), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n943), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G66));
  AOI21_X1  g766(.A(new_n883), .B1(new_n553), .B2(G224), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT124), .ZN(new_n954));
  INV_X1    g768(.A(new_n227), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n876), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n892), .B1(G898), .B2(new_n227), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  AND2_X1   g772(.A1(new_n337), .A2(new_n341), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n533), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n705), .A2(new_n673), .A3(new_n732), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n689), .B2(new_n690), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n961), .C1(new_n689), .C2(new_n690), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n686), .B(KEYINPUT105), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n743), .B1(new_n618), .B2(new_n806), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n367), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n782), .A2(new_n968), .A3(new_n772), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n963), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n960), .B1(new_n970), .B2(new_n227), .ZN(new_n971));
  INV_X1    g785(.A(new_n683), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n367), .A2(new_n501), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n762), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT126), .Z(new_n975));
  AND3_X1   g789(.A1(new_n772), .A2(new_n801), .A3(new_n961), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n975), .A2(new_n976), .A3(new_n227), .A4(new_n782), .ZN(new_n977));
  INV_X1    g791(.A(new_n960), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(G900), .B2(new_n955), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n977), .B2(new_n979), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n971), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(G227), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n955), .B1(new_n985), .B2(new_n665), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n980), .A2(new_n987), .ZN(new_n988));
  OAI22_X1  g802(.A1(new_n984), .A2(new_n986), .B1(new_n971), .B2(new_n988), .ZN(G72));
  INV_X1    g803(.A(new_n675), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n963), .A2(new_n876), .A3(new_n965), .A4(new_n969), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  AOI21_X1  g807(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  AND4_X1   g808(.A1(new_n363), .A2(new_n828), .A3(new_n990), .A4(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n975), .A2(new_n976), .A3(new_n782), .A4(new_n876), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n363), .B1(new_n996), .B2(new_n993), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n994), .A2(new_n995), .A3(new_n888), .A4(new_n997), .ZN(G57));
endmodule


