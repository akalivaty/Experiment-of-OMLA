//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT64), .Z(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT65), .Z(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n462), .B2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n460), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G137), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n459), .B2(new_n472), .ZN(G160));
  AND2_X1   g048(.A1(new_n469), .A2(new_n463), .ZN(new_n474));
  AND4_X1   g049(.A1(KEYINPUT67), .A2(new_n474), .A3(new_n459), .A4(new_n468), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n468), .A2(new_n463), .A3(new_n469), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n476), .B2(new_n459), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n476), .A2(G124), .A3(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT68), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT69), .Z(G162));
  XOR2_X1   g061(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n461), .A2(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(new_n469), .A3(new_n490), .A4(new_n463), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n474), .A2(new_n496), .A3(new_n468), .A4(new_n490), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n468), .A2(new_n469), .A3(G126), .A4(new_n463), .ZN(new_n499));
  NAND2_X1  g074(.A1(G114), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n460), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G102), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n498), .A2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n514), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT72), .B(G88), .Z(new_n520));
  OAI22_X1  g095(.A1(new_n512), .A2(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n510), .A2(new_n521), .ZN(G166));
  XNOR2_X1  g097(.A(KEYINPUT73), .B(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n511), .A2(new_n523), .A3(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n507), .A2(new_n511), .A3(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n507), .A2(G63), .ZN(new_n530));
  NAND3_X1  g105(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n509), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G168));
  NAND3_X1  g108(.A1(new_n511), .A2(G52), .A3(G543), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OAI221_X1 g111(.A(new_n534), .B1(new_n535), .B2(new_n519), .C1(new_n536), .C2(new_n509), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(G43), .ZN(new_n539));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n512), .A2(new_n539), .B1(new_n519), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n507), .A2(G56), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n509), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(new_n519), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n509), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n554), .A3(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  NAND2_X1  g134(.A1(new_n553), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(G288));
  OAI21_X1  g138(.A(G61), .B1(new_n517), .B2(new_n518), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G73), .B2(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n507), .A2(KEYINPUT74), .A3(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n509), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G48), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n512), .A2(new_n569), .B1(new_n519), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n509), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n512), .A2(new_n576), .B1(new_n519), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G54), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n582), .A2(new_n509), .B1(new_n583), .B2(new_n512), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI221_X1 g161(.A(KEYINPUT76), .B1(new_n512), .B2(new_n583), .C1(new_n582), .C2(new_n509), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n553), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n581), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n581), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  XOR2_X1   g173(.A(G280), .B(KEYINPUT77), .Z(G297));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n476), .A2(G2105), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G123), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n610));
  INV_X1    g185(.A(G135), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n610), .C1(new_n478), .C2(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(G2096), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(G2427), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G14), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n631), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT79), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n635), .A2(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT80), .ZN(new_n641));
  NOR2_X1   g216(.A1(G2072), .A2(G2078), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n442), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n639), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n643), .B(KEYINPUT17), .Z(new_n646));
  OAI21_X1  g221(.A(new_n645), .B1(new_n646), .B2(new_n641), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n643), .A2(new_n639), .A3(new_n640), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT18), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n641), .A3(new_n639), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(G227));
  XNOR2_X1  g228(.A(G1971), .B(G1976), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT81), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n664), .C1(new_n655), .C2(new_n663), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1981), .B(G1986), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT84), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n671), .B1(new_n669), .B2(new_n672), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n677), .B1(new_n674), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(G29), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G32), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n476), .A2(G129), .A3(G2105), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT26), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n690), .A2(new_n691), .B1(G105), .B2(new_n503), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n479), .A2(G141), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT92), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n684), .B1(new_n696), .B2(new_n683), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT27), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G6), .A2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n572), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G23), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT85), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G288), .B2(new_n704), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT33), .B(G1976), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n708), .A2(new_n712), .A3(new_n713), .A4(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n704), .A2(G24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n579), .B2(new_n704), .ZN(new_n722));
  INV_X1    g297(.A(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G25), .A2(G29), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n727));
  INV_X1    g302(.A(G119), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n606), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n479), .B2(G131), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT35), .B(G1991), .Z(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n724), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n731), .B2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n720), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(KEYINPUT86), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n737), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n683), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n683), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT29), .B(G2090), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n704), .A2(G20), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT23), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n597), .B2(new_n704), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n704), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n704), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1961), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n704), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n545), .B2(new_n704), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1341), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n704), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n704), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1966), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n683), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n683), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n748), .B(new_n758), .C1(G2078), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n683), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  OR2_X1    g338(.A1(G104), .A2(G2105), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n764), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n765));
  INV_X1    g340(.A(G128), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n606), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n479), .B2(G140), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(new_n683), .ZN(new_n769));
  INV_X1    g344(.A(G2067), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G160), .B2(new_n683), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  OAI221_X1 g353(.A(new_n771), .B1(G2078), .B2(new_n760), .C1(new_n772), .C2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n761), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n772), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  INV_X1    g358(.A(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(KEYINPUT30), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n784), .B2(KEYINPUT30), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n612), .A2(new_n683), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n744), .A2(new_n781), .A3(new_n783), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n683), .A2(G33), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT25), .Z(new_n798));
  INV_X1    g373(.A(G139), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n478), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT88), .Z(new_n801));
  NAND2_X1  g376(.A1(G115), .A2(G2104), .ZN(new_n802));
  INV_X1    g377(.A(G127), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n488), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n459), .B1(new_n804), .B2(KEYINPUT89), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT89), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n796), .B1(new_n808), .B2(new_n683), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(G2072), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n704), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n593), .B2(new_n704), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT87), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1348), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(G2072), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n698), .B2(new_n700), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n703), .A2(new_n740), .A3(new_n795), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  AND2_X1   g394(.A1(new_n507), .A2(G67), .ZN(new_n820));
  AND2_X1   g395(.A1(G80), .A2(G543), .ZN(new_n821));
  OAI21_X1  g396(.A(G651), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT98), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n514), .A2(new_n516), .A3(G55), .A4(G543), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n823), .B(new_n824), .C1(new_n519), .C2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n507), .A2(new_n511), .A3(G93), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(new_n824), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n822), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n541), .A2(new_n544), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n545), .B(new_n822), .C1(new_n829), .C2(new_n827), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT38), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n593), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n830), .A2(G860), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n612), .B(G160), .ZN(new_n844));
  XNOR2_X1  g419(.A(G162), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n696), .A2(new_n808), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n807), .A2(new_n695), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n501), .A2(G2105), .B1(G102), .B2(new_n503), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n498), .B2(KEYINPUT99), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT99), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n850), .B(new_n492), .C1(new_n497), .C2(new_n495), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n846), .A2(new_n847), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n857));
  INV_X1    g432(.A(G106), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n459), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n859), .B1(new_n607), .B2(G130), .ZN(new_n860));
  INV_X1    g435(.A(G142), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n478), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n616), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n730), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n730), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n768), .ZN(new_n867));
  INV_X1    g442(.A(new_n768), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n864), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n854), .B1(new_n846), .B2(new_n847), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n856), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n854), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n695), .B(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(new_n807), .ZN(new_n876));
  INV_X1    g451(.A(new_n847), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n878), .A2(new_n855), .B1(new_n867), .B2(new_n869), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n845), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n870), .B1(new_n856), .B2(new_n871), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n878), .A2(new_n867), .A3(new_n869), .A4(new_n855), .ZN(new_n883));
  INV_X1    g458(.A(new_n845), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g462(.A(new_n602), .B(new_n834), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n592), .A2(new_n597), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n588), .A2(G299), .A3(new_n591), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  INV_X1    g468(.A(new_n890), .ZN(new_n894));
  AOI21_X1  g469(.A(G299), .B1(new_n588), .B2(new_n591), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n892), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(KEYINPUT42), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G288), .B(KEYINPUT101), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n572), .ZN(new_n905));
  XNOR2_X1  g480(.A(G166), .B(new_n579), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n903), .B(new_n908), .ZN(new_n909));
  MUX2_X1   g484(.A(new_n830), .B(new_n909), .S(G868), .Z(G295));
  MUX2_X1   g485(.A(new_n830), .B(new_n909), .S(G868), .Z(G331));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT102), .B1(new_n529), .B2(new_n532), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G301), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n912), .A3(G301), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n834), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n913), .A2(new_n912), .A3(G301), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n832), .B(new_n833), .C1(new_n918), .C2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g496(.A1(G168), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n917), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n898), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT104), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n923), .A2(new_n898), .A3(new_n928), .A4(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(new_n925), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n924), .B1(new_n917), .B2(new_n919), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n891), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n908), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n927), .A2(new_n907), .A3(new_n929), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n881), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n923), .A2(new_n898), .A3(new_n940), .A4(new_n925), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n932), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n908), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n936), .A2(new_n881), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n946), .A3(new_n908), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n948), .B2(KEYINPUT43), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n946), .B1(new_n942), .B2(new_n908), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n953), .A2(new_n937), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n952), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n934), .A2(new_n952), .A3(new_n881), .A4(new_n936), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n957), .A2(KEYINPUT44), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT107), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n951), .B1(new_n959), .B2(new_n962), .ZN(G397));
  INV_X1    g538(.A(KEYINPUT127), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT112), .B(G8), .ZN(new_n965));
  NOR2_X1   g540(.A1(G168), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(G8), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n849), .B2(new_n851), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n472), .A2(new_n459), .ZN(new_n973));
  INV_X1    g548(.A(new_n466), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(G40), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n969), .B(new_n981), .C1(new_n498), .C2(new_n505), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G1966), .B1(new_n972), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n969), .B1(new_n498), .B2(new_n505), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n985), .A2(KEYINPUT50), .B1(new_n977), .B2(new_n978), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(new_n969), .C1(new_n849), .C2(new_n851), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n986), .A2(new_n988), .A3(new_n772), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n968), .B1(new_n984), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n988), .A3(new_n772), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n979), .A2(new_n982), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n971), .B2(new_n970), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n991), .B(new_n967), .C1(new_n993), .C2(G1966), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(KEYINPUT51), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT62), .ZN(new_n996));
  INV_X1    g571(.A(new_n965), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n984), .B2(new_n989), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n966), .A2(KEYINPUT51), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n995), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n986), .A2(new_n988), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n986), .A2(new_n988), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT126), .B(G1961), .Z(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n985), .A2(new_n980), .B1(new_n977), .B2(new_n978), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT45), .B(new_n969), .C1(new_n849), .C2(new_n851), .ZN(new_n1012));
  INV_X1    g587(.A(G2078), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1008), .A2(new_n1009), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n1013), .ZN(new_n1016));
  AOI21_X1  g591(.A(G301), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n1018));
  OAI211_X1 g593(.A(KEYINPUT55), .B(G8), .C1(new_n510), .C2(new_n521), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT110), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1019), .A2(KEYINPUT110), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(KEYINPUT110), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(KEYINPUT111), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  NOR2_X1   g601(.A1(G166), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1027), .A2(KEYINPUT55), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1971), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n987), .B(new_n969), .C1(new_n498), .C2(new_n505), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n979), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(KEYINPUT50), .B2(new_n970), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1018), .B(new_n1030), .C1(new_n1036), .C2(new_n965), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1031), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1034), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n1032), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n965), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT117), .B1(new_n1042), .B2(new_n1029), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n560), .A2(G1976), .A3(new_n561), .A4(new_n562), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n977), .A2(new_n978), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n997), .B(new_n1044), .C1(new_n970), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n979), .B(new_n969), .C1(new_n851), .C2(new_n849), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n564), .A2(new_n565), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G73), .A2(G543), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n567), .ZN(new_n1052));
  OAI21_X1  g627(.A(G651), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  INV_X1    g629(.A(new_n571), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(G1981), .B1(new_n568), .B2(new_n571), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT49), .B1(new_n1059), .B2(KEYINPUT115), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT114), .B1(KEYINPUT115), .B2(KEYINPUT49), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n997), .B(new_n1048), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT113), .B(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1048), .A2(new_n997), .A3(new_n1044), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1047), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n986), .A2(new_n988), .A3(new_n1032), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1026), .B1(new_n1038), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1029), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1017), .A2(new_n1037), .A3(new_n1043), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n964), .B1(new_n1003), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1014), .A2(new_n1010), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1016), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n995), .A2(new_n1000), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1082), .A3(KEYINPUT127), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1072), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1348), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n986), .A2(new_n988), .A3(new_n1006), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1006), .B1(new_n986), .B2(new_n988), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1048), .A2(G2067), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n593), .A2(KEYINPUT125), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n592), .B(KEYINPUT125), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1089), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1092), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(G299), .B(KEYINPUT57), .Z(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT121), .B(G1956), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1011), .A2(new_n1012), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1100), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1099), .B(new_n1105), .C1(new_n1035), .C2(new_n1102), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(KEYINPUT61), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT61), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n831), .B1(new_n1112), .B2(KEYINPUT59), .ZN(new_n1113));
  INV_X1    g688(.A(G1996), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1011), .A2(new_n1012), .A3(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n970), .B2(new_n1045), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT123), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT123), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1113), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1121), .B(new_n1113), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1098), .A2(new_n1111), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1107), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1108), .A2(new_n593), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(new_n1095), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G301), .B(KEYINPUT54), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1076), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1012), .ZN(new_n1133));
  NOR4_X1   g708(.A1(new_n1133), .A2(new_n1010), .A3(G2078), .A4(new_n975), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n970), .A2(new_n980), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1015), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1132), .A2(new_n995), .A3(new_n1000), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n1073), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1130), .A2(new_n1139), .ZN(new_n1140));
  NOR4_X1   g715(.A1(new_n1060), .A2(G1976), .A3(G288), .A4(new_n1062), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1056), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n997), .B(new_n1048), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1068), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1029), .B(G8), .C1(new_n1144), .C2(new_n1031), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1145), .B2(new_n1067), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(KEYINPUT63), .ZN(new_n1148));
  OAI211_X1 g723(.A(G168), .B(new_n997), .C1(new_n984), .C2(new_n989), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(KEYINPUT118), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(new_n1144), .B2(new_n1031), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1067), .B1(new_n1030), .B2(new_n1153), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1152), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1158));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1149), .B(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1158), .B1(new_n1073), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1147), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1084), .A2(new_n1140), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1135), .A2(new_n1045), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n696), .A2(new_n1114), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n695), .A2(G1996), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n768), .B(G2067), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n730), .A2(new_n732), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n730), .A2(new_n732), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1165), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n579), .B(new_n723), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1164), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1175), .A2(new_n1169), .B1(G2067), .B2(new_n868), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1164), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT47), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1167), .A2(new_n694), .A3(new_n693), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1164), .A2(new_n1114), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT46), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1164), .A2(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1181), .B2(new_n1180), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1171), .A2(new_n1164), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1164), .A2(new_n723), .A3(new_n579), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT48), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1189));
  OAI221_X1 g764(.A(new_n1177), .B1(new_n1178), .B2(new_n1183), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1190), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1174), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(G319), .ZN(new_n1194));
  NOR2_X1   g768(.A1(G227), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1195), .B1(new_n635), .B2(new_n637), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n679), .B2(new_n680), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n1197), .A2(new_n886), .A3(new_n949), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


