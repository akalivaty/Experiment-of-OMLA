

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G164), .A2(G1384), .ZN(n782) );
  OR2_X1 U551 ( .A1(n779), .A2(n778), .ZN(n517) );
  XOR2_X2 U552 ( .A(KEYINPUT17), .B(n520), .Z(n990) );
  NAND2_X1 U553 ( .A1(n780), .A2(n782), .ZN(n736) );
  NAND2_X1 U554 ( .A1(n736), .A2(G8), .ZN(n724) );
  NOR2_X1 U555 ( .A1(n814), .A2(n813), .ZN(n518) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n732) );
  NOR2_X1 U557 ( .A1(n759), .A2(G1966), .ZN(n749) );
  INV_X1 U558 ( .A(n939), .ZN(n758) );
  XNOR2_X1 U559 ( .A(n754), .B(KEYINPUT105), .ZN(n775) );
  AND2_X1 U560 ( .A1(n761), .A2(n760), .ZN(n765) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(n724), .Z(n777) );
  NOR2_X2 U562 ( .A1(G2105), .A2(n523), .ZN(n989) );
  NOR2_X1 U563 ( .A1(G651), .A2(n642), .ZN(n648) );
  AND2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n985) );
  NAND2_X1 U565 ( .A1(G114), .A2(n985), .ZN(n519) );
  XNOR2_X1 U566 ( .A(n519), .B(KEYINPUT94), .ZN(n522) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n990), .A2(G138), .ZN(n521) );
  NAND2_X1 U569 ( .A1(n522), .A2(n521), .ZN(n527) );
  INV_X1 U570 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U571 ( .A1(G102), .A2(n989), .ZN(n525) );
  AND2_X1 U572 ( .A1(n523), .A2(G2105), .ZN(n986) );
  NAND2_X1 U573 ( .A1(G126), .A2(n986), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U575 ( .A1(n527), .A2(n526), .ZN(G164) );
  XOR2_X1 U576 ( .A(G2427), .B(G2446), .Z(n529) );
  XNOR2_X1 U577 ( .A(G1341), .B(G2430), .ZN(n528) );
  XNOR2_X1 U578 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U579 ( .A(n530), .B(G2435), .Z(n532) );
  XNOR2_X1 U580 ( .A(G1348), .B(G2438), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n532), .B(n531), .ZN(n536) );
  XOR2_X1 U582 ( .A(G2454), .B(G2451), .Z(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(G2443), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U585 ( .A(n536), .B(n535), .Z(n537) );
  AND2_X1 U586 ( .A1(G14), .A2(n537), .ZN(G401) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NAND2_X1 U588 ( .A1(n648), .A2(G52), .ZN(n541) );
  XNOR2_X1 U589 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n539) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(G651), .ZN(n542) );
  NOR2_X1 U591 ( .A1(G543), .A2(n542), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n539), .B(n538), .ZN(n650) );
  NAND2_X1 U593 ( .A1(G64), .A2(n650), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n548) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U596 ( .A1(G90), .A2(n649), .ZN(n545) );
  NOR2_X1 U597 ( .A1(n642), .A2(n542), .ZN(n543) );
  XNOR2_X1 U598 ( .A(KEYINPUT66), .B(n543), .ZN(n653) );
  NAND2_X1 U599 ( .A1(G77), .A2(n653), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U602 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U604 ( .A1(G111), .A2(n985), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G99), .A2(n989), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G135), .A2(n990), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n986), .A2(G123), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT18), .B(n551), .Z(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT78), .ZN(n996) );
  XNOR2_X1 U613 ( .A(n996), .B(G2096), .ZN(n557) );
  OR2_X1 U614 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  NAND2_X1 U617 ( .A1(G50), .A2(n648), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT84), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n650), .A2(G62), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT83), .B(n559), .Z(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G88), .A2(n649), .ZN(n562) );
  XNOR2_X1 U623 ( .A(KEYINPUT85), .B(n562), .ZN(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n653), .A2(G75), .ZN(n565) );
  NAND2_X1 U626 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT86), .B(n567), .Z(G166) );
  INV_X1 U628 ( .A(G166), .ZN(G303) );
  NAND2_X1 U629 ( .A1(G101), .A2(n989), .ZN(n568) );
  XOR2_X1 U630 ( .A(KEYINPUT64), .B(n568), .Z(n569) );
  XNOR2_X1 U631 ( .A(n569), .B(KEYINPUT23), .ZN(n695) );
  NAND2_X1 U632 ( .A1(G137), .A2(n990), .ZN(n693) );
  NAND2_X1 U633 ( .A1(n695), .A2(n693), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G113), .A2(n985), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G125), .A2(n986), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n691) );
  NOR2_X1 U637 ( .A1(n572), .A2(n691), .ZN(G160) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U640 ( .A(G223), .B(KEYINPUT71), .ZN(n830) );
  NAND2_X1 U641 ( .A1(n830), .A2(G567), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n576) );
  NAND2_X1 U644 ( .A1(G56), .A2(n650), .ZN(n575) );
  XNOR2_X1 U645 ( .A(n576), .B(n575), .ZN(n584) );
  XOR2_X1 U646 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n578) );
  NAND2_X1 U647 ( .A1(G81), .A2(n649), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U649 ( .A(KEYINPUT73), .B(n579), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n653), .A2(G68), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n648), .A2(G43), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n963) );
  INV_X1 U656 ( .A(G860), .ZN(n619) );
  OR2_X1 U657 ( .A1(n963), .A2(n619), .ZN(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G92), .A2(n649), .ZN(n594) );
  NAND2_X1 U661 ( .A1(G79), .A2(n653), .ZN(n588) );
  NAND2_X1 U662 ( .A1(G54), .A2(n648), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U664 ( .A(KEYINPUT76), .B(n589), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G66), .A2(n650), .ZN(n590) );
  XNOR2_X1 U666 ( .A(KEYINPUT75), .B(n590), .ZN(n591) );
  NOR2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n595) );
  XNOR2_X1 U670 ( .A(n596), .B(n595), .ZN(n962) );
  OR2_X1 U671 ( .A1(n962), .A2(G868), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U673 ( .A1(n649), .A2(G89), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n599), .B(KEYINPUT4), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G76), .A2(n653), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT5), .ZN(n607) );
  NAND2_X1 U678 ( .A1(n648), .A2(G51), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G63), .A2(n650), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT6), .B(n605), .Z(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U684 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U685 ( .A1(n648), .A2(G53), .ZN(n610) );
  NAND2_X1 U686 ( .A1(G65), .A2(n650), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U688 ( .A(KEYINPUT69), .B(n611), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G91), .A2(n649), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G78), .A2(n653), .ZN(n612) );
  AND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(G299) );
  INV_X1 U693 ( .A(G868), .ZN(n616) );
  NOR2_X1 U694 ( .A1(G286), .A2(n616), .ZN(n618) );
  NOR2_X1 U695 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U696 ( .A1(n618), .A2(n617), .ZN(G297) );
  NAND2_X1 U697 ( .A1(n619), .A2(G559), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n620), .A2(n962), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n621), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U700 ( .A1(G868), .A2(n963), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G868), .A2(n962), .ZN(n622) );
  NOR2_X1 U702 ( .A1(G559), .A2(n622), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(G282) );
  NAND2_X1 U704 ( .A1(G559), .A2(n962), .ZN(n625) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(n625), .Z(n626) );
  XNOR2_X1 U706 ( .A(n963), .B(n626), .ZN(n668) );
  NOR2_X1 U707 ( .A1(n668), .A2(G860), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G93), .A2(n649), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n627), .B(KEYINPUT80), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G67), .A2(n650), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G80), .A2(n653), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G55), .A2(n648), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n671) );
  XNOR2_X1 U716 ( .A(n634), .B(n671), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G85), .A2(n649), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G72), .A2(n653), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n650), .A2(G60), .ZN(n637) );
  XOR2_X1 U721 ( .A(KEYINPUT68), .B(n637), .Z(n638) );
  NOR2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n648), .A2(G47), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U725 ( .A1(G87), .A2(n642), .ZN(n644) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U728 ( .A1(n650), .A2(n645), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(G49), .ZN(n646) );
  NAND2_X1 U730 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U731 ( .A1(n648), .A2(G48), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n649), .A2(G86), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n657) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n655) );
  NAND2_X1 U736 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U737 ( .A(n655), .B(n654), .Z(n656) );
  NOR2_X1 U738 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n660), .B(KEYINPUT82), .ZN(G305) );
  XNOR2_X1 U741 ( .A(G303), .B(n671), .ZN(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n662) );
  XNOR2_X1 U743 ( .A(G288), .B(KEYINPUT19), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U746 ( .A(G290), .B(n665), .ZN(n667) );
  INV_X1 U747 ( .A(G299), .ZN(n703) );
  XNOR2_X1 U748 ( .A(G305), .B(n703), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n959) );
  XNOR2_X1 U750 ( .A(n959), .B(n668), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n669), .A2(G868), .ZN(n670) );
  XOR2_X1 U752 ( .A(KEYINPUT89), .B(n670), .Z(n673) );
  OR2_X1 U753 ( .A1(n671), .A2(G868), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U758 ( .A(n676), .B(KEYINPUT91), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n677) );
  XNOR2_X1 U760 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U763 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT22), .B(KEYINPUT92), .ZN(n680) );
  XNOR2_X1 U766 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n682), .A2(G96), .ZN(n683) );
  NOR2_X1 U768 ( .A1(G218), .A2(n683), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT93), .B(n684), .ZN(n834) );
  NAND2_X1 U770 ( .A1(n834), .A2(G2106), .ZN(n688) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U772 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U773 ( .A1(G108), .A2(n686), .ZN(n835) );
  NAND2_X1 U774 ( .A1(n835), .A2(G567), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n1018) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n1018), .A2(n689), .ZN(n833) );
  NAND2_X1 U778 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G40), .ZN(n690) );
  NOR2_X1 U780 ( .A1(n691), .A2(n690), .ZN(n692) );
  AND2_X1 U781 ( .A1(n693), .A2(n692), .ZN(n694) );
  AND2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n780) );
  INV_X1 U783 ( .A(G1961), .ZN(n869) );
  NAND2_X1 U784 ( .A1(n736), .A2(n869), .ZN(n697) );
  INV_X1 U785 ( .A(n736), .ZN(n710) );
  XNOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .ZN(n850) );
  NAND2_X1 U787 ( .A1(n710), .A2(n850), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n729) );
  NAND2_X1 U789 ( .A1(n729), .A2(G171), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G2072), .A2(n710), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT27), .ZN(n699) );
  XNOR2_X1 U792 ( .A(KEYINPUT102), .B(n699), .ZN(n701) );
  AND2_X1 U793 ( .A1(n736), .A2(G1956), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n702) );
  XOR2_X1 U796 ( .A(n702), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n718) );
  INV_X1 U798 ( .A(G1996), .ZN(n848) );
  NOR2_X1 U799 ( .A1(n736), .A2(n848), .ZN(n705) );
  XOR2_X1 U800 ( .A(n705), .B(KEYINPUT26), .Z(n707) );
  NAND2_X1 U801 ( .A1(n736), .A2(G1341), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n963), .A2(n708), .ZN(n709) );
  OR2_X1 U804 ( .A1(n962), .A2(n709), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n962), .A2(n709), .ZN(n714) );
  NAND2_X1 U806 ( .A1(G1348), .A2(n736), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n710), .A2(G2067), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U813 ( .A(KEYINPUT29), .B(n721), .Z(n722) );
  NAND2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n735) );
  XNOR2_X1 U815 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n727) );
  INV_X1 U816 ( .A(n777), .ZN(n759) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n736), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n749), .A2(n745), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n725), .A2(G8), .ZN(n726) );
  XOR2_X1 U820 ( .A(n727), .B(n726), .Z(n728) );
  NOR2_X1 U821 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U822 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n733) );
  XNOR2_X1 U824 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n747) );
  NAND2_X1 U826 ( .A1(G286), .A2(n747), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n736), .ZN(n737) );
  XNOR2_X1 U828 ( .A(n737), .B(KEYINPUT104), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n759), .A2(G1971), .ZN(n738) );
  NOR2_X1 U830 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U831 ( .A1(G303), .A2(n740), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(n743), .A2(G8), .ZN(n744) );
  XNOR2_X1 U834 ( .A(n744), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U835 ( .A1(G8), .A2(n745), .ZN(n746) );
  XOR2_X1 U836 ( .A(KEYINPUT101), .B(n746), .Z(n751) );
  INV_X1 U837 ( .A(n747), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  INV_X1 U841 ( .A(n775), .ZN(n757) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n938) );
  NOR2_X1 U843 ( .A1(G303), .A2(G1971), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n938), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n761) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NOR2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT24), .ZN(n763) );
  AND2_X1 U850 ( .A1(n763), .A2(n777), .ZN(n766) );
  OR2_X1 U851 ( .A1(KEYINPUT33), .A2(n766), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n772) );
  INV_X1 U853 ( .A(n766), .ZN(n770) );
  AND2_X1 U854 ( .A1(n938), .A2(KEYINPUT33), .ZN(n767) );
  AND2_X1 U855 ( .A1(n767), .A2(n777), .ZN(n768) );
  XNOR2_X1 U856 ( .A(G1981), .B(G305), .ZN(n948) );
  OR2_X1 U857 ( .A1(n768), .A2(n948), .ZN(n769) );
  AND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n779) );
  NAND2_X1 U860 ( .A1(G8), .A2(G166), .ZN(n773) );
  NOR2_X1 U861 ( .A1(G2090), .A2(n773), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U864 ( .A(G1986), .B(G290), .ZN(n946) );
  INV_X1 U865 ( .A(n780), .ZN(n781) );
  NOR2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n825) );
  AND2_X1 U867 ( .A1(n946), .A2(n825), .ZN(n814) );
  NAND2_X1 U868 ( .A1(G104), .A2(n989), .ZN(n784) );
  NAND2_X1 U869 ( .A1(G140), .A2(n990), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n785), .ZN(n791) );
  NAND2_X1 U872 ( .A1(n985), .A2(G116), .ZN(n786) );
  XOR2_X1 U873 ( .A(KEYINPUT95), .B(n786), .Z(n788) );
  NAND2_X1 U874 ( .A1(n986), .A2(G128), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U876 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n792), .ZN(n1002) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  NOR2_X1 U880 ( .A1(n1002), .A2(n823), .ZN(n903) );
  NAND2_X1 U881 ( .A1(n903), .A2(n825), .ZN(n821) );
  NAND2_X1 U882 ( .A1(G107), .A2(n985), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G119), .A2(n986), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U885 ( .A(KEYINPUT96), .B(n795), .Z(n799) );
  NAND2_X1 U886 ( .A1(n989), .A2(G95), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G131), .A2(n990), .ZN(n796) );
  AND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n998) );
  NAND2_X1 U890 ( .A1(G1991), .A2(n998), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT97), .B(n800), .Z(n810) );
  XOR2_X1 U892 ( .A(KEYINPUT98), .B(KEYINPUT38), .Z(n802) );
  NAND2_X1 U893 ( .A1(G105), .A2(n989), .ZN(n801) );
  XNOR2_X1 U894 ( .A(n802), .B(n801), .ZN(n806) );
  NAND2_X1 U895 ( .A1(G141), .A2(n990), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G117), .A2(n985), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n986), .A2(G129), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n1008) );
  NAND2_X1 U901 ( .A1(G1996), .A2(n1008), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n902) );
  NAND2_X1 U903 ( .A1(n902), .A2(n825), .ZN(n811) );
  XOR2_X1 U904 ( .A(KEYINPUT99), .B(n811), .Z(n812) );
  NAND2_X1 U905 ( .A1(n821), .A2(n812), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n517), .A2(n518), .ZN(n828) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n1008), .ZN(n907) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n998), .ZN(n899) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n815) );
  XNOR2_X1 U910 ( .A(KEYINPUT106), .B(n815), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n899), .A2(n816), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT107), .B(n817), .Z(n818) );
  NOR2_X1 U913 ( .A1(n902), .A2(n818), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n907), .A2(n819), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n1002), .A2(n823), .ZN(n904) );
  NAND2_X1 U918 ( .A1(n824), .A2(n904), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT40), .B(n829), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  NOR2_X1 U927 ( .A1(n835), .A2(n834), .ZN(G325) );
  XNOR2_X1 U928 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  NAND2_X1 U930 ( .A1(G124), .A2(n986), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n836), .B(KEYINPUT44), .ZN(n839) );
  NAND2_X1 U932 ( .A1(G136), .A2(n990), .ZN(n837) );
  XOR2_X1 U933 ( .A(KEYINPUT111), .B(n837), .Z(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(n845) );
  NAND2_X1 U935 ( .A1(n989), .A2(G100), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n840), .B(KEYINPUT112), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G112), .A2(n985), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(KEYINPUT113), .B(n843), .Z(n844) );
  NOR2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G162) );
  INV_X1 U941 ( .A(KEYINPUT55), .ZN(n929) );
  XNOR2_X1 U942 ( .A(G2090), .B(G35), .ZN(n861) );
  XNOR2_X1 U943 ( .A(G2067), .B(G26), .ZN(n847) );
  XNOR2_X1 U944 ( .A(G1991), .B(G25), .ZN(n846) );
  NOR2_X1 U945 ( .A1(n847), .A2(n846), .ZN(n855) );
  XNOR2_X1 U946 ( .A(G32), .B(n848), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n849), .A2(G28), .ZN(n853) );
  XOR2_X1 U948 ( .A(G27), .B(n850), .Z(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT120), .B(n851), .ZN(n852) );
  NOR2_X1 U950 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U951 ( .A1(n855), .A2(n854), .ZN(n858) );
  XOR2_X1 U952 ( .A(KEYINPUT119), .B(G2072), .Z(n856) );
  XNOR2_X1 U953 ( .A(G33), .B(n856), .ZN(n857) );
  NOR2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U955 ( .A(KEYINPUT53), .B(n859), .ZN(n860) );
  NOR2_X1 U956 ( .A1(n861), .A2(n860), .ZN(n864) );
  XOR2_X1 U957 ( .A(G2084), .B(G34), .Z(n862) );
  XNOR2_X1 U958 ( .A(KEYINPUT54), .B(n862), .ZN(n863) );
  NAND2_X1 U959 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U960 ( .A(n929), .B(n865), .ZN(n867) );
  INV_X1 U961 ( .A(G29), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G11), .A2(n868), .ZN(n897) );
  XNOR2_X1 U964 ( .A(G5), .B(n869), .ZN(n890) );
  XOR2_X1 U965 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n876) );
  XNOR2_X1 U966 ( .A(G1976), .B(G23), .ZN(n871) );
  XNOR2_X1 U967 ( .A(G1986), .B(G24), .ZN(n870) );
  NOR2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n874) );
  XOR2_X1 U969 ( .A(G1971), .B(KEYINPUT124), .Z(n872) );
  XNOR2_X1 U970 ( .A(G22), .B(n872), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n876), .B(n875), .ZN(n888) );
  XNOR2_X1 U973 ( .A(G1956), .B(KEYINPUT122), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n877), .B(G20), .ZN(n882) );
  XNOR2_X1 U975 ( .A(G1981), .B(G6), .ZN(n879) );
  XNOR2_X1 U976 ( .A(G19), .B(G1341), .ZN(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n880), .B(KEYINPUT123), .ZN(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n885) );
  XNOR2_X1 U980 ( .A(G1348), .B(KEYINPUT59), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(G4), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT60), .B(n886), .ZN(n887) );
  NOR2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n892) );
  XNOR2_X1 U986 ( .A(G21), .B(G1966), .ZN(n891) );
  NOR2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U988 ( .A(KEYINPUT61), .B(n893), .Z(n894) );
  NOR2_X1 U989 ( .A1(G16), .A2(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n895), .B(KEYINPUT126), .ZN(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n933) );
  XOR2_X1 U992 ( .A(G2084), .B(G160), .Z(n898) );
  NOR2_X1 U993 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U994 ( .A1(n996), .A2(n900), .ZN(n901) );
  NOR2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n914) );
  INV_X1 U996 ( .A(n903), .ZN(n905) );
  NAND2_X1 U997 ( .A1(n905), .A2(n904), .ZN(n912) );
  XOR2_X1 U998 ( .A(G2090), .B(G162), .Z(n906) );
  NOR2_X1 U999 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1000 ( .A(KEYINPUT51), .B(n908), .Z(n910) );
  XNOR2_X1 U1001 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1003 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1004 ( .A1(n914), .A2(n913), .ZN(n927) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n989), .ZN(n916) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n990), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1008 ( .A(KEYINPUT114), .B(n917), .ZN(n922) );
  NAND2_X1 U1009 ( .A1(G115), .A2(n985), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(G127), .A2(n986), .ZN(n918) );
  NAND2_X1 U1011 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1013 ( .A1(n922), .A2(n921), .ZN(n1001) );
  XOR2_X1 U1014 ( .A(G2072), .B(n1001), .Z(n924) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1016 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1017 ( .A(KEYINPUT50), .B(n925), .Z(n926) );
  NOR2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(KEYINPUT52), .B(n928), .ZN(n930) );
  NAND2_X1 U1020 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1021 ( .A1(n931), .A2(G29), .ZN(n932) );
  NAND2_X1 U1022 ( .A1(n933), .A2(n932), .ZN(n957) );
  XOR2_X1 U1023 ( .A(G16), .B(KEYINPUT56), .Z(n955) );
  XNOR2_X1 U1024 ( .A(G1348), .B(n962), .ZN(n937) );
  XNOR2_X1 U1025 ( .A(G301), .B(G1961), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(n963), .B(G1341), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n937), .A2(n936), .ZN(n953) );
  XNOR2_X1 U1029 ( .A(G1971), .B(G166), .ZN(n944) );
  XNOR2_X1 U1030 ( .A(KEYINPUT121), .B(n938), .ZN(n940) );
  NAND2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n942) );
  XNOR2_X1 U1032 ( .A(G1956), .B(G299), .ZN(n941) );
  NOR2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n951) );
  XOR2_X1 U1036 ( .A(G168), .B(G1966), .Z(n947) );
  NOR2_X1 U1037 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1038 ( .A(KEYINPUT57), .B(n949), .Z(n950) );
  NAND2_X1 U1039 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1040 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1041 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1042 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1043 ( .A(n958), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1044 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1045 ( .A(G120), .ZN(G236) );
  INV_X1 U1046 ( .A(G96), .ZN(G221) );
  INV_X1 U1047 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1048 ( .A(KEYINPUT115), .B(n959), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G171), .B(G286), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1051 ( .A(n963), .B(n962), .Z(n964) );
  XNOR2_X1 U1052 ( .A(n965), .B(n964), .ZN(n966) );
  NOR2_X1 U1053 ( .A1(G37), .A2(n966), .ZN(G397) );
  XNOR2_X1 U1054 ( .A(G1976), .B(KEYINPUT110), .ZN(n976) );
  XOR2_X1 U1055 ( .A(G1986), .B(G1956), .Z(n968) );
  XNOR2_X1 U1056 ( .A(G1981), .B(G1966), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(n968), .B(n967), .ZN(n972) );
  XOR2_X1 U1058 ( .A(G2474), .B(KEYINPUT41), .Z(n970) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G1991), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1061 ( .A(n972), .B(n971), .Z(n974) );
  XNOR2_X1 U1062 ( .A(G1961), .B(G1971), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(G229) );
  XOR2_X1 U1065 ( .A(G2100), .B(G2096), .Z(n978) );
  XNOR2_X1 U1066 ( .A(G2090), .B(G2072), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(n978), .B(n977), .ZN(n982) );
  XOR2_X1 U1068 ( .A(G2678), .B(KEYINPUT42), .Z(n980) );
  XNOR2_X1 U1069 ( .A(G2067), .B(KEYINPUT43), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1071 ( .A(n982), .B(n981), .Z(n984) );
  XNOR2_X1 U1072 ( .A(G2078), .B(G2084), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n984), .B(n983), .ZN(G227) );
  NAND2_X1 U1074 ( .A1(G118), .A2(n985), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(G130), .A2(n986), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n995) );
  NAND2_X1 U1077 ( .A1(G106), .A2(n989), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(G142), .A2(n990), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1080 ( .A(KEYINPUT45), .B(n993), .Z(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1000) );
  XOR2_X1 U1082 ( .A(G162), .B(n996), .Z(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(n1000), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1085 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1086 ( .A(n1004), .B(n1003), .ZN(n1010) );
  XOR2_X1 U1087 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1006) );
  XNOR2_X1 U1088 ( .A(G160), .B(G164), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(n1008), .B(n1007), .Z(n1009) );
  XNOR2_X1 U1091 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1011), .ZN(G395) );
  NOR2_X1 U1093 ( .A1(G229), .A2(G227), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(KEYINPUT49), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1095 ( .A1(G397), .A2(n1013), .ZN(n1017) );
  NOR2_X1 U1096 ( .A1(n1018), .A2(G401), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(KEYINPUT116), .B(n1014), .Z(n1015) );
  NOR2_X1 U1098 ( .A1(G395), .A2(n1015), .ZN(n1016) );
  NAND2_X1 U1099 ( .A1(n1017), .A2(n1016), .ZN(G225) );
  INV_X1 U1100 ( .A(G225), .ZN(G308) );
  INV_X1 U1101 ( .A(n1018), .ZN(G319) );
  INV_X1 U1102 ( .A(G108), .ZN(G238) );
endmodule

