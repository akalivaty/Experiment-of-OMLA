//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1252, new_n1253, new_n1254;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT64), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n466), .A2(new_n463), .A3(G101), .A4(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT67), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n469), .A2(new_n470), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n482), .A2(new_n463), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n463), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n463), .A2(KEYINPUT68), .A3(G138), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n482), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(G126), .A3(G2105), .ZN(new_n496));
  AND3_X1   g071(.A1(new_n463), .A2(KEYINPUT68), .A3(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n494), .A2(new_n496), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT69), .A3(G651), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n507), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(G62), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT71), .B1(new_n524), .B2(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  AOI211_X1 g101(.A(new_n526), .B(new_n504), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n525), .A2(new_n527), .B1(KEYINPUT70), .B2(new_n509), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n519), .A2(new_n528), .ZN(G166));
  NAND4_X1  g104(.A1(new_n513), .A2(G51), .A3(G543), .A4(new_n514), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n517), .A2(new_n531), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n530), .B(new_n536), .C1(new_n518), .C2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G168));
  AND2_X1   g116(.A1(new_n508), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n504), .ZN(new_n545));
  INV_X1    g120(.A(new_n518), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G90), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n542), .A2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n504), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n546), .A2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT73), .ZN(G188));
  NAND4_X1  g136(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n508), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n508), .A2(G91), .A3(new_n517), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n515), .B2(new_n516), .ZN(new_n568));
  AND2_X1   g143(.A1(G78), .A2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  AOI22_X1  g147(.A1(new_n546), .A2(G88), .B1(new_n509), .B2(KEYINPUT70), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n524), .A2(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(new_n526), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n524), .A2(KEYINPUT71), .A3(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n510), .A2(new_n511), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(G303));
  NAND3_X1  g154(.A1(new_n508), .A2(G49), .A3(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n508), .A2(G87), .A3(new_n517), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n515), .B2(new_n516), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n513), .A2(G86), .A3(new_n517), .A4(new_n514), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n513), .A2(G48), .A3(G543), .A4(new_n514), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n504), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n599), .B(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(G47), .A2(new_n542), .B1(new_n546), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n520), .A2(new_n521), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n508), .A2(G543), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n546), .A2(KEYINPUT10), .A3(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n518), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n612), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n604), .B1(new_n617), .B2(G868), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NOR2_X1   g194(.A1(G299), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g196(.A(new_n620), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n554), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n617), .A2(new_n623), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g205(.A1(new_n463), .A2(G2104), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n495), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT13), .Z(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT78), .Z(new_n638));
  INV_X1    g213(.A(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n484), .A2(G135), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n641), .A2(new_n642), .B1(new_n644), .B2(G2105), .ZN(new_n645));
  AOI22_X1  g220(.A1(new_n486), .A2(G123), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g222(.A1(new_n635), .A2(new_n636), .B1(new_n639), .B2(new_n647), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n638), .B(new_n648), .C1(new_n639), .C2(new_n647), .ZN(G156));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2430), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n660), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT82), .Z(G401));
  INV_X1    g241(.A(KEYINPUT18), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n636), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n639), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n690), .B(new_n689), .S(new_n682), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1981), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n693), .A2(G1986), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n694), .B2(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n680), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n703), .A2(new_n699), .A3(new_n679), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(G229));
  INV_X1    g280(.A(G29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G32), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n486), .A2(G129), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G141), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT26), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n714), .A2(new_n715), .B1(G105), .B2(new_n631), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n707), .B1(new_n717), .B2(new_n706), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1961), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(G1961), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n718), .A2(new_n720), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n721), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT84), .B(G29), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G27), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(G26), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n484), .A2(G140), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G116), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G2105), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n486), .B2(G128), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(new_n706), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n730), .A2(G35), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n730), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2090), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n734), .B1(new_n745), .B2(G2067), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n647), .A2(new_n730), .ZN(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n745), .A2(G2067), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT24), .B(G34), .ZN(new_n761));
  AOI22_X1  g336(.A1(G160), .A2(G29), .B1(new_n729), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n751), .A2(new_n759), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n728), .A2(new_n750), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G168), .A2(G16), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(KEYINPUT91), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G16), .B2(G21), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n768), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n495), .A2(G127), .ZN(new_n774));
  NAND2_X1  g349(.A1(G115), .A2(G2104), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n463), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n480), .A2(new_n483), .A3(G139), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(KEYINPUT89), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n777), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n776), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G29), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G29), .B2(G33), .ZN(new_n786));
  INV_X1    g361(.A(G2072), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g364(.A1(G299), .A2(G16), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n722), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT23), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n788), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n722), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n617), .B2(new_n722), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1348), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n722), .A2(G19), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT87), .Z(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n554), .B2(G16), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1341), .Z(new_n802));
  NOR2_X1   g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n766), .A2(new_n773), .A3(new_n795), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n484), .A2(G131), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G107), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(G2105), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n486), .B2(G119), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G25), .B(new_n810), .S(new_n730), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT35), .B(G1991), .Z(new_n812));
  XOR2_X1   g387(.A(new_n811), .B(new_n812), .Z(new_n813));
  OR2_X1    g388(.A1(G16), .A2(G24), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT85), .ZN(new_n815));
  XNOR2_X1  g390(.A(G290), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n814), .B1(new_n816), .B2(new_n722), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G1986), .ZN(new_n818));
  INV_X1    g393(.A(G1986), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n819), .B(new_n814), .C1(new_n816), .C2(new_n722), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n813), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G6), .A2(G16), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT86), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT32), .B(G1981), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n722), .A2(G23), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n584), .B2(new_n722), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT33), .B(G1976), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(G16), .A2(G22), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G166), .B2(G16), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n831), .A2(new_n832), .B1(new_n834), .B2(G1971), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(G1971), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT34), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(KEYINPUT34), .B1(new_n827), .B2(new_n837), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n821), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n821), .A2(new_n840), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n804), .B1(new_n843), .B2(new_n845), .ZN(G311));
  NOR2_X1   g421(.A1(G311), .A2(KEYINPUT93), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT93), .ZN(new_n848));
  AOI211_X1 g423(.A(new_n848), .B(new_n804), .C1(new_n843), .C2(new_n845), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(G150));
  NAND2_X1  g425(.A1(new_n542), .A2(G55), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n504), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n546), .A2(G93), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n617), .A2(G559), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT38), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(KEYINPUT94), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n851), .A2(new_n853), .A3(new_n854), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n555), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n555), .B1(new_n860), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n859), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n857), .B1(new_n868), .B2(new_n870), .ZN(G145));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n717), .B1(new_n784), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n874));
  INV_X1    g449(.A(new_n783), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n782), .B1(new_n777), .B2(new_n779), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g452(.A(KEYINPUT96), .B(new_n874), .C1(new_n877), .C2(new_n776), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n873), .A2(new_n878), .A3(new_n743), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n743), .B1(new_n873), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n501), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n744), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n873), .A2(new_n878), .A3(new_n743), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(G164), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n634), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(new_n805), .A3(new_n809), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n805), .B2(new_n809), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n484), .A2(G142), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n463), .A2(G118), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(KEYINPUT97), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n891), .B2(KEYINPUT97), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n892), .A2(new_n894), .B1(new_n486), .B2(G130), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n888), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n896), .B1(new_n888), .B2(new_n889), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(KEYINPUT98), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n901));
  INV_X1    g476(.A(new_n896), .ZN(new_n902));
  INV_X1    g477(.A(new_n889), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n887), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n881), .A2(new_n885), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n881), .B2(new_n885), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT99), .A4(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G160), .B(KEYINPUT95), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(new_n490), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n647), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n881), .A2(new_n885), .A3(new_n898), .A4(new_n899), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n881), .A2(new_n885), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n915), .B(new_n918), .C1(new_n919), .C2(new_n906), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT40), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n915), .B1(new_n910), .B2(new_n911), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n921), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n923), .A2(new_n927), .ZN(G395));
  NAND2_X1  g503(.A1(new_n855), .A2(new_n625), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n627), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n866), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n930), .B(new_n932), .C1(new_n864), .C2(new_n865), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n617), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(G299), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n566), .A2(new_n570), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n940), .A2(new_n564), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n617), .A2(new_n941), .A3(new_n565), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT41), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n936), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n934), .A2(new_n944), .A3(new_n935), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(G290), .B(new_n584), .ZN(new_n949));
  XNOR2_X1  g524(.A(G303), .B(G305), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G290), .B(new_n583), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(KEYINPUT101), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(KEYINPUT101), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n956), .A2(KEYINPUT101), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n952), .A2(new_n954), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n948), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n960), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n947), .A3(new_n946), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n929), .B1(new_n964), .B2(new_n625), .ZN(G295));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n929), .C1(new_n964), .C2(new_n625), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n625), .B1(new_n961), .B2(new_n963), .ZN(new_n968));
  INV_X1    g543(.A(new_n929), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT102), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(G331));
  NAND3_X1  g546(.A1(G171), .A2(new_n539), .A3(new_n540), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G171), .B1(new_n539), .B2(new_n540), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n864), .A2(new_n865), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n860), .A2(new_n862), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n554), .ZN(new_n977));
  NAND2_X1  g552(.A1(G168), .A2(G301), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n863), .A3(new_n978), .A4(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n945), .A2(new_n943), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n975), .A2(new_n979), .A3(new_n938), .A4(new_n942), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n955), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n982), .A2(new_n955), .A3(KEYINPUT105), .A4(new_n983), .ZN(new_n987));
  INV_X1    g562(.A(new_n955), .ZN(new_n988));
  INV_X1    g563(.A(new_n983), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n979), .A2(new_n975), .B1(new_n945), .B2(new_n943), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n986), .A2(new_n921), .A3(new_n987), .A4(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n987), .A2(new_n921), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n945), .A2(new_n943), .A3(KEYINPUT106), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n980), .C1(KEYINPUT106), .C2(new_n945), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n983), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n988), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n996), .A2(new_n986), .A3(new_n1000), .A4(new_n993), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n995), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n996), .A2(new_n986), .A3(new_n1000), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n996), .A2(new_n986), .A3(new_n991), .A4(new_n993), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(KEYINPUT44), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(G397));
  XNOR2_X1  g584(.A(new_n874), .B(G1996), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n743), .B(G2067), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n810), .B(new_n812), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n501), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n479), .A2(G137), .B1(new_n465), .B2(new_n467), .ZN(new_n1019));
  INV_X1    g594(.A(G125), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n477), .B2(new_n478), .ZN(new_n1021));
  INV_X1    g596(.A(new_n474), .ZN(new_n1022));
  OAI21_X1  g597(.A(G2105), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT107), .B(G40), .Z(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1018), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1014), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G290), .A2(G1986), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n1029), .B(KEYINPUT108), .Z(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(G1986), .B2(G290), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1027), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1956), .ZN(new_n1036));
  NOR2_X1   g611(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n501), .A2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n472), .A2(new_n475), .A3(new_n1024), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n501), .B2(new_n1015), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1036), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1017), .A2(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1026), .B1(new_n501), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1018), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n940), .A2(new_n1050), .A3(new_n565), .A4(new_n564), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT120), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1039), .A2(new_n1059), .A3(new_n1015), .A4(new_n501), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2067), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n1064));
  INV_X1    g639(.A(G1348), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1026), .B1(new_n501), .B2(new_n1037), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1063), .A2(new_n1064), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G2067), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT119), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(new_n937), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1057), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  NAND3_X1  g651(.A1(new_n1058), .A2(new_n1060), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1996), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1045), .A2(new_n1018), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n554), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1069), .A2(KEYINPUT60), .A3(new_n937), .A4(new_n1071), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT121), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1043), .A4(new_n1047), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1084), .A2(new_n1056), .A3(KEYINPUT61), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1085), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1073), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1082), .A2(new_n1083), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1071), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1068), .A2(new_n1065), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1070), .B2(KEYINPUT119), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1098), .A2(KEYINPUT60), .A3(new_n1071), .A4(new_n1095), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(new_n617), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1075), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n580), .A2(new_n581), .A3(G1976), .A4(new_n582), .ZN(new_n1103));
  OAI211_X1 g678(.A(G8), .B(new_n1103), .C1(new_n1016), .C2(new_n1026), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(KEYINPUT112), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1039), .A2(new_n1015), .A3(new_n501), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(G8), .A4(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT113), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1105), .A2(new_n1111), .A3(new_n1108), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1114));
  OAI211_X1 g689(.A(G8), .B(new_n1114), .C1(new_n519), .C2(new_n528), .ZN(new_n1115));
  INV_X1    g690(.A(G8), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n575), .A2(new_n576), .B1(new_n510), .B2(new_n511), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1116), .B1(new_n1117), .B2(new_n573), .ZN(new_n1118));
  XOR2_X1   g693(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1971), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n501), .A2(new_n1044), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1039), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT45), .B1(new_n501), .B2(new_n1015), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1040), .A2(G2090), .A3(new_n1042), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(KEYINPUT110), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT110), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1068), .A2(new_n1128), .A3(G2090), .ZN(new_n1129));
  OAI211_X1 g704(.A(G8), .B(new_n1120), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(G61), .B1(new_n520), .B2(new_n521), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n504), .B1(new_n1131), .B2(new_n592), .ZN(new_n1132));
  OAI21_X1  g707(.A(G1981), .B1(new_n1132), .B2(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n823), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1981), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n594), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G305), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT49), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(G8), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1134), .A2(new_n1138), .A3(KEYINPUT49), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1143));
  INV_X1    g718(.A(G1976), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n585), .A2(new_n1144), .A3(new_n587), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1115), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1119), .B1(G303), .B2(G8), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(G1971), .B1(new_n1045), .B2(new_n1018), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1150), .B2(new_n1126), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1113), .A2(new_n1130), .A3(new_n1146), .A4(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n772), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1066), .A2(new_n1067), .A3(new_n763), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(new_n1155), .A3(G168), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT51), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1156), .A2(new_n1157), .A3(G8), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G286), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(G8), .A3(new_n1156), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1161), .B2(KEYINPUT51), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1045), .A2(new_n1018), .A3(new_n733), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1961), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1068), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1045), .A2(new_n1018), .A3(KEYINPUT53), .A4(new_n733), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(G171), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n473), .A2(new_n474), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n463), .B1(new_n1171), .B2(KEYINPUT122), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(KEYINPUT122), .B2(new_n1171), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n733), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n472), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1018), .A2(new_n1122), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1165), .A2(new_n1167), .A3(G301), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT54), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1153), .A2(new_n1162), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1165), .A2(new_n1167), .A3(new_n1176), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(G171), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1181), .B(KEYINPUT54), .C1(G171), .C2(new_n1169), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(KEYINPUT123), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1169), .A2(G171), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT54), .A4(new_n1181), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1101), .A2(new_n1179), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1189), .A2(new_n1144), .A3(new_n588), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n823), .A2(new_n1135), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1140), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT115), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1113), .B2(new_n1146), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1105), .A2(new_n1111), .A3(new_n1108), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1111), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1146), .B(new_n1193), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1130), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1192), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1156), .A2(G8), .ZN(new_n1203));
  AOI21_X1  g778(.A(G168), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1204));
  OAI21_X1  g779(.A(KEYINPUT51), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1156), .A2(new_n1157), .A3(G8), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1206), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1130), .A2(new_n1152), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1146), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1211), .A2(new_n1212), .A3(new_n1170), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1202), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1162), .A2(new_n1206), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(KEYINPUT62), .ZN(new_n1217));
  AND4_X1   g792(.A1(new_n1202), .A2(new_n1213), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1188), .B(new_n1201), .C1(new_n1214), .C2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1153), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1159), .A2(G8), .A3(G168), .ZN(new_n1221));
  AND2_X1   g796(.A1(new_n1221), .A2(KEYINPUT116), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1221), .A2(KEYINPUT116), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g799(.A(KEYINPUT63), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g800(.A(KEYINPUT63), .B(new_n1130), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1226));
  OAI21_X1  g801(.A(G8), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1149), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1228), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT117), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1226), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1199), .A2(KEYINPUT117), .A3(new_n1228), .ZN(new_n1232));
  AOI21_X1  g807(.A(new_n1225), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1035), .B1(new_n1219), .B2(new_n1233), .ZN(new_n1234));
  AND2_X1   g809(.A1(new_n1030), .A2(new_n1027), .ZN(new_n1235));
  OR2_X1    g810(.A1(new_n1235), .A2(KEYINPUT48), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(KEYINPUT48), .ZN(new_n1237));
  NAND3_X1  g812(.A1(new_n1236), .A2(new_n1028), .A3(new_n1237), .ZN(new_n1238));
  NAND4_X1  g813(.A1(new_n1012), .A2(new_n812), .A3(new_n805), .A4(new_n809), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n744), .A2(new_n1062), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1032), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(KEYINPUT125), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1027), .A2(new_n1078), .ZN(new_n1243));
  XNOR2_X1  g818(.A(new_n1243), .B(KEYINPUT46), .ZN(new_n1244));
  OAI21_X1  g819(.A(new_n1027), .B1(new_n1011), .B2(new_n874), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  XNOR2_X1  g821(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1247));
  XNOR2_X1  g822(.A(new_n1246), .B(new_n1247), .ZN(new_n1248));
  AND3_X1   g823(.A1(new_n1238), .A2(new_n1242), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1234), .A2(new_n1249), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g825(.A1(new_n917), .A2(new_n922), .ZN(new_n1252));
  OR3_X1    g826(.A1(new_n665), .A2(new_n461), .A3(G227), .ZN(new_n1253));
  AOI21_X1  g827(.A(new_n1253), .B1(new_n702), .B2(new_n704), .ZN(new_n1254));
  AND3_X1   g828(.A1(new_n1252), .A2(new_n1254), .A3(new_n1002), .ZN(G308));
  NAND3_X1  g829(.A1(new_n1252), .A2(new_n1254), .A3(new_n1002), .ZN(G225));
endmodule


