//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT64), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(KEYINPUT66), .A3(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n462), .A2(new_n463), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  AOI21_X1  g051(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT67), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n481), .B1(new_n483), .B2(G136), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n461), .B2(G114), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n486), .A2(new_n488), .A3(new_n489), .A4(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(KEYINPUT69), .A3(new_n491), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n466), .B2(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n467), .C2(new_n466), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n461), .A2(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n464), .A2(new_n468), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n494), .A2(new_n495), .B1(new_n502), .B2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n510), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(G166));
  NAND3_X1  g099(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n526), .A2(new_n528), .A3(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AND4_X1   g109(.A1(new_n513), .A2(new_n515), .A3(new_n526), .A4(new_n528), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(new_n530), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n517), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n522), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n535), .A2(G81), .B1(new_n530), .B2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n513), .A2(new_n515), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT73), .ZN(G188));
  AOI21_X1  g133(.A(KEYINPUT76), .B1(new_n513), .B2(new_n515), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT76), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G65), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n522), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g141(.A(G53), .B1(new_n566), .B2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n529), .A2(new_n567), .B1(new_n568), .B2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(new_n567), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n568), .A2(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n570), .A2(new_n507), .A3(G543), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n535), .A2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G168), .ZN(G286));
  OAI221_X1 g154(.A(new_n510), .B1(new_n511), .B2(new_n517), .C1(new_n522), .C2(new_n521), .ZN(G303));
  AND3_X1   g155(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT77), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n535), .A2(G87), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  INV_X1    g161(.A(G48), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n517), .A2(new_n586), .B1(new_n587), .B2(new_n529), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n516), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n522), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n535), .A2(G85), .B1(new_n530), .B2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n547), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n595), .B1(new_n599), .B2(KEYINPUT79), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n598), .A2(KEYINPUT79), .A3(G651), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n600), .A2(KEYINPUT80), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT80), .B1(new_n600), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n535), .A2(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n606), .B(KEYINPUT81), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n560), .A2(G66), .A3(new_n561), .ZN(new_n613));
  INV_X1    g188(.A(G79), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(new_n514), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n615), .A2(G651), .B1(G54), .B2(new_n530), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n609), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n605), .B1(new_n618), .B2(G868), .ZN(G321));
  XOR2_X1   g194(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n576), .ZN(G297));
  XOR2_X1   g198(.A(G297), .B(KEYINPUT84), .Z(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  OR3_X1    g201(.A1(new_n617), .A2(KEYINPUT85), .A3(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT85), .B1(new_n617), .B2(G559), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(G868), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n551), .A2(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT11), .Z(G282));
  INV_X1    g207(.A(new_n631), .ZN(G323));
  AND2_X1   g208(.A1(new_n464), .A2(new_n468), .ZN(new_n634));
  INV_X1    g209(.A(G2104), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n635), .A2(G2105), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n461), .A2(G111), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT87), .Z(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n644), .B1(KEYINPUT88), .B2(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(KEYINPUT88), .ZN(new_n648));
  INV_X1    g223(.A(new_n477), .ZN(new_n649));
  INV_X1    g224(.A(G123), .ZN(new_n650));
  OR3_X1    g225(.A1(new_n649), .A2(KEYINPUT86), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(KEYINPUT86), .B1(new_n649), .B2(new_n650), .ZN(new_n652));
  AOI22_X1  g227(.A1(new_n647), .A2(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n483), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n641), .A2(new_n642), .A3(new_n657), .ZN(G156));
  XOR2_X1   g233(.A(KEYINPUT15), .B(G2435), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XOR2_X1   g235(.A(G2427), .B(G2430), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT89), .B(KEYINPUT14), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1341), .B(G1348), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT90), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(G14), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(G401));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT17), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n679), .A2(new_n677), .A3(new_n680), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n677), .A3(new_n680), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT18), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n656), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(G227));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n691), .B2(new_n692), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT93), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n694), .A2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT20), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n695), .A2(new_n699), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n700), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(G1981), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n708), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G1971), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n714), .A2(G23), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G288), .B2(G16), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT33), .B(G1976), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n714), .A2(G6), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n593), .B2(new_n714), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n719), .A2(new_n720), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n716), .B2(G1971), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n721), .A2(new_n725), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT34), .Z(new_n730));
  MUX2_X1   g305(.A(G24), .B(G290), .S(G16), .Z(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1986), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G25), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT94), .Z(new_n735));
  OR2_X1    g310(.A1(G95), .A2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G107), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n635), .B1(new_n737), .B2(G2105), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n477), .A2(G119), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n483), .B2(G131), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT35), .B(G1991), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n742), .B(new_n744), .Z(new_n745));
  NAND3_X1  g320(.A1(new_n730), .A2(new_n732), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n733), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n733), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G2090), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n714), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT23), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n576), .B2(new_n714), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n733), .A2(G33), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT25), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n634), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n461), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(G139), .C2(new_n483), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n733), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2072), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n714), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1966), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT31), .B(G11), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT103), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(G28), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(G28), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n551), .A2(G16), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n714), .A2(G19), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n775), .B1(new_n733), .B2(new_n655), .C1(new_n779), .C2(G1341), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n766), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G164), .A2(new_n733), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G27), .B2(new_n733), .ZN(new_n783));
  INV_X1    g358(.A(G2078), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n733), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G2084), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n783), .A2(new_n784), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(G2084), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n785), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n714), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n714), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n779), .A2(G1341), .B1(G1961), .B2(new_n796), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n797), .B1(G1961), .B2(new_n796), .C1(new_n750), .C2(G2090), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n781), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n733), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT100), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT28), .ZN(new_n802));
  NOR2_X1   g377(.A1(G104), .A2(G2105), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT98), .Z(new_n804));
  INV_X1    g379(.A(G116), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n635), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n804), .A2(new_n806), .B1(G128), .B2(new_n477), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n483), .A2(KEYINPUT97), .A3(G140), .ZN(new_n808));
  AOI21_X1  g383(.A(KEYINPUT97), .B1(new_n483), .B2(G140), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G29), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(KEYINPUT99), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n483), .A2(G141), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT101), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT26), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n477), .A2(G129), .B1(G105), .B2(new_n636), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n733), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT102), .Z(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G29), .B2(G32), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT27), .B(G1996), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(G4), .A2(G16), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n617), .B2(new_n714), .ZN(new_n830));
  INV_X1    g405(.A(G1348), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  AND4_X1   g408(.A1(new_n758), .A2(new_n799), .A3(new_n816), .A4(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n747), .A2(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n747), .A2(new_n834), .ZN(G150));
  NAND2_X1  g411(.A1(new_n530), .A2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n517), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n516), .A2(G67), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n522), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n551), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n552), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n618), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT105), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n843), .A2(G860), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT37), .Z(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  INV_X1    g432(.A(new_n741), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n822), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n503), .B1(new_n462), .B2(new_n463), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT4), .B1(new_n861), .B2(new_n500), .ZN(new_n862));
  INV_X1    g437(.A(new_n501), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n505), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n492), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n810), .B(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n764), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n477), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(G106), .A2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n483), .B2(G142), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n638), .B(new_n873), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n868), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n868), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n859), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n655), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  AOI21_X1  g459(.A(G37), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n884), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n878), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT40), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G395));
  NAND2_X1  g465(.A1(new_n617), .A2(new_n576), .ZN(new_n891));
  NAND4_X1  g466(.A1(G299), .A2(new_n609), .A3(new_n612), .A4(new_n616), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT41), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n844), .A2(new_n846), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n627), .A2(new_n628), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n627), .B2(new_n628), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n891), .A2(new_n892), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT108), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G303), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n593), .A2(new_n603), .A3(new_n602), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n593), .B1(new_n603), .B2(new_n602), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G305), .A2(G290), .ZN(new_n911));
  XNOR2_X1  g486(.A(G303), .B(G288), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(KEYINPUT107), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n908), .A2(new_n909), .A3(new_n906), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n912), .B1(new_n911), .B2(new_n907), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n917), .A2(KEYINPUT107), .B1(new_n921), .B2(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n901), .A2(KEYINPUT108), .A3(new_n903), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n904), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND4_X1   g501(.A1(new_n904), .A2(new_n925), .A3(new_n918), .A4(new_n922), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n845), .ZN(G331));
  XNOR2_X1  g505(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G171), .B(G168), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n897), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n902), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n847), .A3(KEYINPUT110), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n933), .B(new_n847), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(KEYINPUT110), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n921), .B(new_n935), .C1(new_n896), .C2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n934), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n895), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n893), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n944), .A2(new_n946), .B1(new_n902), .B2(new_n934), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(new_n921), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n932), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n947), .B2(new_n921), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n938), .A2(new_n902), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n894), .A2(new_n895), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n937), .B1(new_n945), .B2(KEYINPUT111), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n914), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n950), .A2(new_n956), .A3(new_n931), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n949), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n934), .B1(new_n952), .B2(new_n895), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n945), .A2(KEYINPUT111), .A3(new_n893), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n960), .A2(new_n961), .B1(new_n938), .B2(new_n902), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n939), .B(new_n940), .C1(new_n962), .C2(new_n921), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n935), .B1(new_n896), .B2(new_n938), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n914), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n950), .A2(new_n931), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n958), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n959), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n949), .A2(new_n957), .A3(new_n958), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n941), .A2(new_n948), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n972), .A2(new_n931), .B1(new_n963), .B2(KEYINPUT43), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n970), .B(new_n971), .C1(new_n973), .C2(new_n958), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(G397));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n864), .B2(new_n865), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT45), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n810), .B(new_n815), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(new_n822), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n984));
  INV_X1    g559(.A(new_n978), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(G1996), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n822), .B(G1996), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n741), .B(new_n744), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n978), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  NOR3_X1   g569(.A1(G290), .A2(new_n985), .A3(G1986), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT48), .Z(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n858), .A2(new_n744), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(new_n990), .B2(new_n985), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n810), .A2(G2067), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(KEYINPUT126), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT126), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n985), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT63), .ZN(new_n1008));
  INV_X1    g583(.A(G40), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n471), .A2(new_n475), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n977), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT117), .B1(new_n592), .B2(new_n710), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NOR4_X1   g590(.A1(new_n588), .A2(new_n591), .A3(new_n1015), .A4(G1981), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1014), .A2(new_n1016), .B1(new_n710), .B2(new_n592), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1013), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n1018), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n905), .A2(new_n1025), .A3(G1976), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT116), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n1029), .B2(new_n1012), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1013), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n905), .B2(G1976), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1024), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT45), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(G164), .B2(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1010), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT113), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n866), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT114), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n977), .A2(new_n1057), .A3(new_n1053), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1056), .A2(new_n1010), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1050), .B(new_n1052), .C1(G2090), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1043), .A2(new_n1061), .A3(G8), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1010), .B1(new_n977), .B2(new_n1053), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n494), .A2(new_n495), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT50), .B(G1384), .C1(new_n1065), .C2(new_n864), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1064), .A2(new_n1066), .A3(G2090), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1042), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1035), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT119), .B(G2084), .Z(new_n1071));
  NOR2_X1   g646(.A1(new_n976), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1056), .A2(new_n1072), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1010), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n1075));
  NOR3_X1   g650(.A1(G164), .A2(new_n1044), .A3(G1384), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(G8), .A3(G168), .ZN(new_n1079));
  XOR2_X1   g654(.A(new_n1079), .B(KEYINPUT120), .Z(new_n1080));
  OAI21_X1  g655(.A(new_n1008), .B1(new_n1070), .B2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1079), .A2(KEYINPUT120), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(KEYINPUT120), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1008), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1061), .A2(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1042), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(new_n1086), .A3(new_n1062), .A4(new_n1035), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1062), .A2(new_n1024), .A3(new_n1034), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n905), .A2(new_n1027), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1024), .A2(new_n1090), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1091), .B2(new_n1013), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1078), .A2(KEYINPUT124), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1073), .A2(new_n1077), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G168), .A2(new_n1063), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1078), .A2(G286), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G8), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1097), .A2(new_n1099), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G286), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT51), .B1(new_n1105), .B2(new_n1063), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1096), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1095), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1110));
  OAI21_X1  g685(.A(G168), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1101), .B1(new_n1111), .B2(G8), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT62), .B1(new_n1112), .B2(new_n1103), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1047), .A2(G2078), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  INV_X1    g690(.A(G1961), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1114), .A2(new_n1115), .B1(new_n1116), .B2(new_n1060), .ZN(new_n1117));
  OR4_X1    g692(.A1(new_n1115), .A2(new_n1075), .A3(new_n1076), .A4(G2078), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1108), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n565), .A2(new_n575), .A3(KEYINPUT121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT76), .ZN(new_n1124));
  INV_X1    g699(.A(G65), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n559), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n564), .ZN(new_n1127));
  OAI21_X1  g702(.A(G651), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n569), .A2(new_n572), .B1(new_n535), .B2(G91), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1121), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n565), .B2(new_n575), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n755), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT56), .B(G2072), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1045), .A2(new_n1046), .A3(new_n1010), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1060), .A2(new_n831), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1011), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n815), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n618), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT57), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1144), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1142), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n618), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n617), .A4(new_n1142), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n1149), .B2(new_n1139), .ZN(new_n1157));
  OAI21_X1  g732(.A(KEYINPUT122), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1135), .A2(new_n1160), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1045), .A2(new_n1046), .A3(new_n982), .A4(new_n1010), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT58), .B(G1341), .Z(new_n1164));
  NAND2_X1  g739(.A1(new_n1011), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n551), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1166), .B(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1157), .A2(new_n1162), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1155), .B1(new_n1169), .B2(KEYINPUT123), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1157), .A2(new_n1162), .A3(new_n1168), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1150), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1117), .A2(G301), .A3(new_n1118), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1046), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1175), .A2(new_n1075), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1117), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(KEYINPUT54), .B(new_n1174), .C1(new_n1177), .C2(G301), .ZN(new_n1178));
  XOR2_X1   g753(.A(KEYINPUT125), .B(KEYINPUT54), .Z(new_n1179));
  AND3_X1   g754(.A1(new_n1117), .A2(G301), .A3(new_n1176), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(new_n1119), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1178), .B(new_n1181), .C1(new_n1112), .C2(new_n1103), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1120), .B1(new_n1173), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1070), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1093), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n992), .ZN(new_n1186));
  XOR2_X1   g761(.A(G290), .B(G1986), .Z(new_n1187));
  AOI21_X1  g762(.A(new_n985), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1007), .B1(new_n1185), .B2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g764(.A(new_n459), .B(G227), .C1(new_n673), .C2(new_n675), .ZN(new_n1191));
  AND2_X1   g765(.A1(new_n712), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n885), .A2(new_n887), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n957), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(G308));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(G225));
endmodule


