//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n187));
  NOR2_X1   g001(.A1(G475), .A2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT93), .Z(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT69), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G237), .ZN(new_n195));
  AND4_X1   g009(.A1(G143), .A2(new_n194), .A3(G214), .A4(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(G237), .B1(new_n191), .B2(new_n193), .ZN(new_n197));
  AOI21_X1  g011(.A(G143), .B1(new_n197), .B2(G214), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(G214), .A3(new_n195), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n197), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n199), .A2(new_n200), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT79), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(KEYINPUT16), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n214), .A2(new_n211), .A3(KEYINPUT79), .A4(G125), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n209), .A2(G146), .A3(new_n213), .A4(new_n215), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n204), .B1(new_n203), .B2(new_n205), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G113), .B(G122), .ZN(new_n224));
  INV_X1    g038(.A(G104), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n203), .B(new_n205), .C1(new_n204), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G125), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G140), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n208), .A2(new_n217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n228), .B(new_n234), .C1(new_n199), .C2(new_n227), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n223), .A2(new_n226), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT91), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n223), .A2(new_n238), .A3(new_n226), .A4(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n199), .A2(new_n206), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT90), .B1(new_n231), .B2(KEYINPUT19), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT19), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n208), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT89), .B1(new_n208), .B2(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(new_n247), .A3(KEYINPUT19), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n242), .A2(new_n245), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n217), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n219), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n226), .B1(new_n251), .B2(new_n235), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n240), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT92), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n189), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n187), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n189), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n240), .B2(new_n253), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT92), .B(new_n252), .C1(new_n237), .C2(new_n239), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n189), .A2(KEYINPUT20), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n240), .B2(new_n253), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n190), .A2(G952), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(G234), .B2(G237), .ZN(new_n272));
  INV_X1    g086(.A(new_n194), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n274), .B1(G234), .B2(G237), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n276), .B(KEYINPUT98), .Z(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT21), .B(G898), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G128), .B(G143), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT14), .A3(G122), .ZN(new_n285));
  XNOR2_X1  g099(.A(G116), .B(G122), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(G107), .B(new_n285), .C1(new_n287), .C2(KEYINPUT14), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n283), .B(new_n288), .C1(G107), .C2(new_n287), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n202), .A2(G128), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n290), .A2(KEYINPUT13), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n282), .B(new_n291), .C1(KEYINPUT13), .C2(new_n281), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT96), .ZN(new_n293));
  INV_X1    g107(.A(G107), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n286), .B(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n281), .A2(new_n282), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n289), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT77), .B(G217), .Z(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT9), .B(G234), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n300), .A2(new_n302), .A3(G953), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n298), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n274), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT97), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT15), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G478), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n309), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n226), .B1(new_n223), .B2(new_n235), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT95), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n240), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n274), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G475), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n270), .A2(new_n280), .A3(new_n312), .A4(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n225), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n294), .A3(G104), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n225), .A2(G107), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G119), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT2), .B(G113), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n328), .A2(KEYINPUT4), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n323), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n225), .A2(G107), .ZN(new_n339));
  OAI21_X1  g153(.A(G101), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT5), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G116), .ZN(new_n343));
  OAI211_X1 g157(.A(G113), .B(new_n343), .C1(new_n331), .C2(new_n341), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n326), .A2(new_n333), .A3(new_n340), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G122), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n345), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n217), .B2(G143), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n202), .A2(KEYINPUT65), .A3(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(KEYINPUT0), .A2(G128), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n202), .A2(G146), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  OR2_X1    g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n217), .A2(G143), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n356), .B(new_n361), .C1(new_n358), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n358), .B1(new_n353), .B2(new_n354), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G128), .ZN(new_n368));
  OAI21_X1  g182(.A(G128), .B1(new_n358), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n358), .B2(new_n362), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(new_n229), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n190), .A2(G224), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n346), .A2(new_n375), .A3(new_n348), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n351), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT85), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n365), .A2(new_n371), .B1(KEYINPUT7), .B2(new_n373), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n365), .A2(KEYINPUT84), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT84), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n381), .B1(new_n372), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n347), .B(KEYINPUT8), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n326), .A2(new_n340), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n344), .A2(new_n333), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n385), .B1(new_n388), .B2(new_n345), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n378), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n345), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n384), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n372), .A2(new_n382), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(KEYINPUT85), .A3(new_n393), .A4(new_n381), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n394), .A3(new_n350), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n377), .A2(new_n395), .A3(new_n274), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT86), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  INV_X1    g214(.A(new_n398), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n377), .A2(new_n395), .A3(new_n274), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(G214), .B1(G237), .B2(G902), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n398), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n318), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT32), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n368), .A2(new_n370), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n282), .B2(G137), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n282), .A2(G137), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n410), .B(new_n414), .C1(new_n282), .C2(G137), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n412), .A2(new_n204), .A3(new_n413), .A4(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n413), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n282), .A2(G137), .ZN(new_n418));
  OAI21_X1  g232(.A(G131), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n416), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(KEYINPUT67), .A3(G131), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n420), .B1(new_n426), .B2(new_n364), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT68), .B1(new_n360), .B2(new_n363), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n360), .A2(KEYINPUT68), .A3(new_n363), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n424), .B(new_n425), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n335), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(G101), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n197), .A2(G210), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n335), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n439), .A3(new_n420), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT31), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n443));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n438), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n432), .A2(KEYINPUT28), .A3(new_n439), .A4(new_n420), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n427), .A2(new_n335), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n450));
  INV_X1    g264(.A(new_n438), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n442), .B(new_n444), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G472), .A2(G902), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT72), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n454), .A2(KEYINPUT73), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT73), .B1(new_n454), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n408), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT74), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n432), .A2(new_n420), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n335), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n446), .A2(new_n463), .A3(KEYINPUT29), .A4(new_n447), .ZN(new_n464));
  OR3_X1    g278(.A1(new_n464), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT75), .B1(new_n464), .B2(new_n451), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n274), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT76), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n465), .A2(new_n469), .A3(new_n466), .A4(new_n274), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n434), .A2(new_n440), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n451), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT29), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(new_n473), .C1(new_n451), .C2(new_n449), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n468), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n454), .A2(KEYINPUT32), .A3(new_n457), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT74), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n408), .C1(new_n458), .C2(new_n459), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n461), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT80), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n218), .A2(new_n219), .ZN(new_n482));
  XOR2_X1   g296(.A(KEYINPUT24), .B(G110), .Z(new_n483));
  XNOR2_X1  g297(.A(G119), .B(G128), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT78), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n342), .A2(G128), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n342), .A2(G128), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G110), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n482), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n491), .A2(G110), .B1(new_n484), .B2(new_n483), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n219), .A3(new_n233), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT22), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(G137), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n500), .B(G137), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n481), .B(KEYINPUT25), .C1(new_n505), .C2(G902), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n300), .B1(G234), .B2(new_n274), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT80), .B(KEYINPUT25), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n502), .A2(new_n504), .A3(new_n274), .A4(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n505), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n507), .A2(G902), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n386), .A2(new_n370), .A3(new_n368), .ZN(new_n517));
  INV_X1    g331(.A(new_n369), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n368), .B1(new_n366), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n326), .A2(new_n519), .A3(new_n340), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n426), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n521), .B(KEYINPUT12), .Z(new_n522));
  INV_X1    g336(.A(KEYINPUT10), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT83), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(KEYINPUT83), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n329), .B(new_n336), .C1(new_n430), .C2(new_n431), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n409), .A4(new_n340), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n528), .A2(new_n426), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n194), .A2(G227), .ZN(new_n532));
  XNOR2_X1  g346(.A(G110), .B(G140), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n522), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n527), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT83), .B1(new_n520), .B2(new_n523), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n529), .B(new_n530), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n425), .A3(new_n424), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n534), .B1(new_n540), .B2(new_n531), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n516), .B(new_n274), .C1(new_n536), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n516), .A2(new_n274), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n534), .ZN(new_n545));
  INV_X1    g359(.A(new_n531), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(new_n531), .A3(new_n534), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(G469), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT81), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n407), .A2(new_n480), .A3(new_n515), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(G101), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(G3));
  AOI21_X1  g370(.A(G478), .B1(new_n305), .B2(new_n274), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT101), .B1(new_n305), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n298), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n303), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n298), .A2(new_n560), .A3(new_n304), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT33), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(KEYINPUT101), .A3(KEYINPUT33), .A4(new_n563), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n557), .B1(new_n567), .B2(G478), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n270), .B2(new_n317), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n399), .A2(new_n402), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n404), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n279), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n458), .A2(new_n459), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n454), .A2(new_n274), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G472), .ZN(new_n576));
  AND4_X1   g390(.A1(new_n574), .A2(new_n553), .A3(new_n515), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT34), .B(G104), .Z(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G6));
  NAND2_X1  g394(.A1(new_n310), .A2(new_n311), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n266), .B1(new_n262), .B2(new_n263), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n582), .A2(KEYINPUT102), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(KEYINPUT102), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n260), .A2(new_n583), .A3(new_n265), .A4(new_n584), .ZN(new_n585));
  AND4_X1   g399(.A1(new_n581), .A2(new_n572), .A3(new_n585), .A4(new_n317), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G107), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G9));
  AND2_X1   g403(.A1(new_n574), .A2(new_n576), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT103), .B1(new_n503), .B2(KEYINPUT36), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n501), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n591), .A2(new_n497), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n497), .B1(new_n594), .B2(new_n591), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n512), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n510), .A2(new_n597), .A3(KEYINPUT104), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT104), .B1(new_n510), .B2(new_n597), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n407), .A2(new_n553), .A3(new_n590), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT105), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT37), .B(G110), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G12));
  INV_X1    g418(.A(G900), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n272), .B1(new_n277), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND4_X1   g421(.A1(new_n581), .A2(new_n585), .A3(new_n317), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n550), .A2(new_n552), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n571), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n480), .A2(new_n608), .A3(new_n600), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G128), .ZN(G30));
  XNOR2_X1  g426(.A(new_n606), .B(KEYINPUT39), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n553), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n615), .A2(KEYINPUT40), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n270), .A2(new_n317), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n312), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(KEYINPUT40), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n404), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n471), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n451), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n463), .A2(new_n451), .A3(new_n440), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n274), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n461), .A2(new_n477), .A3(new_n479), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n403), .A2(new_n405), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT38), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n621), .A2(new_n600), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(new_n202), .ZN(G45));
  AOI211_X1 g446(.A(new_n606), .B(new_n568), .C1(new_n270), .C2(new_n317), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n480), .A2(new_n633), .A3(new_n600), .A4(new_n610), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G146), .ZN(G48));
  NAND2_X1  g449(.A1(new_n480), .A2(new_n515), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n274), .B1(new_n536), .B2(new_n541), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(G469), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n552), .A3(new_n542), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n573), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT41), .B(G113), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G15));
  NAND4_X1  g457(.A1(new_n480), .A2(new_n586), .A3(new_n515), .A4(new_n640), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G116), .ZN(G18));
  AND2_X1   g459(.A1(new_n480), .A2(new_n600), .ZN(new_n646));
  INV_X1    g460(.A(new_n318), .ZN(new_n647));
  INV_X1    g461(.A(new_n404), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n399), .B2(new_n402), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n639), .A3(new_n552), .A4(new_n542), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G119), .ZN(G21));
  INV_X1    g467(.A(new_n576), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n446), .A2(new_n447), .A3(new_n463), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n442), .B(new_n444), .C1(new_n438), .C2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n457), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n654), .A2(new_n514), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n619), .A2(new_n280), .A3(new_n651), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G122), .ZN(G24));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n661));
  INV_X1    g475(.A(new_n568), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n264), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT94), .B1(new_n264), .B2(KEYINPUT20), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n664), .A3(new_n268), .ZN(new_n665));
  INV_X1    g479(.A(new_n317), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n662), .B(new_n607), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n657), .B1(G472), .B2(new_n575), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n640), .A2(new_n668), .A3(new_n649), .A4(new_n600), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n661), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n657), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n600), .A2(new_n576), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n650), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(new_n569), .A3(KEYINPUT106), .A4(new_n607), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G125), .ZN(G27));
  NAND2_X1  g490(.A1(new_n629), .A2(new_n404), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n609), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n569), .A3(new_n607), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n454), .A2(new_n457), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n408), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n476), .A2(new_n477), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n515), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT42), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n633), .A2(new_n685), .A3(new_n678), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n684), .B1(new_n636), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n204), .ZN(G33));
  NAND3_X1  g502(.A1(new_n637), .A2(new_n608), .A3(new_n678), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G134), .ZN(G36));
  NOR3_X1   g504(.A1(new_n617), .A2(KEYINPUT43), .A3(new_n568), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n617), .A2(KEYINPUT108), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n617), .A2(KEYINPUT108), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n662), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n691), .B1(new_n695), .B2(KEYINPUT43), .ZN(new_n696));
  INV_X1    g510(.A(new_n590), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(new_n600), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT109), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n547), .A2(new_n548), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT107), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n706), .A3(G469), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n543), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n708), .A2(KEYINPUT46), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n542), .B1(new_n708), .B2(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n552), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(new_n613), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n677), .B1(new_n698), .B2(new_n699), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n701), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G137), .ZN(G39));
  INV_X1    g530(.A(KEYINPUT47), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT47), .B(new_n552), .C1(new_n709), .C2(new_n710), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n667), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n677), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n480), .A2(new_n515), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G140), .ZN(G42));
  NAND2_X1  g538(.A1(new_n639), .A2(new_n542), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n718), .B(new_n719), .C1(new_n552), .C2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n691), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n568), .B1(new_n692), .B2(new_n693), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n272), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n658), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n726), .A2(new_n721), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n721), .A2(new_n640), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n627), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n515), .A2(new_n272), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n735), .A2(KEYINPUT117), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT117), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n617), .A4(new_n662), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n740));
  INV_X1    g554(.A(new_n734), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n696), .A2(new_n740), .A3(new_n272), .A4(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT116), .B1(new_n730), .B2(new_n734), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n672), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n739), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n630), .A2(new_n648), .A3(new_n640), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n730), .A2(new_n731), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n747), .A2(new_n748), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n751), .B2(new_n755), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n733), .B(new_n746), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n683), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT119), .B1(new_n744), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n764), .B(new_n683), .C1(new_n742), .C2(new_n743), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n271), .B1(new_n766), .B2(KEYINPUT48), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n746), .B(KEYINPUT118), .C1(new_n757), .C2(new_n758), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n733), .ZN(new_n769));
  INV_X1    g583(.A(new_n758), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n756), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT118), .B1(new_n771), .B2(new_n746), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n761), .B(new_n767), .C1(new_n769), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n617), .A2(new_n662), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n737), .A2(new_n738), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n730), .A2(new_n650), .A3(new_n731), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT48), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n763), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n581), .A2(new_n606), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n585), .A2(new_n781), .A3(new_n317), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n585), .A2(new_n781), .A3(new_n784), .A4(new_n317), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n480), .A2(new_n783), .A3(new_n600), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n480), .A2(new_n608), .A3(new_n515), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n633), .A2(new_n745), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n687), .B1(new_n678), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n641), .A2(new_n652), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n270), .A2(new_n581), .A3(new_n317), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n774), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n406), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n577), .A3(new_n794), .A4(new_n280), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n554), .A3(new_n644), .A4(new_n601), .ZN(new_n796));
  INV_X1    g610(.A(new_n659), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n791), .A3(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n571), .B(new_n312), .C1(new_n270), .C2(new_n317), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n510), .A2(new_n597), .A3(new_n607), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n627), .A2(new_n800), .A3(new_n553), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n675), .A2(new_n611), .A3(new_n634), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n608), .A2(new_n610), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n646), .A2(new_n808), .B1(new_n670), .B2(new_n674), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT111), .A3(new_n634), .A4(new_n802), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n803), .A2(new_n804), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n799), .B1(new_n807), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n813), .B1(new_n811), .B2(new_n803), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n790), .A2(new_n791), .A3(new_n798), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n814), .B2(KEYINPUT53), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n811), .B1(new_n810), .B2(new_n812), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(KEYINPUT112), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n817), .A2(KEYINPUT53), .A3(new_n818), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n780), .B1(new_n820), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n820), .A2(new_n780), .A3(new_n830), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n777), .B(new_n779), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OR2_X1    g647(.A1(G952), .A2(G953), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n515), .B(new_n552), .C1(new_n725), .C2(KEYINPUT49), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n836), .B(new_n695), .C1(KEYINPUT49), .C2(new_n725), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n404), .A3(new_n628), .A4(new_n630), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n835), .A2(new_n838), .ZN(G75));
  NAND3_X1  g653(.A1(new_n822), .A2(new_n829), .A3(new_n827), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(G902), .A3(new_n398), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n351), .A2(new_n376), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(new_n374), .Z(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n194), .A2(G952), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n847), .A2(KEYINPUT120), .A3(new_n849), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(G51));
  NAND2_X1  g670(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n830), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n840), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n543), .B(KEYINPUT57), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n862), .B1(new_n541), .B2(new_n536), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n840), .A2(G902), .A3(new_n705), .A4(new_n707), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n848), .B1(new_n863), .B2(new_n864), .ZN(G54));
  NAND4_X1  g679(.A1(new_n840), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n255), .A2(new_n257), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n868), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n869), .A2(new_n870), .A3(new_n848), .ZN(G60));
  NAND2_X1  g685(.A1(new_n565), .A2(new_n566), .ZN(new_n872));
  NAND2_X1  g686(.A1(G478), .A2(G902), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT59), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n859), .A2(new_n872), .A3(new_n860), .A4(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n832), .A2(new_n831), .A3(new_n874), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n849), .B(new_n876), .C1(new_n877), .C2(new_n872), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(G63));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n880));
  NAND2_X1  g694(.A1(G217), .A2(G902), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT60), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n595), .A2(new_n596), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT122), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n840), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n849), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n511), .B1(new_n840), .B2(new_n882), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n880), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n849), .B(new_n885), .C1(new_n887), .C2(new_n889), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT124), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n840), .A2(new_n882), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n895), .B2(new_n505), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n886), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n888), .B1(new_n893), .B2(new_n898), .ZN(G66));
  INV_X1    g713(.A(G224), .ZN(new_n900));
  OAI21_X1  g714(.A(G953), .B1(new_n278), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n798), .A2(new_n791), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n903), .B2(new_n273), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n844), .B1(G898), .B2(new_n194), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(G69));
  NAND2_X1  g720(.A1(new_n429), .A2(new_n433), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n249), .ZN(new_n908));
  INV_X1    g722(.A(G227), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n273), .A2(G900), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n637), .A2(new_n614), .A3(new_n678), .ZN(new_n911));
  INV_X1    g725(.A(new_n793), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT126), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n911), .A2(KEYINPUT126), .A3(new_n912), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n715), .A2(new_n194), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n809), .A2(new_n634), .ZN(new_n917));
  OR4_X1    g731(.A1(new_n916), .A2(new_n631), .A3(new_n917), .A4(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n631), .A2(new_n917), .B1(new_n916), .B2(KEYINPUT62), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n723), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  OAI221_X1 g735(.A(new_n908), .B1(new_n909), .B2(new_n910), .C1(new_n915), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n701), .A2(new_n714), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n762), .A2(new_n800), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n712), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n723), .A2(new_n634), .A3(new_n689), .A4(new_n809), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n687), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n273), .ZN(new_n928));
  INV_X1    g742(.A(new_n908), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(G227), .B2(new_n910), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n922), .B1(new_n928), .B2(new_n930), .ZN(G72));
  NOR4_X1   g745(.A1(new_n925), .A2(new_n926), .A3(new_n687), .A4(new_n902), .ZN(new_n932));
  NAND2_X1  g746(.A1(G472), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT63), .Z(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n451), .B(new_n622), .C1(new_n932), .C2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n816), .B2(new_n819), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n472), .B2(new_n441), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT127), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n715), .A2(new_n903), .A3(new_n913), .A4(new_n914), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n940), .B2(new_n921), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n848), .B1(new_n941), .B2(new_n623), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n936), .A2(new_n939), .A3(new_n942), .ZN(G57));
endmodule


