//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT91), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n203), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G57gat), .A2(G64gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(new_n205), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT92), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n215), .A3(new_n210), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n214), .A2(new_n202), .A3(new_n208), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G231gat), .A2(G233gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G127gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(KEYINPUT16), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n224), .A2(new_n225), .ZN(new_n228));
  OAI211_X1 g027(.A(KEYINPUT88), .B(G8gat), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n231));
  OR2_X1    g030(.A1(KEYINPUT88), .A2(G8gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(new_n226), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n229), .A2(KEYINPUT89), .A3(new_n233), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n236), .B(new_n237), .C1(new_n219), .C2(new_n218), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n223), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n240));
  INV_X1    g039(.A(G155gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G183gat), .B(G211gat), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n239), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(G232gat), .A2(G233gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT41), .ZN(new_n248));
  XNOR2_X1  g047(.A(G134gat), .B(G162gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G29gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT14), .B(G29gat), .Z(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(G36gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G43gat), .B(G50gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT87), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT15), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n259), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n259), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n255), .A2(new_n264), .B1(new_n258), .B2(new_n261), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G85gat), .ZN(new_n268));
  INV_X1    g067(.A(G92gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(KEYINPUT8), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT7), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(new_n268), .B2(new_n269), .ZN(new_n272));
  NAND3_X1  g071(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G99gat), .B(G106gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n270), .A2(new_n275), .A3(new_n272), .A4(new_n273), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT95), .A3(new_n278), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n278), .A2(KEYINPUT95), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n266), .A2(new_n281), .B1(KEYINPUT41), .B2(new_n247), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT17), .B1(new_n263), .B2(new_n265), .ZN(new_n283));
  INV_X1    g082(.A(new_n281), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n255), .A2(new_n264), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n258), .A2(new_n261), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(new_n288), .A3(new_n262), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n283), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G190gat), .B(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT96), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n251), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(new_n293), .B(new_n250), .C1(new_n282), .C2(new_n290), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(KEYINPUT96), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OR3_X1    g099(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(new_n295), .B2(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n277), .A2(new_n278), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n218), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n281), .A2(new_n218), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT10), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n212), .A4(new_n217), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT97), .ZN(new_n313));
  INV_X1    g112(.A(new_n305), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g117(.A(KEYINPUT10), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n218), .A2(new_n306), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n279), .A2(new_n280), .B1(new_n212), .B2(new_n217), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n314), .B1(new_n322), .B2(new_n310), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT97), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n313), .A2(new_n315), .A3(new_n318), .A4(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n318), .B1(new_n312), .B2(new_n315), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n246), .A2(new_n304), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G169gat), .A2(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  NAND2_X1  g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(G190gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n339), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n336), .B(new_n343), .C1(new_n344), .C2(KEYINPUT25), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n332), .A2(new_n344), .A3(new_n335), .A4(new_n333), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n337), .A2(G190gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n341), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n331), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT65), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n333), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n355), .B2(new_n331), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT27), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G183gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(new_n339), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n367), .A2(new_n368), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n361), .B(new_n362), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  INV_X1    g172(.A(G233gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  INV_X1    g181(.A(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n381), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n380), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(KEYINPUT68), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT69), .B(KEYINPUT29), .Z(new_n394));
  AOI21_X1  g193(.A(new_n375), .B1(new_n372), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n377), .B2(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(G8gat), .B(G36gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT70), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n392), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n380), .A2(new_n391), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n377), .A2(new_n395), .A3(new_n393), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT37), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT38), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n396), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n400), .B1(new_n408), .B2(KEYINPUT37), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n402), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n393), .ZN(new_n411));
  INV_X1    g210(.A(new_n395), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n376), .ZN(new_n413));
  INV_X1    g212(.A(new_n391), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n377), .A2(new_n379), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n400), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT37), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(new_n401), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(KEYINPUT37), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n406), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G141gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT72), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT72), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(G141gat), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n430), .A3(G148gat), .ZN(new_n431));
  INV_X1    g230(.A(G148gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G141gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(KEYINPUT73), .A3(new_n433), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT75), .B(G155gat), .Z(new_n438));
  AND2_X1   g237(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT2), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n241), .A2(G162gat), .ZN(new_n443));
  INV_X1    g242(.A(G162gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(G155gat), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT74), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(G155gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n241), .A2(G162gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n437), .A3(new_n442), .A4(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G127gat), .B(G134gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G113gat), .B(G120gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(KEYINPUT1), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n455), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT1), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n453), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT71), .B(KEYINPUT2), .Z(new_n461));
  XNOR2_X1  g260(.A(G141gat), .B(G148gat), .ZN(new_n462));
  OAI22_X1  g261(.A1(new_n461), .A2(new_n462), .B1(new_n443), .B2(new_n445), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n452), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT4), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n460), .A3(KEYINPUT78), .A4(new_n463), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g270(.A(new_n460), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n473), .A3(new_n463), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n464), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g275(.A1(G225gat), .A2(G233gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT77), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AND4_X1   g278(.A1(new_n469), .A2(new_n475), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n472), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n468), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n478), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT5), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT79), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT5), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n480), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n475), .A2(new_n479), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n467), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n466), .A2(new_n468), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n426), .B1(new_n488), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n469), .A3(new_n476), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n486), .B1(new_n483), .B2(KEYINPUT5), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT79), .B(new_n494), .C1(new_n482), .C2(new_n478), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n425), .A3(new_n495), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n425), .B1(new_n503), .B2(new_n495), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n498), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n421), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n479), .B1(new_n493), .B2(new_n475), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n466), .A2(new_n481), .A3(new_n468), .A4(new_n479), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n511), .A2(KEYINPUT84), .A3(KEYINPUT39), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT84), .B1(new_n511), .B2(KEYINPUT39), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n510), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(new_n475), .A3(new_n490), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT39), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n478), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n425), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n509), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n416), .A2(new_n402), .A3(KEYINPUT30), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n392), .A2(new_n523), .A3(new_n396), .A4(new_n401), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n506), .A2(new_n525), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n514), .A2(new_n519), .A3(new_n509), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n509), .C1(new_n514), .C2(new_n519), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n521), .A2(new_n526), .A3(new_n527), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G228gat), .A2(G233gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n473), .B1(new_n414), .B2(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n470), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n474), .A2(new_n394), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n411), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n531), .B(KEYINPUT81), .Z(new_n536));
  AOI21_X1  g335(.A(new_n391), .B1(new_n474), .B2(new_n394), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT3), .B1(new_n391), .B2(new_n394), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n463), .B2(new_n452), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G78gat), .B(G106gat), .Z(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G50gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(G22gat), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n541), .B2(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(G22gat), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n535), .A2(new_n540), .A3(KEYINPUT82), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n542), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT83), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n554), .A2(new_n555), .A3(new_n546), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n554), .B2(new_n546), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n508), .A2(new_n530), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n546), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT83), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n555), .A3(new_n546), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n548), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI211_X1 g362(.A(new_n425), .B(new_n499), .C1(new_n503), .C2(new_n495), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n506), .A2(new_n498), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(new_n504), .ZN(new_n566));
  INV_X1    g365(.A(new_n525), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G227gat), .A2(G233gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n372), .A2(new_n472), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n353), .A2(new_n371), .A3(new_n460), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT66), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G15gat), .B(G43gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G99gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n569), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n353), .A2(new_n460), .A3(new_n371), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n460), .B1(new_n353), .B2(new_n371), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n577), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT66), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT32), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n574), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT34), .B1(new_n587), .B2(new_n578), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT34), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n589), .A3(new_n569), .A4(new_n571), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(new_n581), .B(KEYINPUT32), .C1(new_n582), .C2(new_n577), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n586), .B2(new_n592), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT67), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT67), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n596), .B1(new_n601), .B2(new_n595), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n559), .A2(new_n568), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT35), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n593), .A2(new_n594), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n561), .A2(new_n562), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n608), .B2(new_n549), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n567), .B1(new_n505), .B2(new_n507), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n505), .A2(new_n507), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n597), .A2(new_n605), .A3(new_n600), .ZN(new_n613));
  AND4_X1   g412(.A1(new_n612), .A2(new_n613), .A3(new_n558), .A4(new_n525), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n229), .A2(KEYINPUT89), .A3(new_n233), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT89), .B1(new_n229), .B2(new_n233), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n266), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n283), .A2(new_n289), .A3(new_n234), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT18), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n287), .A2(new_n262), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n236), .A2(new_n624), .A3(new_n237), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n620), .B(KEYINPUT13), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n618), .A2(new_n619), .A3(KEYINPUT18), .A4(new_n620), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT86), .B(G197gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(KEYINPUT11), .B(G169gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n623), .A2(new_n628), .A3(new_n629), .A4(new_n636), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n615), .A2(KEYINPUT90), .A3(new_n640), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n330), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n566), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT98), .B(G1gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n567), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G8gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(KEYINPUT42), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(G8gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(KEYINPUT42), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(G1325gat));
  NAND2_X1  g455(.A1(new_n643), .A2(new_n644), .ZN(new_n657));
  INV_X1    g456(.A(new_n330), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n659), .B2(new_n603), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n601), .A2(G15gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n563), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n245), .A2(new_n329), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n304), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT101), .Z(new_n673));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n252), .A3(new_n566), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT45), .Z(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n640), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n638), .A2(KEYINPUT102), .A3(new_n639), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n304), .A2(KEYINPUT44), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n611), .A2(new_n614), .A3(KEYINPUT104), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n503), .A2(new_n425), .A3(new_n495), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n506), .A3(new_n498), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n525), .B1(new_n686), .B2(new_n564), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n558), .A2(new_n606), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT35), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n610), .A2(new_n558), .A3(new_n613), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n604), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n602), .B1(new_n687), .B2(new_n563), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(KEYINPUT103), .A3(new_n559), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n682), .B1(new_n692), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n699), .B1(new_n615), .B2(new_n303), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n681), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n252), .B1(new_n702), .B2(new_n566), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n675), .A2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n567), .ZN(new_n705));
  INV_X1    g504(.A(new_n682), .ZN(new_n706));
  AND4_X1   g505(.A1(KEYINPUT103), .A2(new_n559), .A3(new_n603), .A4(new_n568), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT103), .B1(new_n695), .B2(new_n559), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT104), .B1(new_n611), .B2(new_n614), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n684), .A3(new_n690), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n706), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n567), .B(new_n680), .C1(new_n713), .C2(new_n700), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n705), .A2(new_n716), .A3(G36gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n525), .A2(G36gat), .ZN(new_n718));
  INV_X1    g517(.A(new_n644), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT90), .B1(new_n615), .B2(new_n640), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n673), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n657), .A2(new_n673), .A3(new_n724), .A4(new_n718), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n717), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  NAND2_X1  g530(.A1(new_n657), .A2(new_n673), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(G43gat), .A3(new_n601), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n602), .B(new_n680), .C1(new_n713), .C2(new_n700), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G43gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(KEYINPUT47), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n735), .A2(new_n740), .A3(G43gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n735), .B2(G43gat), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n741), .A2(new_n733), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n743), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g543(.A(new_n563), .B(new_n680), .C1(new_n713), .C2(new_n700), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT110), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n698), .A2(new_n701), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n563), .A4(new_n680), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(new_n749), .A3(G50gat), .ZN(new_n750));
  INV_X1    g549(.A(G50gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n563), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n657), .A2(new_n673), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n745), .A2(G50gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n754), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n757), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n751), .B1(new_n745), .B2(KEYINPUT110), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n755), .B1(new_n764), .B2(new_n749), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT48), .B1(new_n758), .B2(new_n754), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT111), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(G1331gat));
  NAND2_X1  g567(.A1(new_n709), .A2(new_n712), .ZN(new_n769));
  INV_X1    g568(.A(new_n679), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n770), .A2(new_n245), .A3(new_n303), .A4(new_n329), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n612), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(G57gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1332gat));
  INV_X1    g574(.A(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777));
  INV_X1    g576(.A(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n567), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT113), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n778), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1333gat));
  XOR2_X1   g582(.A(new_n601), .B(KEYINPUT114), .Z(new_n784));
  AOI21_X1  g583(.A(G71gat), .B1(new_n776), .B2(new_n784), .ZN(new_n785));
  AND4_X1   g584(.A1(G71gat), .A2(new_n769), .A3(new_n602), .A4(new_n771), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n558), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT115), .B(G78gat), .Z(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1335gat));
  NOR3_X1   g590(.A1(new_n246), .A2(new_n304), .A3(new_n770), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n692), .B2(new_n697), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n329), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n268), .A3(new_n566), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n246), .A2(new_n329), .A3(new_n770), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n747), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n566), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n268), .B2(new_n799), .ZN(G1336gat));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT118), .B1(new_n793), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT117), .B1(new_n805), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n793), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n329), .A2(G92gat), .A3(new_n525), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n747), .A2(new_n567), .A3(new_n797), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(KEYINPUT116), .A3(G92gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT116), .B1(new_n810), .B2(G92gat), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(G92gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  INV_X1    g615(.A(new_n808), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n815), .B(new_n816), .C1(new_n794), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(G1337gat));
  INV_X1    g618(.A(G99gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n601), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n795), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n798), .A2(new_n602), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n820), .B2(new_n823), .ZN(G1338gat));
  NAND3_X1  g623(.A1(new_n747), .A2(new_n563), .A3(new_n797), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  OR3_X1    g626(.A1(new_n558), .A2(new_n329), .A3(G106gat), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n826), .B(new_n827), .C1(new_n794), .C2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n828), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n804), .A2(new_n807), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n826), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n829), .B1(new_n832), .B2(new_n827), .ZN(G1339gat));
  NAND4_X1  g632(.A1(new_n246), .A2(new_n304), .A3(new_n329), .A4(new_n679), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n318), .B1(new_n323), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n313), .A2(KEYINPUT54), .A3(new_n325), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n322), .A2(new_n314), .A3(new_n310), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT119), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n836), .B(KEYINPUT55), .C1(new_n837), .C2(new_n839), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n326), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n626), .A2(new_n627), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n620), .B1(new_n618), .B2(new_n619), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n635), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n303), .A2(new_n639), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n639), .B(new_n847), .C1(new_n327), .C2(new_n328), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n844), .B2(new_n679), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n851), .B2(new_n304), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n834), .B1(new_n852), .B2(new_n246), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n566), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n854), .A2(new_n525), .A3(new_n609), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n770), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n853), .A2(new_n558), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(new_n566), .A3(new_n525), .A4(new_n821), .ZN(new_n858));
  INV_X1    g657(.A(G113gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n640), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n856), .A2(new_n861), .ZN(G1340gat));
  INV_X1    g661(.A(new_n329), .ZN(new_n863));
  AOI21_X1  g662(.A(G120gat), .B1(new_n855), .B2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(G120gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n858), .A2(new_n865), .A3(new_n329), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(G1341gat));
  INV_X1    g666(.A(G127gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n855), .A2(new_n868), .A3(new_n246), .ZN(new_n869));
  OAI21_X1  g668(.A(G127gat), .B1(new_n858), .B2(new_n245), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT120), .Z(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n873), .A3(new_n303), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n858), .B2(new_n304), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n428), .A2(new_n430), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n602), .A2(new_n612), .A3(new_n567), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n853), .B2(new_n563), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n563), .A2(KEYINPUT57), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n842), .A2(new_n326), .A3(new_n640), .A4(new_n843), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n303), .B1(new_n884), .B2(new_n850), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n245), .B1(new_n885), .B2(new_n849), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n886), .B2(new_n834), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n881), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n879), .B(new_n880), .C1(new_n888), .C2(new_n860), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n602), .A2(new_n558), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n854), .A2(new_n525), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n427), .A3(new_n640), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n889), .B(new_n892), .C1(KEYINPUT122), .C2(new_n879), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT122), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n888), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT121), .B(new_n881), .C1(new_n882), .C2(new_n887), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n770), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(new_n880), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n893), .B1(new_n900), .B2(new_n879), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n891), .A2(new_n863), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(KEYINPUT59), .A3(new_n432), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n881), .A2(KEYINPUT59), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n853), .A2(KEYINPUT57), .A3(new_n563), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n886), .B1(new_n640), .B2(new_n330), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n563), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n863), .B(new_n904), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n863), .A3(new_n897), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n912), .B2(new_n432), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT123), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n915), .B(new_n903), .C1(new_n912), .C2(new_n432), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1345gat));
  NAND3_X1  g716(.A1(new_n891), .A2(new_n438), .A3(new_n246), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n898), .A2(new_n246), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n438), .ZN(G1346gat));
  NAND3_X1  g719(.A1(new_n891), .A2(new_n441), .A3(new_n303), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n898), .A2(new_n303), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n922), .A2(KEYINPUT124), .B1(new_n440), .B2(new_n439), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n922), .A2(KEYINPUT124), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(G1347gat));
  AND2_X1   g724(.A1(new_n853), .A2(new_n612), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(new_n567), .A3(new_n609), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n770), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n857), .A2(new_n612), .A3(new_n567), .A4(new_n784), .ZN(new_n929));
  INV_X1    g728(.A(G169gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n929), .A2(new_n930), .A3(new_n860), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n928), .A2(new_n931), .ZN(G1348gat));
  INV_X1    g731(.A(G176gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n933), .A3(new_n863), .ZN(new_n934));
  OAI21_X1  g733(.A(G176gat), .B1(new_n929), .B2(new_n329), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1349gat));
  NAND4_X1  g735(.A1(new_n927), .A2(new_n364), .A3(new_n366), .A4(new_n246), .ZN(new_n937));
  OAI21_X1  g736(.A(G183gat), .B1(new_n929), .B2(new_n245), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n929), .B2(new_n304), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n339), .A3(new_n303), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1351gat));
  AND3_X1   g743(.A1(new_n926), .A2(new_n567), .A3(new_n890), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n770), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n905), .A2(new_n907), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n602), .A2(new_n566), .A3(new_n525), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT125), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT126), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n640), .A2(G197gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n946), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  INV_X1    g753(.A(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n945), .A2(new_n955), .A3(new_n863), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT62), .Z(new_n957));
  NAND2_X1  g756(.A1(new_n947), .A2(new_n863), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n958), .B2(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(G1353gat));
  OR2_X1    g759(.A1(new_n950), .A2(new_n245), .ZN(new_n961));
  OAI21_X1  g760(.A(G211gat), .B1(new_n948), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g761(.A1(new_n962), .A2(KEYINPUT63), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(KEYINPUT63), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n383), .A3(new_n246), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n945), .B2(new_n303), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n304), .A2(new_n384), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n952), .B2(new_n969), .ZN(G1355gat));
endmodule


