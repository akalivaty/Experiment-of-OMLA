//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g002(.A(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n208), .A2(KEYINPUT77), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(new_n208), .B2(KEYINPUT77), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT22), .ZN(new_n213));
  INV_X1    g012(.A(G211gat), .ZN(new_n214));
  INV_X1    g013(.A(G218gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT74), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n219));
  XNOR2_X1  g018(.A(G197gat), .B(G204gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G211gat), .B(G218gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n217), .A2(new_n222), .A3(new_n219), .A4(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT29), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n212), .B1(new_n226), .B2(KEYINPUT3), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n210), .B2(new_n211), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n225), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G228gat), .ZN(new_n235));
  INV_X1    g034(.A(G233gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n227), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n230), .B1(new_n225), .B2(KEYINPUT82), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n224), .A2(KEYINPUT82), .A3(new_n225), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n208), .A2(KEYINPUT77), .ZN(new_n244));
  INV_X1    g043(.A(new_n209), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n208), .A2(KEYINPUT77), .A3(new_n209), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n234), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n238), .B1(new_n239), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT83), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n253));
  INV_X1    g052(.A(G50gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G78gat), .ZN(new_n256));
  INV_X1    g055(.A(G106gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n227), .A2(new_n234), .A3(new_n237), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n232), .B1(new_n230), .B2(new_n229), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n224), .A2(KEYINPUT82), .A3(new_n225), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n228), .B1(new_n261), .B2(new_n240), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n262), .B2(new_n212), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n251), .B(new_n259), .C1(new_n263), .C2(new_n237), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n259), .B1(new_n263), .B2(new_n237), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G22gat), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n252), .A2(new_n258), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT83), .ZN(new_n268));
  AND4_X1   g067(.A1(new_n268), .A2(new_n266), .A3(new_n264), .A4(new_n258), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT40), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT39), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273));
  XNOR2_X1  g072(.A(G127gat), .B(G134gat), .ZN(new_n274));
  INV_X1    g073(.A(G113gat), .ZN(new_n275));
  OR2_X1    g074(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT69), .A2(G120gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n275), .A2(G120gat), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n273), .B(new_n274), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n274), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G120gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n281), .B1(KEYINPUT1), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n248), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n283), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n212), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n284), .B2(new_n248), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n212), .A2(new_n286), .A3(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n246), .A2(KEYINPUT3), .A3(new_n247), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n229), .A2(new_n298), .A3(new_n286), .ZN(new_n299));
  INV_X1    g098(.A(new_n295), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n248), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n212), .A2(new_n286), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n301), .B(KEYINPUT79), .C1(new_n302), .C2(new_n293), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n297), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  AOI211_X1 g103(.A(new_n272), .B(new_n291), .C1(new_n304), .C2(new_n290), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n272), .A3(new_n290), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  INV_X1    g106(.A(G85gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT0), .B(G57gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n271), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n297), .A2(new_n303), .A3(new_n315), .A4(new_n299), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n302), .B1(new_n299), .B2(new_n295), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n285), .A2(new_n293), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n317), .A2(new_n290), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n288), .A2(new_n290), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n316), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n290), .ZN(new_n324));
  INV_X1    g123(.A(new_n291), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(KEYINPUT39), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n326), .A2(KEYINPUT40), .A3(new_n312), .A4(new_n306), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n314), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT30), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  OR2_X1    g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n332), .A2(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(G176gat), .ZN(new_n339));
  AND2_X1   g138(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT65), .B(G169gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n345), .A2(KEYINPUT66), .A3(new_n339), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n333), .A2(KEYINPUT67), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n354), .B2(new_n332), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n334), .A2(new_n338), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n334), .B2(new_n336), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n361));
  INV_X1    g160(.A(G183gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(KEYINPUT27), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT27), .B(G183gat), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n360), .B(new_n363), .C1(new_n364), .C2(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(KEYINPUT28), .A3(new_n360), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n334), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT26), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT26), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n335), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n371), .B(new_n331), .C1(new_n373), .C2(new_n370), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n359), .A2(new_n376), .B1(new_n230), .B2(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n347), .A2(new_n348), .B1(new_n355), .B2(new_n357), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n367), .B2(new_n368), .ZN(new_n380));
  INV_X1    g179(.A(new_n377), .ZN(new_n381));
  NOR3_X1   g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n233), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n359), .A2(new_n376), .A3(new_n377), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n379), .A2(new_n380), .B1(KEYINPUT29), .B2(new_n381), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n232), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT75), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n233), .C1(new_n378), .C2(new_n382), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT76), .B(new_n329), .C1(new_n390), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n393), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n387), .B2(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT30), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n270), .B1(new_n328), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT80), .B1(new_n323), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n322), .A2(new_n403), .A3(KEYINPUT6), .A4(new_n311), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n316), .B(new_n312), .C1(new_n319), .C2(new_n321), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n323), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n389), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT37), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n387), .A2(KEYINPUT37), .A3(new_n389), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n393), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n396), .B1(new_n412), .B2(KEYINPUT38), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n383), .A2(new_n386), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT38), .B1(new_n414), .B2(KEYINPUT37), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n393), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n407), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n404), .A3(new_n406), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n418), .A2(new_n395), .A3(new_n398), .A4(new_n394), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n400), .A2(new_n417), .B1(new_n419), .B2(new_n270), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT36), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n359), .A2(new_n376), .A3(new_n284), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT70), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT70), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n359), .A2(new_n376), .A3(new_n424), .A4(new_n284), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n286), .B1(new_n379), .B2(new_n380), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT71), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT71), .B(new_n286), .C1(new_n379), .C2(new_n380), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n423), .A2(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT34), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n425), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT34), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .A4(new_n431), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n430), .A2(new_n439), .A3(new_n436), .A4(new_n431), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n433), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  AOI21_X1  g243(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(KEYINPUT33), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT32), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450));
  INV_X1    g249(.A(new_n444), .ZN(new_n451));
  OAI221_X1 g250(.A(KEYINPUT32), .B1(new_n450), .B2(new_n451), .C1(new_n430), .C2(new_n431), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n441), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n438), .A2(new_n440), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT32), .B1(new_n430), .B2(new_n431), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n430), .B2(new_n431), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n444), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n455), .A2(new_n458), .A3(new_n452), .A4(new_n433), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n421), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n459), .A3(KEYINPUT73), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n455), .A2(new_n433), .B1(new_n458), .B2(new_n452), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT73), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n460), .B1(new_n465), .B2(new_n421), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n267), .A2(new_n269), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n407), .A2(new_n399), .A3(KEYINPUT35), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n459), .A3(new_n454), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n470), .B2(new_n419), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n420), .A2(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT16), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(G1gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G22gat), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n477), .B(KEYINPUT87), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n482), .C1(G1gat), .C2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(G1gat), .ZN(new_n485));
  OAI21_X1  g284(.A(G8gat), .B1(new_n485), .B2(new_n480), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT88), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(KEYINPUT90), .B(G57gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G64gat), .ZN(new_n494));
  INV_X1    g293(.A(G64gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G57gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500));
  INV_X1    g299(.A(new_n492), .ZN(new_n501));
  XNOR2_X1  g300(.A(G57gat), .B(G64gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n362), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n362), .B1(new_n491), .B2(new_n508), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n474), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n508), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G183gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n509), .A3(new_n473), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G211gat), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n512), .B2(new_n515), .ZN(new_n519));
  XNOR2_X1  g318(.A(G127gat), .B(G155gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OR3_X1    g322(.A1(new_n518), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT93), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(G85gat), .A3(G92gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(G92gat), .ZN(new_n533));
  AOI22_X1  g332(.A1(KEYINPUT8), .A2(new_n532), .B1(new_n308), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n528), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G99gat), .B(G106gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n531), .A2(new_n534), .A3(new_n537), .A4(new_n535), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n254), .A2(G43gat), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT15), .B1(new_n543), .B2(KEYINPUT85), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  OR3_X1    g345(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n547), .A2(new_n548), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT84), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n549), .A2(new_n552), .A3(new_n551), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n550), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G232gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n236), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n542), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT86), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n559), .A3(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT17), .B1(new_n555), .B2(new_n559), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n558), .B1(new_n563), .B2(new_n542), .ZN(new_n564));
  XNOR2_X1  g363(.A(G190gat), .B(G218gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT95), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n558), .B(new_n566), .C1(new_n563), .C2(new_n542), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n571), .B(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n472), .A2(new_n527), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n486), .B(new_n484), .C1(new_n561), .C2(new_n562), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n489), .A2(new_n555), .A3(new_n490), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n555), .ZN(new_n585));
  INV_X1    g384(.A(new_n490), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT88), .B1(new_n484), .B2(new_n486), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n580), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n582), .B(KEYINPUT13), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT18), .A4(new_n582), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n584), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  INV_X1    g394(.A(G197gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT11), .B(G169gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT12), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n584), .A2(new_n592), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n500), .B1(new_n497), .B2(KEYINPUT91), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n504), .A2(new_n500), .A3(new_n501), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(new_n499), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n542), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n538), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n507), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT10), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n542), .A2(new_n507), .A3(KEYINPUT10), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G230gat), .ZN(new_n615));
  OAI22_X1  g414(.A1(new_n612), .A2(new_n614), .B1(new_n615), .B2(new_n236), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n608), .A2(new_n538), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n608), .B2(new_n542), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n615), .A2(new_n236), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n605), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n577), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n418), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT97), .B(G1gat), .Z(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1324gat));
  INV_X1    g431(.A(new_n399), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(G8gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT16), .B(G8gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT98), .ZN(new_n637));
  NOR2_X1   g436(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  AOI22_X1  g438(.A1(new_n635), .A2(KEYINPUT42), .B1(new_n634), .B2(new_n639), .ZN(G1325gat));
  INV_X1    g439(.A(new_n629), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT36), .B1(new_n461), .B2(new_n464), .ZN(new_n642));
  OAI21_X1  g441(.A(KEYINPUT100), .B1(new_n642), .B2(new_n460), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n642), .A2(KEYINPUT100), .A3(new_n460), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n641), .A2(G15gat), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(G15gat), .B1(new_n641), .B2(new_n465), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(G1326gat));
  OR3_X1    g448(.A1(new_n629), .A2(KEYINPUT101), .A3(new_n467), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT101), .B1(new_n629), .B2(new_n467), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT43), .B(G22gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  INV_X1    g453(.A(G29gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n527), .A2(new_n628), .ZN(new_n656));
  INV_X1    g455(.A(new_n576), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT44), .B1(new_n472), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n465), .A2(new_n421), .ZN(new_n659));
  INV_X1    g458(.A(new_n460), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n420), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n469), .A2(new_n471), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n576), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n656), .B1(new_n658), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n655), .B1(new_n666), .B2(new_n407), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n472), .A2(new_n657), .A3(new_n656), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n655), .A3(new_n407), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT45), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT45), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n671), .A3(new_n655), .A4(new_n407), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT102), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675));
  INV_X1    g474(.A(G36gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n668), .A2(new_n676), .A3(new_n399), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n668), .A2(new_n679), .A3(new_n676), .A4(new_n399), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n675), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n675), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n399), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G36gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .A4(new_n686), .ZN(G1329gat));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  INV_X1    g487(.A(new_n466), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n526), .A2(new_n605), .A3(new_n627), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n664), .B1(new_n663), .B2(new_n576), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT44), .B(new_n657), .C1(new_n661), .C2(new_n662), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G43gat), .ZN(new_n694));
  INV_X1    g493(.A(G43gat), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n663), .A2(new_n695), .A3(new_n576), .A4(new_n690), .ZN(new_n696));
  INV_X1    g495(.A(new_n465), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n688), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n688), .B1(new_n696), .B2(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n666), .A2(new_n646), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(G43gat), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n700), .A2(KEYINPUT105), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n695), .B1(new_n666), .B2(new_n689), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT47), .B1(new_n706), .B2(new_n698), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n466), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n643), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n710), .B(new_n656), .C1(new_n658), .C2(new_n665), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n688), .B(new_n699), .C1(new_n711), .C2(new_n695), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n705), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n704), .A2(new_n713), .ZN(G1330gat));
  OAI211_X1 g513(.A(new_n270), .B(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n663), .A2(new_n254), .A3(new_n576), .A4(new_n690), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n716), .B(KEYINPUT48), .C1(new_n467), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n467), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n668), .A2(KEYINPUT106), .A3(new_n254), .A4(new_n270), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n716), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n254), .B1(new_n666), .B2(new_n270), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n721), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n719), .B(new_n724), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n718), .B1(new_n725), .B2(new_n729), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n527), .A2(new_n576), .ZN(new_n731));
  INV_X1    g530(.A(new_n627), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n604), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n663), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n663), .A2(new_n731), .A3(KEYINPUT108), .A4(new_n733), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n407), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(new_n493), .Z(G1332gat));
  NAND2_X1  g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n399), .B(KEYINPUT109), .Z(new_n742));
  NAND4_X1  g541(.A1(new_n736), .A2(new_n737), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT110), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(KEYINPUT110), .ZN(new_n745));
  OR2_X1    g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n736), .A2(new_n465), .A3(new_n737), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(G71gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n736), .A2(KEYINPUT111), .A3(new_n465), .A4(new_n737), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n738), .A2(G71gat), .A3(new_n646), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT50), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n738), .A2(new_n270), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n472), .B2(new_n657), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n663), .A2(KEYINPUT112), .A3(new_n576), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n526), .A2(new_n604), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT51), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(new_n308), .A3(new_n407), .A4(new_n627), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n527), .A2(new_n733), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n658), .B2(new_n665), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n418), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n742), .A2(new_n533), .A3(new_n627), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT113), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n742), .ZN(new_n782));
  OAI21_X1  g581(.A(G92gat), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n533), .B1(new_n775), .B2(new_n399), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n772), .B2(new_n780), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n781), .A2(new_n785), .B1(new_n787), .B2(new_n784), .ZN(G1337gat));
  NOR2_X1   g587(.A1(new_n697), .A2(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n627), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(G99gat), .B1(new_n776), .B2(new_n710), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1338gat));
  NAND3_X1  g591(.A1(new_n627), .A2(new_n257), .A3(new_n270), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT114), .Z(new_n794));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n257), .B1(new_n775), .B2(new_n270), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n795), .A2(KEYINPUT115), .A3(KEYINPUT53), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g597(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n799));
  NAND2_X1  g598(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n800));
  INV_X1    g599(.A(new_n794), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n770), .B2(new_n771), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n796), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n798), .A2(new_n803), .ZN(G1339gat));
  OAI211_X1 g603(.A(new_n619), .B(new_n613), .C1(new_n618), .C2(KEYINPUT10), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n616), .A3(KEYINPUT54), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  OAI221_X1 g608(.A(new_n809), .B1(new_n615), .B2(new_n236), .C1(new_n612), .C2(new_n614), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n624), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n805), .A2(new_n616), .A3(KEYINPUT116), .A4(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n808), .A2(new_n811), .A3(KEYINPUT55), .A4(new_n812), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n815), .A2(new_n604), .A3(new_n625), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n588), .A2(new_n580), .A3(new_n590), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT117), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n581), .A2(new_n583), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n588), .A2(new_n580), .A3(new_n821), .A4(new_n590), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n599), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n627), .A2(new_n603), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n576), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(new_n625), .A3(new_n816), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n824), .B2(new_n603), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n828), .A3(new_n603), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n576), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n527), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n526), .A2(new_n605), .A3(new_n732), .A4(new_n657), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n418), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n470), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n782), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n275), .A3(new_n604), .ZN(new_n839));
  AOI211_X1 g638(.A(new_n270), .B(new_n697), .C1(new_n833), .C2(new_n834), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n742), .A2(new_n418), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n605), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n839), .A2(new_n843), .ZN(G1340gat));
  NAND2_X1  g643(.A1(new_n276), .A2(new_n277), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n838), .A2(new_n845), .A3(new_n627), .ZN(new_n846));
  OAI21_X1  g645(.A(G120gat), .B1(new_n842), .B2(new_n732), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n838), .B2(new_n526), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n842), .A2(new_n527), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(G127gat), .B2(new_n850), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n657), .A2(new_n399), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n837), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n842), .B2(new_n657), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n841), .A2(new_n466), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT119), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n833), .A2(new_n834), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT57), .B1(new_n862), .B2(new_n270), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n864), .B(new_n467), .C1(new_n833), .C2(new_n834), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n604), .B(new_n861), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n862), .A2(new_n407), .A3(new_n270), .A4(new_n710), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n742), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n204), .A3(new_n604), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1344gat));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n205), .A3(new_n627), .ZN(new_n876));
  INV_X1    g675(.A(new_n861), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n270), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n864), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n862), .A2(KEYINPUT57), .A3(new_n270), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT59), .B(new_n205), .C1(new_n881), .C2(new_n627), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n627), .A3(new_n861), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n876), .B1(new_n882), .B2(new_n886), .ZN(G1345gat));
  NOR3_X1   g686(.A1(new_n868), .A2(new_n527), .A3(new_n742), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT120), .ZN(new_n889));
  INV_X1    g688(.A(G155gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n527), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n889), .A2(new_n890), .B1(new_n881), .B2(new_n891), .ZN(G1346gat));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n576), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G162gat), .ZN(new_n894));
  INV_X1    g693(.A(G162gat), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n853), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n868), .B2(new_n896), .ZN(G1347gat));
  NAND2_X1  g696(.A1(new_n399), .A2(new_n418), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT121), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n840), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n605), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n407), .B1(new_n833), .B2(new_n834), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n902), .A2(new_n836), .A3(new_n742), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n604), .A3(new_n345), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n903), .B2(new_n627), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n900), .A2(new_n732), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(G176gat), .B2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(G183gat), .B1(new_n900), .B2(new_n527), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n903), .A2(new_n364), .A3(new_n526), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n840), .A2(new_n576), .A3(new_n899), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(G190gat), .ZN(new_n914));
  XOR2_X1   g713(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n915));
  OR2_X1    g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n903), .A2(new_n360), .A3(new_n576), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n915), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(G1351gat));
  OAI211_X1 g718(.A(new_n270), .B(new_n742), .C1(new_n644), .C2(new_n645), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n710), .A2(KEYINPUT123), .A3(new_n270), .A4(new_n742), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n902), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT124), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n922), .A2(new_n902), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n596), .A3(new_n604), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n710), .A2(new_n899), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n884), .A2(new_n604), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n596), .B2(new_n932), .ZN(G1352gat));
  OAI211_X1 g732(.A(new_n627), .B(new_n930), .C1(new_n863), .C2(new_n865), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT125), .B(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n924), .A2(new_n732), .A3(new_n938), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1353gat));
  NAND3_X1  g741(.A1(new_n928), .A2(new_n214), .A3(new_n526), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n526), .B(new_n930), .C1(new_n863), .C2(new_n865), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n944), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1354gat));
  NAND4_X1  g746(.A1(new_n925), .A2(new_n215), .A3(new_n576), .A4(new_n927), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n576), .B(new_n930), .C1(new_n863), .C2(new_n865), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G218gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


