//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1156, new_n1157;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n462), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n465), .A2(new_n467), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(G124), .B1(G136), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n492), .B(new_n461), .C1(new_n465), .C2(new_n467), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n461), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT72), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n461), .C1(new_n503), .C2(new_n472), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT4), .A2(G138), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT3), .B1(new_n466), .B2(G2104), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n461), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g086(.A(G126), .B(G2105), .C1(new_n508), .C2(new_n509), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(new_n500), .ZN(new_n514));
  AND3_X1   g089(.A1(new_n502), .A2(new_n511), .A3(new_n514), .ZN(G164));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT74), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT6), .B(G651), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n518), .A2(new_n520), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n526), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n525), .B(new_n530), .C1(new_n531), .C2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  NAND3_X1  g110(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n536), .B(new_n538), .C1(new_n533), .C2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n526), .A2(G543), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT75), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n540), .B1(G51), .B2(new_n542), .ZN(G168));
  INV_X1    g118(.A(new_n533), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n542), .A2(G52), .B1(G90), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n545), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT77), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT77), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT78), .Z(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT79), .B(G81), .Z(new_n557));
  AOI22_X1  g132(.A1(new_n542), .A2(G43), .B1(new_n544), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT80), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n521), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n544), .A2(G91), .B1(G651), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n541), .B2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n526), .A2(KEYINPUT81), .A3(G53), .A4(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT9), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n572), .B(new_n577), .C1(new_n541), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n571), .A2(new_n576), .A3(new_n578), .ZN(G299));
  AND2_X1   g154(.A1(new_n551), .A2(new_n552), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  NAND2_X1  g156(.A1(new_n544), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n527), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n532), .A2(new_n586), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT83), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT82), .B1(new_n521), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n533), .A2(new_n594), .B1(new_n595), .B2(new_n541), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n542), .A2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n544), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n546), .C2(new_n601), .ZN(G290));
  AOI22_X1  g177(.A1(new_n532), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n546), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n542), .B2(G54), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n532), .A2(G92), .A3(new_n526), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(new_n608), .ZN(new_n616));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n484), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n625));
  INV_X1    g200(.A(G123), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n623), .B1(new_n624), .B2(new_n625), .C1(new_n482), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  AND2_X1   g221(.A1(new_n646), .A2(G14), .ZN(G401));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT85), .Z(new_n649));
  XOR2_X1   g224(.A(G2067), .B(G2678), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  INV_X1    g230(.A(new_n650), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n651), .B1(new_n649), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n653), .B(KEYINPUT17), .Z(new_n659));
  AND2_X1   g234(.A1(new_n649), .A2(new_n650), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT87), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n675), .A2(new_n667), .A3(new_n670), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n676), .C1(new_n667), .C2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  INV_X1    g255(.A(G1981), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n679), .B(new_n682), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT89), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NAND2_X1  g261(.A1(new_n484), .A2(G131), .ZN(new_n687));
  NOR2_X1   g262(.A1(G95), .A2(G2105), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(new_n461), .B2(G107), .ZN(new_n689));
  INV_X1    g264(.A(G119), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n687), .B1(new_n688), .B2(new_n689), .C1(new_n690), .C2(new_n482), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n692), .S(G29), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT35), .B(G1991), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G24), .B(G290), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT93), .B(G1971), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(G6), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n596), .B1(G651), .B2(new_n592), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G16), .B2(G23), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT33), .ZN(new_n713));
  INV_X1    g288(.A(G1976), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(KEYINPUT33), .ZN(new_n717));
  AOI21_X1  g292(.A(G1976), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n703), .B(new_n709), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT34), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n698), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n727), .B(new_n698), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G33), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n484), .A2(G139), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n473), .A2(new_n474), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n734), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT97), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n731), .B(new_n733), .C1(new_n736), .C2(new_n461), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT98), .Z(new_n738));
  AOI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G2072), .Z(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G32), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n481), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G2105), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n483), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n741), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT99), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT27), .B(G1996), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n741), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n741), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT29), .Z(new_n756));
  INV_X1    g331(.A(G2090), .ZN(new_n757));
  OR3_X1    g332(.A1(new_n756), .A2(KEYINPUT103), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(G299), .A2(G16), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G20), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G16), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n759), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G1956), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT103), .B1(new_n756), .B2(new_n757), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n758), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT95), .Z(new_n773));
  AOI22_X1  g348(.A1(new_n483), .A2(G128), .B1(G140), .B2(new_n484), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n741), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n741), .A2(G26), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT28), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT28), .B2(new_n779), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(KEYINPUT24), .A2(G34), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT24), .A2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G160), .B2(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(G2084), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n699), .A2(G21), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G168), .B2(new_n699), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1966), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n627), .A2(new_n741), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT100), .Z(new_n794));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G28), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(G28), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n796), .A2(new_n797), .A3(G29), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n789), .A2(new_n792), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n756), .A2(new_n757), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n770), .A2(new_n783), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G5), .A2(G16), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G171), .B2(G16), .ZN(new_n804));
  MUX2_X1   g379(.A(new_n803), .B(new_n804), .S(KEYINPUT101), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1961), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G19), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n560), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT94), .B(G1341), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n788), .A2(G2084), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n616), .A2(new_n699), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G4), .B2(new_n699), .ZN(new_n814));
  INV_X1    g389(.A(G1348), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n741), .A2(G27), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G164), .B2(new_n741), .ZN(new_n818));
  INV_X1    g393(.A(G2078), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT31), .B(G11), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n814), .A2(new_n815), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n816), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR4_X1   g398(.A1(new_n802), .A2(new_n806), .A3(new_n812), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n729), .A2(new_n740), .A3(new_n753), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(new_n802), .ZN(new_n829));
  INV_X1    g404(.A(new_n812), .ZN(new_n830));
  INV_X1    g405(.A(new_n823), .ZN(new_n831));
  INV_X1    g406(.A(new_n806), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n726), .B2(new_n728), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n834), .A2(new_n826), .A3(new_n740), .A4(new_n753), .ZN(G150));
  AOI22_X1  g410(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  INV_X1    g411(.A(G93), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n836), .A2(new_n546), .B1(new_n837), .B2(new_n533), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G55), .B2(new_n542), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT106), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n559), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n559), .A2(new_n839), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n616), .A2(G559), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT39), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n844), .B1(new_n852), .B2(G860), .ZN(G145));
  NAND2_X1  g428(.A1(new_n506), .A2(new_n510), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n512), .A2(new_n500), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n776), .A2(new_n777), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n857), .B1(new_n776), .B2(new_n777), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n859), .A2(new_n748), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n776), .A2(new_n777), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n856), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n749), .B1(new_n863), .B2(new_n858), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT108), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n748), .B1(new_n859), .B2(new_n860), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT108), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n749), .A3(new_n858), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n738), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n861), .B2(new_n864), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(KEYINPUT109), .A3(new_n868), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n737), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n484), .A2(G142), .ZN(new_n876));
  NOR2_X1   g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n878));
  INV_X1    g453(.A(G130), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n876), .B1(new_n877), .B2(new_n878), .C1(new_n879), .C2(new_n482), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n630), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n691), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT110), .ZN(new_n884));
  INV_X1    g459(.A(new_n882), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n870), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n627), .B(KEYINPUT107), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n479), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G162), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n885), .B1(new_n870), .B2(new_n874), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(KEYINPUT110), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n883), .A2(new_n886), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT111), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G395));
  NAND2_X1  g477(.A1(new_n842), .A2(new_n609), .ZN(new_n903));
  XNOR2_X1  g478(.A(G305), .B(G288), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(G290), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(G166), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n847), .B(new_n619), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n608), .B(G299), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(KEYINPUT41), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(KEYINPUT112), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT112), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n616), .A2(new_n912), .A3(G299), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n914), .B2(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n908), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n907), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n903), .B1(new_n919), .B2(new_n609), .ZN(G295));
  XOR2_X1   g495(.A(G295), .B(KEYINPUT113), .Z(G331));
  INV_X1    g496(.A(new_n909), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(G301), .A2(G168), .ZN(new_n924));
  NAND2_X1  g499(.A1(G171), .A2(G286), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n847), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n924), .A2(new_n846), .A3(new_n845), .A4(new_n925), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT114), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n926), .B2(new_n847), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n928), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n914), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT41), .B(new_n909), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n906), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n915), .B1(new_n927), .B2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n931), .B1(new_n933), .B2(new_n930), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(new_n917), .ZN(new_n940));
  INV_X1    g515(.A(new_n906), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n937), .A2(KEYINPUT43), .A3(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n929), .A2(new_n914), .A3(new_n931), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n906), .B1(new_n944), .B2(new_n938), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT43), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT44), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n937), .A2(new_n948), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n939), .A2(new_n917), .ZN(new_n950));
  INV_X1    g525(.A(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n945), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n958), .ZN(G397));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n854), .B2(new_n855), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n470), .A2(new_n477), .A3(G40), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT46), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n862), .B(new_n782), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n749), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n970), .B2(new_n965), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n748), .B(new_n966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n694), .B(new_n692), .C1(new_n974), .C2(new_n965), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n862), .A2(G2067), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n965), .ZN(new_n978));
  INV_X1    g553(.A(new_n965), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n691), .B(new_n694), .Z(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT126), .Z(new_n982));
  NOR3_X1   g557(.A1(new_n979), .A2(G1986), .A3(G290), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n972), .B(new_n977), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT127), .Z(new_n986));
  INV_X1    g561(.A(KEYINPUT54), .ZN(new_n987));
  INV_X1    g562(.A(new_n963), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT116), .B1(new_n988), .B2(new_n964), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  INV_X1    g565(.A(new_n964), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n963), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n502), .A2(new_n511), .A3(new_n514), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n960), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n989), .B(new_n992), .C1(new_n962), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n996));
  OR3_X1    g571(.A1(new_n995), .A2(new_n996), .A3(G2078), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n995), .B2(G2078), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(KEYINPUT53), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n961), .B2(new_n962), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n994), .B2(new_n962), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n819), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  INV_X1    g578(.A(new_n961), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n964), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n994), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1006), .B1(new_n1007), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(G1961), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1002), .A2(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G301), .B1(new_n999), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(G301), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OR4_X1    g588(.A1(new_n1003), .A2(new_n988), .A3(new_n1000), .A4(G2078), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n987), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G168), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1018), .B2(KEYINPUT121), .ZN(new_n1019));
  INV_X1    g594(.A(G1966), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n995), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1008), .ZN(new_n1022));
  INV_X1    g597(.A(G2084), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(G8), .B(new_n1019), .C1(new_n1025), .C2(G286), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1018), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1019), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n995), .A2(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1027), .B(new_n1028), .C1(new_n1029), .C2(new_n1017), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(G8), .A3(G286), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n705), .A2(new_n681), .ZN(new_n1034));
  NOR2_X1   g609(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n961), .A2(new_n964), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n1017), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1035), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n714), .B2(G288), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(G288), .B2(new_n714), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1038), .B(new_n1043), .C1(new_n714), .C2(G288), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  AND3_X1   g621(.A1(G303), .A2(new_n1046), .A3(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(G303), .B2(G8), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1001), .A2(G1971), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1008), .A2(G2090), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(G8), .C1(new_n1050), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n993), .A2(new_n1005), .A3(new_n960), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n964), .B1(new_n961), .B2(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1001), .A2(G1971), .B1(G2090), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1049), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT123), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1058), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1052), .A4(new_n1045), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n999), .A2(new_n1013), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT124), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1010), .A2(new_n1067), .A3(new_n1014), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(G171), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1069), .A3(KEYINPUT54), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1016), .A2(new_n1032), .A3(new_n1063), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1001), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1056), .B2(new_n765), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT117), .B(G1956), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n570), .A2(G651), .ZN(new_n1079));
  INV_X1    g654(.A(G91), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n578), .B(new_n1079), .C1(new_n1080), .C2(new_n533), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT118), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n571), .A2(new_n576), .A3(new_n1084), .A4(new_n578), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1083), .A2(KEYINPUT57), .A3(new_n1085), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1078), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1090), .B(new_n1074), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT119), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1092), .A2(new_n1096), .A3(new_n1093), .A4(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1001), .A2(new_n966), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT58), .B(G1341), .Z(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n961), .B2(new_n964), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n559), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT59), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1098), .A2(KEYINPUT120), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT120), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1008), .A2(new_n815), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1037), .A2(new_n782), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n608), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n616), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1114), .B1(new_n1113), .B2(new_n1110), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1106), .A2(new_n1107), .A3(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1111), .A2(new_n608), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1092), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1093), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1072), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1026), .A2(new_n1030), .A3(new_n1123), .A4(new_n1031), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1063), .A2(new_n1122), .A3(new_n1011), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1053), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1029), .A2(new_n1017), .A3(G286), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  OAI21_X1  g703(.A(G8), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1049), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1127), .A3(new_n1131), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1060), .A2(new_n1127), .A3(new_n1052), .A4(new_n1045), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(KEYINPUT63), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1052), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1045), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1040), .A2(new_n714), .A3(new_n710), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1038), .B1(new_n1137), .B2(new_n1033), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1125), .A2(new_n1134), .A3(new_n1136), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1121), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G290), .B(G1986), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n981), .B1(new_n965), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT125), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1098), .A2(new_n1105), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1098), .A2(new_n1105), .A3(KEYINPUT120), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1115), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1071), .B1(new_n1150), .B2(new_n1119), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT125), .B(new_n1143), .C1(new_n1151), .C2(new_n1139), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n986), .B1(new_n1144), .B2(new_n1153), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g729(.A(G227), .B1(new_n646), .B2(G14), .ZN(new_n1156));
  AND2_X1   g730(.A1(new_n896), .A2(new_n1156), .ZN(new_n1157));
  AND4_X1   g731(.A1(G319), .A2(new_n956), .A3(new_n685), .A4(new_n1157), .ZN(G308));
  NAND4_X1  g732(.A1(new_n956), .A2(new_n1157), .A3(G319), .A4(new_n685), .ZN(G225));
endmodule


