//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT73), .ZN(new_n194));
  XNOR2_X1  g008(.A(G110), .B(G140), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n199), .B1(KEYINPUT11), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G134), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT65), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT65), .B(new_n204), .C1(new_n200), .C2(G137), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n202), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n202), .B(new_n210), .C1(new_n205), .C2(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT12), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(KEYINPUT77), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n232), .A3(G146), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  AND4_X1   g049(.A1(new_n228), .A2(new_n233), .A3(G128), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n235), .ZN(new_n237));
  AOI21_X1  g051(.A(G146), .B1(new_n230), .B2(new_n232), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n228), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n236), .B1(new_n241), .B2(KEYINPUT74), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT74), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(new_n237), .C1(new_n239), .C2(new_n240), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n227), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n229), .A2(G146), .ZN(new_n247));
  OAI21_X1  g061(.A(G128), .B1(new_n247), .B2(new_n228), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n234), .A2(G143), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(KEYINPUT66), .C1(new_n238), .C2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n249), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(G143), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT66), .B1(new_n254), .B2(new_n248), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n246), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n227), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n215), .B1(new_n245), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT77), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT12), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(KEYINPUT76), .A3(KEYINPUT10), .A4(new_n257), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT76), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n230), .A2(new_n232), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n249), .B1(new_n266), .B2(new_n234), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n240), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n236), .B1(new_n269), .B2(new_n250), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n257), .A2(KEYINPUT10), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n267), .A2(new_n276), .B1(new_n237), .B2(new_n273), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G101), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n282), .A3(G101), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n263), .A2(new_n272), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n231), .A2(G143), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n234), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n240), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n247), .B1(new_n253), .B2(G146), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT74), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n246), .A3(new_n244), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n257), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n286), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI211_X1 g110(.A(KEYINPUT75), .B(KEYINPUT10), .C1(new_n293), .C2(new_n257), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n285), .B(new_n213), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n197), .B1(new_n262), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n285), .B1(new_n296), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n212), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(KEYINPUT78), .A3(new_n212), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(new_n305), .B2(new_n197), .ZN(new_n306));
  OAI21_X1  g120(.A(G469), .B1(new_n306), .B2(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n196), .A3(new_n304), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n262), .A2(new_n197), .A3(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G469), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n190), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n191), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(G234), .B2(new_n190), .ZN(new_n315));
  XOR2_X1   g129(.A(G119), .B(G128), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT24), .B(G110), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G128), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(G119), .C2(new_n240), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n318), .B1(G110), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT71), .A3(G140), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n328), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n329), .A2(KEYINPUT71), .A3(G140), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT72), .B1(new_n339), .B2(new_n328), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(G146), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n336), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n324), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n323), .A2(G110), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n316), .A2(new_n317), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n345), .A2(new_n346), .B1(new_n234), .B2(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n349), .B(new_n350), .Z(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  INV_X1    g167(.A(new_n324), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n332), .A2(new_n333), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n356));
  INV_X1    g170(.A(new_n327), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n334), .A2(new_n335), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n234), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n354), .B1(new_n360), .B2(new_n341), .ZN(new_n361));
  INV_X1    g175(.A(new_n348), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n352), .A2(new_n363), .A3(new_n190), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n315), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n352), .A2(new_n363), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n315), .A2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G472), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n320), .A2(G116), .ZN(new_n376));
  INV_X1    g190(.A(G116), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G119), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT2), .B(G113), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT2), .B(G113), .Z(new_n385));
  XNOR2_X1  g199(.A(G116), .B(G119), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT67), .A3(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n199), .B2(new_n201), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n211), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n269), .A2(new_n250), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(new_n246), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n277), .B1(new_n211), .B2(new_n209), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT30), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n397));
  INV_X1    g211(.A(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n256), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n212), .A2(new_n278), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n397), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n390), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G237), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n192), .A3(G210), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n404), .B(KEYINPUT27), .Z(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT26), .B(G101), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n399), .A2(new_n400), .A3(new_n389), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT31), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n394), .A2(new_n390), .A3(new_n395), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT30), .B1(new_n394), .B2(new_n395), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n399), .A2(new_n397), .A3(new_n400), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n413), .B1(new_n416), .B2(new_n390), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT31), .A3(new_n408), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n389), .B1(new_n399), .B2(new_n400), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT28), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n407), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n374), .B1(new_n419), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n407), .B1(new_n422), .B2(new_n425), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n389), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n431), .A2(new_n408), .A3(new_n413), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n429), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n409), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT28), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n438), .A2(KEYINPUT29), .A3(new_n408), .A4(new_n425), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n439), .A3(new_n190), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n428), .A2(KEYINPUT32), .B1(new_n440), .B2(G472), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT31), .B1(new_n417), .B2(new_n408), .ZN(new_n442));
  NOR4_X1   g256(.A1(new_n431), .A2(new_n411), .A3(new_n407), .A4(new_n413), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n427), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n373), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT69), .B(KEYINPUT32), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n372), .B1(new_n441), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G210), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n384), .A2(new_n281), .A3(new_n388), .A4(new_n283), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n227), .A2(new_n383), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n386), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n460));
  INV_X1    g274(.A(new_n376), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n462), .A3(G113), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n452), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n452), .A2(new_n466), .A3(new_n464), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n471), .A3(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n246), .B(new_n329), .C1(new_n251), .C2(new_n255), .ZN(new_n474));
  INV_X1    g288(.A(G224), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(G953), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n277), .A2(G125), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n474), .B2(new_n478), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n473), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n477), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n479), .B2(new_n480), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n452), .A2(new_n464), .ZN(new_n490));
  INV_X1    g304(.A(G113), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n460), .B2(new_n461), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n383), .B1(new_n459), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT83), .B1(new_n493), .B2(new_n257), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n463), .A2(new_n387), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT83), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n227), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n492), .B1(new_n454), .B2(new_n379), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n453), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n466), .B(KEYINPUT8), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n490), .A2(new_n466), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n474), .A2(new_n478), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n487), .A3(new_n477), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n489), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n190), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n451), .B1(new_n486), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n476), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n481), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n472), .B(new_n470), .C1(new_n483), .C2(new_n511), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n512), .A2(new_n190), .A3(new_n450), .A4(new_n505), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(KEYINPUT84), .B(new_n451), .C1(new_n486), .C2(new_n506), .ZN(new_n515));
  OAI21_X1  g329(.A(G214), .B1(G237), .B2(G902), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n516), .B(KEYINPUT79), .Z(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G952), .A3(new_n192), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(G902), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n192), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n515), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(G104), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n403), .A2(new_n192), .A3(G214), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n530), .A2(new_n229), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n253), .A2(new_n530), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n210), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n531), .A2(new_n532), .A3(new_n210), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n360), .A2(new_n341), .A3(new_n534), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n531), .A2(new_n532), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT18), .A3(G131), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT85), .B1(new_n338), .B2(new_n234), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n355), .B2(new_n234), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n339), .A2(KEYINPUT85), .A3(G146), .ZN(new_n544));
  NAND2_X1  g358(.A1(KEYINPUT18), .A2(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n531), .A2(new_n532), .A3(new_n545), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n529), .B1(new_n539), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n529), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n535), .A2(new_n537), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n341), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n355), .A2(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(KEYINPUT19), .B2(new_n338), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT86), .A3(new_n234), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT86), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n338), .A2(KEYINPUT19), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n355), .B2(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n557), .B2(G146), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n549), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n548), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT20), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n527), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n539), .A2(new_n547), .ZN(new_n566));
  INV_X1    g380(.A(new_n529), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n560), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n561), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n564), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n566), .B1(new_n574), .B2(new_n567), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n529), .A4(new_n547), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n190), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(G475), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n377), .A2(G122), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT14), .Z(new_n582));
  INV_X1    g396(.A(KEYINPUT89), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n377), .B2(G122), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT89), .A3(G116), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n219), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n581), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(KEYINPUT90), .A3(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n588), .B1(new_n593), .B2(new_n219), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n230), .A2(new_n232), .A3(G128), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT91), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT91), .A4(G128), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n229), .A2(G128), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT93), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n603), .B(new_n600), .C1(new_n597), .C2(new_n598), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n602), .A2(new_n604), .A3(new_n200), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT91), .B1(new_n253), .B2(G128), .ZN(new_n606));
  AND4_X1   g420(.A1(KEYINPUT91), .A2(new_n230), .A3(new_n232), .A4(G128), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n603), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(KEYINPUT93), .A3(new_n601), .ZN(new_n610));
  AOI21_X1  g424(.A(G134), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n594), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n188), .A2(new_n314), .A3(G953), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT13), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n600), .B1(new_n599), .B2(new_n614), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(KEYINPUT92), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT13), .B1(new_n597), .B2(new_n598), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n600), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n200), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n200), .B1(new_n602), .B2(new_n604), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n593), .A2(new_n219), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n591), .A2(G107), .A3(new_n592), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n612), .B(new_n613), .C1(new_n621), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT94), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n599), .A2(new_n614), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT92), .A3(new_n601), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n630), .B(new_n620), .C1(new_n614), .C2(new_n599), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(G134), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n622), .A2(new_n625), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n612), .A4(new_n613), .ZN(new_n636));
  INV_X1    g450(.A(new_n613), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n621), .A2(new_n626), .ZN(new_n638));
  INV_X1    g452(.A(new_n588), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n623), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n609), .A2(G134), .A3(new_n610), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n622), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n637), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n628), .A2(new_n636), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n190), .ZN(new_n645));
  INV_X1    g459(.A(G478), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(KEYINPUT15), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n644), .B(new_n190), .C1(KEYINPUT15), .C2(new_n646), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n526), .A2(new_n580), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n313), .A2(new_n449), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  AOI21_X1  g468(.A(G478), .B1(new_n644), .B2(new_n190), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n642), .B1(new_n632), .B2(new_n633), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n613), .A2(KEYINPUT95), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n644), .A2(new_n656), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n646), .A2(G902), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n655), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n573), .A2(new_n579), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n654), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n644), .A2(new_n656), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g482(.A(KEYINPUT96), .B(new_n580), .C1(new_n668), .C2(new_n655), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n516), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n507), .B2(new_n513), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n524), .ZN(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n444), .B2(new_n190), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n676), .A2(new_n428), .A3(new_n372), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n313), .A2(new_n670), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G104), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G6));
  INV_X1    g495(.A(new_n524), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n578), .B1(new_n648), .B2(new_n649), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n565), .A2(new_n571), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n684), .B1(new_n565), .B2(new_n571), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n572), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n682), .A2(new_n683), .A3(new_n687), .A4(new_n672), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n313), .A2(new_n688), .A3(new_n677), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT35), .B(G107), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  NOR2_X1   g505(.A1(new_n676), .A2(new_n428), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n344), .A2(new_n348), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n370), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n368), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n313), .A2(new_n651), .A3(new_n692), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  NOR2_X1   g514(.A1(new_n192), .A2(G900), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OR3_X1    g516(.A1(new_n702), .A2(KEYINPUT99), .A3(new_n521), .ZN(new_n703));
  OAI21_X1  g517(.A(KEYINPUT99), .B1(new_n702), .B2(new_n521), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n519), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n683), .A2(new_n687), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT100), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n683), .A2(new_n687), .A3(new_n708), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(G469), .A2(G902), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n298), .A2(new_n302), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT75), .B1(new_n245), .B2(KEYINPUT10), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n294), .A2(new_n286), .A3(new_n295), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n213), .B1(new_n716), .B2(new_n285), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n304), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n197), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT12), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n215), .B(new_n261), .C1(new_n245), .C2(new_n258), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n298), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n196), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n720), .A2(G469), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n312), .A2(new_n712), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n191), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n444), .A2(KEYINPUT32), .A3(new_n373), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n440), .A2(G472), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n448), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n672), .A3(new_n697), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n711), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n697), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n441), .B2(new_n448), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n313), .A2(new_n738), .A3(new_n672), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT101), .B1(new_n739), .B2(new_n710), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT102), .B(G128), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G30));
  NAND2_X1  g557(.A1(new_n448), .A2(new_n730), .ZN(new_n744));
  INV_X1    g558(.A(new_n436), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n409), .A2(new_n434), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n407), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n408), .B1(new_n431), .B2(new_n413), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n190), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(KEYINPUT103), .A3(G472), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT103), .B1(new_n749), .B2(G472), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n737), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n650), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n664), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n753), .A2(new_n756), .A3(new_n671), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n514), .A2(new_n515), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT38), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT104), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n705), .B(KEYINPUT39), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n313), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT40), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n266), .B(KEYINPUT105), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G45));
  NOR2_X1   g581(.A1(new_n663), .A2(new_n664), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n705), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n739), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n234), .ZN(G48));
  AOI21_X1  g585(.A(new_n311), .B1(new_n310), .B2(new_n190), .ZN(new_n772));
  AOI211_X1 g586(.A(G469), .B(G902), .C1(new_n308), .C2(new_n309), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n191), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n670), .A3(new_n449), .A4(new_n674), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT41), .B(G113), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT107), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT106), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n775), .B(new_n778), .ZN(G15));
  NAND3_X1  g593(.A1(new_n774), .A2(new_n449), .A3(new_n688), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G116), .ZN(G18));
  NOR3_X1   g595(.A1(new_n650), .A2(new_n580), .A3(new_n524), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT108), .B1(new_n774), .B2(new_n672), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n310), .A2(new_n190), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(G469), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n728), .A3(new_n312), .A4(new_n672), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n738), .B(new_n782), .C1(new_n783), .C2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G119), .ZN(G21));
  NAND2_X1  g604(.A1(new_n438), .A2(new_n425), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n407), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n374), .B1(new_n419), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n676), .A2(new_n793), .A3(new_n372), .A4(new_n524), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n772), .A2(new_n773), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n650), .A2(new_n580), .A3(new_n672), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n728), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G122), .ZN(G24));
  NOR2_X1   g612(.A1(new_n676), .A2(new_n793), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n768), .A2(new_n697), .A3(new_n799), .A4(new_n705), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n786), .A2(new_n787), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n795), .A2(KEYINPUT108), .A3(new_n728), .A4(new_n672), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n329), .ZN(G27));
  INV_X1    g618(.A(KEYINPUT32), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n445), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n730), .A3(new_n731), .ZN(new_n807));
  INV_X1    g621(.A(new_n372), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n768), .A3(new_n808), .A4(new_n705), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n299), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n725), .A2(KEYINPUT109), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n720), .A2(new_n811), .A3(new_n812), .A4(G469), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n312), .A2(new_n813), .A3(new_n712), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n191), .B(new_n671), .C1(new_n514), .C2(new_n515), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT42), .B1(new_n809), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n705), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n663), .A2(new_n664), .A3(KEYINPUT42), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n449), .A2(new_n819), .A3(new_n815), .A4(new_n814), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G131), .ZN(G33));
  NAND4_X1  g636(.A1(new_n814), .A2(new_n732), .A3(new_n815), .A4(new_n808), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n710), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(new_n200), .ZN(G36));
  NAND4_X1  g639(.A1(new_n720), .A2(new_n811), .A3(new_n812), .A4(KEYINPUT45), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(G469), .C1(KEYINPUT45), .C2(new_n306), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n827), .A2(new_n712), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT46), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n312), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(KEYINPUT110), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(KEYINPUT110), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n728), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n762), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n671), .B1(new_n514), .B2(new_n515), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n661), .A2(new_n662), .ZN(new_n839));
  INV_X1    g653(.A(new_n655), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n664), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT43), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n843), .A2(new_n692), .A3(new_n737), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT44), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n836), .B(new_n846), .C1(new_n845), .C2(new_n844), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G137), .ZN(G39));
  NAND2_X1  g662(.A1(new_n835), .A2(KEYINPUT47), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT47), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n834), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n769), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n838), .A2(new_n732), .A3(new_n808), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(G140), .ZN(G42));
  NOR4_X1   g670(.A1(new_n759), .A2(new_n191), .A3(new_n517), .A4(new_n842), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n744), .A2(new_n372), .A3(new_n752), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n795), .B(KEYINPUT49), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n843), .A2(new_n519), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n795), .A3(new_n815), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n807), .A2(new_n808), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT48), .Z(new_n865));
  NAND4_X1  g679(.A1(new_n858), .A2(new_n520), .A3(new_n795), .A4(new_n815), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n665), .B2(new_n669), .ZN(new_n867));
  INV_X1    g681(.A(G952), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n867), .A2(new_n868), .A3(G953), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n783), .A2(new_n788), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n861), .A2(new_n808), .A3(new_n799), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n865), .B(new_n869), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n795), .A2(new_n191), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n849), .A2(new_n851), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n871), .A2(new_n838), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT115), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n759), .A2(new_n516), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n774), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT50), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n862), .A2(new_n676), .A3(new_n737), .A4(new_n793), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n866), .A2(new_n580), .A3(new_n841), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n887));
  OAI211_X1 g701(.A(KEYINPUT51), .B(new_n882), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n873), .B1(new_n878), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n882), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n882), .B2(new_n885), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n875), .A2(new_n877), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n889), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n818), .A2(new_n191), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n650), .A2(new_n580), .A3(new_n672), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n753), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n734), .A2(new_n853), .B1(new_n899), .B2(new_n814), .ZN(new_n900));
  INV_X1    g714(.A(new_n800), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n783), .B2(new_n788), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n735), .B1(new_n711), .B2(new_n734), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n739), .A2(new_n710), .A3(KEYINPUT101), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n900), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n803), .B1(new_n736), .B2(new_n740), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .A3(new_n900), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT111), .B1(new_n841), .B2(new_n580), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n650), .A2(new_n664), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n664), .B2(new_n663), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(KEYINPUT111), .ZN(new_n914));
  INV_X1    g728(.A(new_n526), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n727), .A2(new_n915), .A3(new_n728), .A4(new_n677), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n652), .B(new_n797), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n775), .A2(new_n698), .A3(new_n780), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n920), .A3(new_n789), .ZN(new_n921));
  OAI22_X1  g735(.A1(new_n710), .A2(new_n823), .B1(new_n816), .B2(new_n800), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n727), .A2(new_n732), .A3(new_n728), .A4(new_n697), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT112), .ZN(new_n924));
  INV_X1    g738(.A(new_n572), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n565), .A2(new_n571), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT98), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n565), .A2(new_n571), .A3(new_n684), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n578), .A2(new_n818), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n648), .A2(new_n930), .A3(new_n649), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n932), .B2(new_n837), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n648), .A2(new_n930), .A3(new_n649), .ZN(new_n934));
  AND4_X1   g748(.A1(new_n924), .A2(new_n837), .A3(new_n934), .A4(new_n687), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n923), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n922), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n821), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n921), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n910), .A2(KEYINPUT53), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT114), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n917), .A2(new_n919), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n789), .A3(new_n821), .A4(new_n937), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n907), .B2(new_n909), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT114), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT53), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT54), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT113), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n944), .B2(KEYINPUT53), .ZN(new_n950));
  AND4_X1   g764(.A1(KEYINPUT52), .A2(new_n741), .A3(new_n902), .A4(new_n900), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT52), .B1(new_n908), .B2(new_n900), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n939), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT53), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n953), .A2(KEYINPUT113), .A3(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n940), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n944), .A2(KEYINPUT53), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT54), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n896), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT118), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n868), .A2(new_n192), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n961), .A2(KEYINPUT118), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n860), .B1(new_n964), .B2(new_n965), .ZN(G75));
  NOR2_X1   g780(.A1(new_n192), .A2(G952), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n484), .A2(new_n473), .A3(new_n485), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n512), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT55), .Z(new_n970));
  AND2_X1   g784(.A1(new_n950), .A2(new_n955), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n190), .B1(new_n971), .B2(new_n947), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(G210), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT56), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n974), .A3(new_n970), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT119), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT119), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(new_n978), .A3(new_n974), .A4(new_n970), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n967), .B(new_n975), .C1(new_n977), .C2(new_n979), .ZN(G51));
  XOR2_X1   g794(.A(new_n712), .B(KEYINPUT57), .Z(new_n981));
  AND4_X1   g795(.A1(new_n945), .A2(new_n910), .A3(KEYINPUT53), .A4(new_n939), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n945), .B1(new_n944), .B2(KEYINPUT53), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n950), .A2(new_n955), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT54), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n948), .B1(new_n971), .B2(new_n947), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n310), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n827), .B(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n972), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n967), .B1(new_n989), .B2(new_n991), .ZN(G54));
  NAND3_X1  g806(.A1(new_n972), .A2(KEYINPUT58), .A3(G475), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n568), .A2(new_n569), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n967), .ZN(G60));
  INV_X1    g811(.A(new_n661), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT59), .Z(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n986), .B2(new_n987), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT121), .ZN(new_n1003));
  INV_X1    g817(.A(new_n967), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1001), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT54), .B1(new_n984), .B2(new_n985), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n956), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT121), .B1(new_n1008), .B2(new_n967), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n998), .B1(new_n960), .B2(new_n1000), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT122), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .A4(KEYINPUT122), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(G63));
  NAND2_X1  g829(.A1(G217), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT60), .Z(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n984), .B2(new_n985), .ZN(new_n1018));
  INV_X1    g832(.A(new_n369), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n695), .B(new_n1017), .C1(new_n984), .C2(new_n985), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1020), .A2(new_n1004), .A3(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1021), .A2(KEYINPUT123), .A3(new_n1004), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT124), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT61), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1023), .B2(KEYINPUT61), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1022), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(KEYINPUT124), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1022), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1023), .A2(new_n1024), .A3(KEYINPUT61), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1027), .A2(new_n1032), .ZN(G66));
  OAI21_X1  g847(.A(G953), .B1(new_n523), .B2(new_n475), .ZN(new_n1034));
  INV_X1    g848(.A(new_n921), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n473), .B1(G898), .B2(new_n192), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(G69));
  OAI21_X1  g852(.A(new_n908), .B1(new_n739), .B2(new_n769), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n821), .B1(new_n710), .B2(new_n823), .ZN(new_n1040));
  NOR3_X1   g854(.A1(new_n756), .A2(new_n863), .A3(new_n673), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n1039), .B(new_n1040), .C1(new_n836), .C2(new_n1041), .ZN(new_n1042));
  AND3_X1   g856(.A1(new_n1042), .A2(new_n847), .A3(new_n855), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n702), .B1(new_n1043), .B2(G953), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n557), .B(KEYINPUT125), .Z(new_n1045));
  XNOR2_X1  g859(.A(new_n416), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g861(.A1(G227), .A2(G900), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(G953), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1046), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n855), .A2(new_n847), .ZN(new_n1051));
  OR3_X1    g865(.A1(new_n765), .A2(KEYINPUT62), .A3(new_n1039), .ZN(new_n1052));
  OAI21_X1  g866(.A(KEYINPUT62), .B1(new_n765), .B2(new_n1039), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n449), .A2(new_n837), .ZN(new_n1054));
  OR3_X1    g868(.A1(new_n914), .A2(new_n763), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1050), .B1(new_n1057), .B2(G953), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1047), .A2(new_n1049), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g873(.A(G953), .B(new_n1048), .C1(new_n1044), .C2(new_n1050), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1059), .A2(new_n1060), .ZN(G72));
  INV_X1    g875(.A(new_n748), .ZN(new_n1062));
  XOR2_X1   g876(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1063));
  NOR2_X1   g877(.A1(new_n675), .A2(new_n190), .ZN(new_n1064));
  XNOR2_X1  g878(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1062), .A2(new_n432), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n957), .B2(new_n958), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1065), .B1(new_n1043), .B2(new_n1035), .ZN(new_n1068));
  INV_X1    g882(.A(new_n432), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1004), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g884(.A1(new_n1051), .A2(new_n921), .A3(new_n1056), .ZN(new_n1071));
  OAI21_X1  g885(.A(new_n1062), .B1(new_n1071), .B2(new_n1065), .ZN(new_n1072));
  OR2_X1    g886(.A1(new_n1072), .A2(KEYINPUT127), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1072), .A2(KEYINPUT127), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(G57));
endmodule


