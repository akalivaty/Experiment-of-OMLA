//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n599, new_n602, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  NOR2_X1   g049(.A1(new_n465), .A2(new_n472), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n465), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND3_X1  g057(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n483));
  NAND2_X1  g058(.A1(G114), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n461), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G102), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n472), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n486), .A2(new_n488), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  XNOR2_X1  g070(.A(KEYINPUT67), .B(G651), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G75), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT68), .A3(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n497), .A2(G62), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n509), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND3_X1  g095(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n504), .A2(new_n505), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n517), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n521), .B(new_n523), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n506), .A2(new_n513), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(new_n514), .A2(new_n516), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n506), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(new_n534), .C1(new_n496), .C2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT69), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n531), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n497), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT70), .Z(new_n543));
  NAND3_X1  g118(.A1(new_n524), .A2(G43), .A3(G543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n524), .A2(G81), .A3(new_n517), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n531), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n532), .A2(G91), .B1(G651), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n528), .A2(new_n561), .A3(G53), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n561), .B1(new_n528), .B2(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n532), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n528), .A2(G49), .ZN(new_n567));
  INV_X1    g142(.A(G74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n500), .B1(new_n531), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT72), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n528), .A2(G48), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n532), .A2(G86), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n517), .A2(KEYINPUT73), .A3(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n531), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(new_n497), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n572), .A2(new_n573), .A3(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(new_n532), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n528), .A2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n496), .C2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n525), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n500), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n528), .A2(G54), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n532), .A2(new_n592), .A3(G92), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n586), .B1(G868), .B2(new_n595), .ZN(G284));
  OAI21_X1  g171(.A(new_n586), .B1(G868), .B2(new_n595), .ZN(G321));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G299), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G297));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(G280));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n602), .B2(G860), .ZN(G148));
  NOR2_X1   g178(.A1(new_n550), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n595), .A2(new_n602), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(G868), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT74), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n475), .A2(G123), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n477), .A2(G135), .ZN(new_n610));
  NOR2_X1   g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(G2096), .Z(new_n614));
  NAND2_X1  g189(.A1(new_n492), .A2(new_n487), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT13), .B(G2100), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n614), .A2(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2430), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2435), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2438), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2451), .B(G2454), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT76), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT16), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT77), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n631), .B2(new_n633), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n635), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT79), .Z(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT17), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT80), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n643), .A2(new_n644), .ZN(new_n649));
  INV_X1    g224(.A(new_n646), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n650), .C1(new_n645), .C2(new_n643), .ZN(new_n651));
  INV_X1    g226(.A(new_n644), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n652), .A2(new_n646), .A3(new_n642), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT18), .Z(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2100), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n661), .A2(new_n664), .A3(new_n668), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G1981), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G35), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G162), .B2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT29), .Z(new_n682));
  INV_X1    g257(.A(G2090), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT96), .ZN(new_n685));
  MUX2_X1   g260(.A(G24), .B(G290), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1986), .ZN(new_n687));
  AOI22_X1  g262(.A1(G119), .A2(new_n475), .B1(new_n477), .B2(G131), .ZN(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n689));
  NOR2_X1   g264(.A1(G95), .A2(G2105), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT83), .Z(new_n691));
  OAI21_X1  g266(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n692), .S(G29), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT35), .B(G1991), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT84), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n693), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(G1971), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G16), .B2(G23), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(G1971), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n703), .B(new_n705), .C1(G16), .C2(G23), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n701), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G6), .B(G305), .S(G16), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n711), .A2(KEYINPUT34), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT34), .B1(new_n711), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n697), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(new_n697), .C1(new_n715), .C2(new_n716), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n685), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT89), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2105), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n477), .A2(G139), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G103), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT25), .Z(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n724), .A2(KEYINPUT90), .A3(new_n725), .A4(new_n727), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n730), .A2(KEYINPUT91), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(KEYINPUT91), .B1(new_n730), .B2(new_n731), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n732), .A2(new_n733), .A3(new_n679), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n679), .A2(G33), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(KEYINPUT92), .B2(G2072), .ZN(new_n736));
  NAND2_X1  g311(.A1(KEYINPUT92), .A2(G2072), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n736), .B(new_n737), .Z(new_n738));
  NOR2_X1   g313(.A1(G5), .A2(G16), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G171), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n698), .A2(KEYINPUT23), .A3(G20), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n744));
  INV_X1    g319(.A(G20), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G16), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n743), .B(new_n746), .C1(new_n599), .C2(new_n698), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT30), .B(G28), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n679), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n721), .A2(new_n738), .A3(new_n742), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n477), .A2(G141), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n475), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n487), .A2(G105), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G32), .B(new_n761), .S(G29), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT27), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1996), .ZN(new_n764));
  INV_X1    g339(.A(G19), .ZN(new_n765));
  OAI21_X1  g340(.A(KEYINPUT85), .B1(new_n765), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n765), .A2(KEYINPUT85), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n550), .C2(new_n698), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT86), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G1341), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(G1341), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n764), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n679), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n679), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n773), .B(new_n774), .S(KEYINPUT95), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n682), .A2(new_n683), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT97), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n698), .A2(G4), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n595), .B2(new_n698), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1348), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n698), .A2(G21), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G168), .B2(new_n698), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1966), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n679), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n475), .A2(new_n790), .A3(G128), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n492), .A2(G2105), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT87), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n477), .A2(G140), .ZN(new_n795));
  OR2_X1    g370(.A1(G104), .A2(G2105), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n796), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n791), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n789), .B1(new_n799), .B2(new_n679), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT31), .B(G11), .Z(new_n802));
  NOR4_X1   g377(.A1(new_n783), .A2(new_n786), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n772), .A2(new_n777), .A3(new_n780), .A4(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G34), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(KEYINPUT24), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(KEYINPUT24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n679), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G160), .B2(new_n679), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G2084), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n613), .A2(new_n679), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n751), .A2(new_n804), .A3(new_n810), .A4(new_n811), .ZN(G311));
  INV_X1    g387(.A(new_n751), .ZN(new_n813));
  INV_X1    g388(.A(new_n810), .ZN(new_n814));
  INV_X1    g389(.A(new_n811), .ZN(new_n815));
  INV_X1    g390(.A(new_n804), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(new_n532), .A2(G93), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT99), .B(G55), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n528), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n496), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n595), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT39), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n818), .A2(new_n822), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(new_n820), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(new_n549), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n823), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n829), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n825), .B1(new_n836), .B2(G860), .ZN(G145));
  NAND2_X1  g412(.A1(new_n799), .A2(new_n494), .ZN(new_n838));
  NAND2_X1  g413(.A1(G164), .A2(new_n798), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n759), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n759), .B1(new_n838), .B2(new_n839), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n760), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n844), .A2(KEYINPUT94), .A3(new_n840), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n845), .C1(new_n732), .C2(new_n733), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n730), .A2(new_n731), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n847), .A2(new_n840), .A3(new_n844), .ZN(new_n848));
  AOI22_X1  g423(.A1(G130), .A2(new_n475), .B1(new_n477), .B2(G142), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n851), .B(new_n852), .C1(G118), .C2(new_n472), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n692), .B(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(new_n617), .Z(new_n856));
  AND3_X1   g431(.A1(new_n846), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n846), .B2(new_n848), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G160), .B(KEYINPUT100), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n613), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT102), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n859), .B2(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  INV_X1    g440(.A(new_n862), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n865), .B(new_n866), .C1(new_n857), .C2(new_n858), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n863), .A2(new_n864), .A3(new_n870), .A4(new_n867), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(KEYINPUT40), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(KEYINPUT40), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(G395));
  NOR2_X1   g449(.A1(new_n823), .A2(G868), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(KEYINPUT104), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(new_n560), .C1(new_n562), .C2(new_n563), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n595), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(G299), .A2(new_n594), .A3(KEYINPUT104), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n879), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n879), .A2(new_n880), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n835), .B(new_n605), .ZN(new_n885));
  MUX2_X1   g460(.A(new_n883), .B(new_n884), .S(new_n885), .Z(new_n886));
  INV_X1    g461(.A(KEYINPUT106), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G303), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G305), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n702), .B(KEYINPUT105), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n886), .B2(new_n887), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n875), .B1(new_n897), .B2(G868), .ZN(G295));
  AOI21_X1  g473(.A(new_n875), .B1(new_n897), .B2(G868), .ZN(G331));
  XOR2_X1   g474(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n900));
  NAND3_X1  g475(.A1(new_n549), .A2(new_n830), .A3(new_n820), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n901), .A2(G286), .A3(new_n833), .ZN(new_n902));
  AOI21_X1  g477(.A(G286), .B1(new_n901), .B2(new_n833), .ZN(new_n903));
  OAI21_X1  g478(.A(G171), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(G168), .B1(new_n832), .B2(new_n834), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(G286), .A3(new_n833), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(G301), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n883), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n909));
  INV_X1    g484(.A(new_n891), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n890), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n904), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n884), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n883), .A2(new_n904), .A3(new_n907), .A4(new_n914), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n909), .A2(new_n911), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n908), .A2(KEYINPUT108), .B1(new_n912), .B2(new_n884), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n911), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n900), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n908), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n892), .ZN(new_n924));
  INV_X1    g499(.A(new_n900), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n924), .A2(new_n916), .A3(new_n917), .A4(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n921), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n915), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n892), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(new_n917), .A3(new_n916), .A4(new_n925), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n916), .A3(new_n917), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n922), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(new_n933), .ZN(G397));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  INV_X1    g510(.A(new_n484), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n492), .B2(G126), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n488), .B1(new_n937), .B2(new_n472), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n491), .A2(new_n493), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n468), .A2(new_n473), .A3(G40), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n692), .B(new_n695), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT111), .Z(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n798), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(G1996), .B1(new_n755), .B2(new_n758), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n948), .B(new_n949), .C1(new_n761), .C2(G1996), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n944), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(G290), .A2(G1986), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n944), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT48), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n942), .A2(G1996), .A3(new_n943), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT46), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n948), .A2(new_n759), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n944), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(KEYINPUT46), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n692), .A2(new_n695), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n950), .A2(new_n963), .B1(G2067), .B2(new_n798), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n944), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n955), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT127), .Z(new_n967));
  NAND2_X1  g542(.A1(G303), .A2(G8), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT55), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n942), .B1(new_n971), .B2(KEYINPUT113), .ZN(new_n972));
  INV_X1    g547(.A(new_n943), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n491), .A2(new_n493), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n485), .A2(G2105), .B1(G102), .B2(new_n487), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n976), .A2(KEYINPUT113), .A3(KEYINPUT45), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1971), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n943), .B1(new_n940), .B2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n981), .B(new_n935), .C1(new_n938), .C2(new_n939), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT114), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n494), .A2(new_n984), .A3(new_n981), .A4(new_n935), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n978), .A2(new_n979), .B1(new_n986), .B2(new_n683), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n969), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n580), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G1981), .ZN(new_n992));
  NOR2_X1   g567(.A1(G305), .A2(KEYINPUT49), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  AOI22_X1  g569(.A1(G86), .A2(new_n532), .B1(new_n579), .B2(new_n497), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(new_n572), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G305), .A2(KEYINPUT49), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(new_n994), .A3(new_n572), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(G1981), .A3(new_n999), .A4(new_n991), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n940), .A2(new_n943), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n988), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n997), .A2(new_n1000), .A3(KEYINPUT117), .A4(new_n1002), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n566), .A2(new_n567), .A3(G1976), .A4(new_n570), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  INV_X1    g585(.A(G1976), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G288), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1002), .A2(new_n1012), .A3(new_n1013), .A4(new_n1008), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n989), .A2(new_n1007), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT119), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n987), .A2(new_n988), .A3(new_n969), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1007), .A2(new_n989), .A3(new_n1017), .A4(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1019), .A2(KEYINPUT63), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1966), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n943), .B1(new_n940), .B2(new_n941), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n970), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n494), .B2(new_n935), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n1028), .A2(KEYINPUT118), .A3(new_n943), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n986), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n988), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G168), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n980), .A2(new_n982), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(G2090), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n978), .B2(new_n979), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n969), .B1(new_n1037), .B2(new_n988), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1020), .A2(new_n1007), .A3(new_n1017), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1023), .A2(new_n1034), .B1(new_n1040), .B2(KEYINPUT63), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(new_n1020), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1007), .A2(new_n1011), .A3(new_n702), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(G1981), .B2(G305), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1002), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT118), .B1(new_n1028), .B2(new_n943), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n942), .A2(new_n1026), .A3(new_n973), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n970), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1050), .A2(new_n1024), .B1(new_n986), .B2(new_n1031), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT125), .B1(new_n1051), .B2(new_n988), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n973), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n971), .B1(new_n1055), .B2(KEYINPUT118), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1966), .B1(new_n1056), .B2(new_n1049), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G2084), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1054), .B(G8), .C1(new_n1057), .C2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(G168), .A2(new_n988), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1052), .A2(new_n1053), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT51), .B(G8), .C1(new_n1064), .C2(G286), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT124), .B(KEYINPUT51), .C1(new_n1033), .C2(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1064), .A2(new_n1061), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n978), .A2(G2078), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1073), .A2(new_n1074), .B1(new_n741), .B2(new_n1058), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1050), .A2(G2078), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT126), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT62), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1069), .A2(new_n1081), .A3(new_n1070), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1072), .A2(G171), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(G1956), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1035), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT120), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  XOR2_X1   g662(.A(new_n1087), .B(KEYINPUT122), .Z(new_n1088));
  OR2_X1    g663(.A1(new_n978), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n560), .B2(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(G299), .B(new_n1092), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1086), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1058), .A2(new_n1096), .B1(new_n947), .B2(new_n1001), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n594), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT58), .B(G1341), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n978), .A2(G1996), .B1(new_n1001), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT123), .A3(new_n550), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1097), .A2(new_n594), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT60), .B1(new_n1105), .B2(new_n1098), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1101), .A2(KEYINPUT123), .A3(KEYINPUT59), .A4(new_n550), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(new_n1108), .A3(new_n595), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1104), .A2(new_n1106), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1095), .A2(KEYINPUT61), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1086), .A2(new_n1089), .A3(new_n1112), .A4(new_n1093), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1094), .B(new_n1099), .C1(new_n1110), .C2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G301), .B(KEYINPUT54), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n1055), .A2(new_n971), .A3(new_n1074), .A4(G2078), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n1075), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1080), .A2(new_n1116), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n1119), .A3(new_n1120), .A4(new_n1071), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1083), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1039), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1047), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n952), .ZN(new_n1125));
  NAND2_X1  g700(.A1(G290), .A2(G1986), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT109), .A3(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n944), .C1(KEYINPUT109), .C2(new_n1126), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT110), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n951), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT112), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n967), .B1(new_n1124), .B2(new_n1131), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g707(.A1(new_n921), .A2(new_n926), .ZN(new_n1134));
  AND3_X1   g708(.A1(new_n868), .A2(new_n640), .A3(new_n657), .ZN(new_n1135));
  NAND4_X1  g709(.A1(new_n1134), .A2(new_n1135), .A3(G319), .A4(new_n677), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


