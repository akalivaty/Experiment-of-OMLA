

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769;

  NOR2_X1 U362 ( .A1(n767), .A2(n765), .ZN(n592) );
  NOR2_X1 U363 ( .A1(n595), .A2(n594), .ZN(n673) );
  XNOR2_X1 U364 ( .A(KEYINPUT39), .B(n579), .ZN(n607) );
  NOR2_X1 U365 ( .A1(n574), .A2(n573), .ZN(n602) );
  BUF_X1 U366 ( .A(n708), .Z(n342) );
  AND2_X1 U367 ( .A1(n539), .A2(n589), .ZN(n571) );
  NAND2_X1 U368 ( .A1(n538), .A2(n563), .ZN(n527) );
  NAND2_X1 U369 ( .A1(n561), .A2(n558), .ZN(n706) );
  OR2_X1 U370 ( .A1(n625), .A2(G902), .ZN(n407) );
  XNOR2_X1 U371 ( .A(n520), .B(n519), .ZN(n708) );
  XNOR2_X1 U372 ( .A(n348), .B(n343), .ZN(n445) );
  XNOR2_X1 U373 ( .A(n397), .B(KEYINPUT71), .ZN(n343) );
  NOR2_X2 U374 ( .A1(G953), .A2(G237), .ZN(n477) );
  XNOR2_X2 U375 ( .A(n442), .B(n441), .ZN(n745) );
  XNOR2_X2 U376 ( .A(KEYINPUT79), .B(KEYINPUT45), .ZN(n551) );
  AND2_X1 U377 ( .A1(n422), .A2(n421), .ZN(n420) );
  XNOR2_X2 U378 ( .A(n344), .B(KEYINPUT35), .ZN(n763) );
  NAND2_X2 U379 ( .A1(n390), .A2(n403), .ZN(n344) );
  NOR2_X2 U380 ( .A1(n706), .A2(n705), .ZN(n538) );
  XNOR2_X2 U381 ( .A(n655), .B(n657), .ZN(n658) );
  XNOR2_X2 U382 ( .A(n634), .B(KEYINPUT122), .ZN(n635) );
  XNOR2_X2 U383 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U384 ( .A(G116), .B(G107), .ZN(n488) );
  BUF_X1 U385 ( .A(G104), .Z(n663) );
  AND2_X2 U386 ( .A1(n375), .A2(n502), .ZN(n399) );
  AND2_X1 U387 ( .A1(n732), .A2(n347), .ZN(n346) );
  XNOR2_X1 U388 ( .A(n408), .B(G143), .ZN(n448) );
  INV_X1 U389 ( .A(G137), .ZN(n410) );
  INV_X1 U390 ( .A(G953), .ZN(n347) );
  XOR2_X1 U391 ( .A(G146), .B(G125), .Z(n482) );
  AND2_X1 U392 ( .A1(n733), .A2(n346), .ZN(n345) );
  NOR2_X1 U393 ( .A1(n728), .A2(n727), .ZN(n733) );
  XNOR2_X1 U394 ( .A(n689), .B(n688), .ZN(n691) );
  AND2_X1 U395 ( .A1(n415), .A2(n414), .ZN(n413) );
  AND2_X1 U396 ( .A1(n400), .A2(n388), .ZN(n386) );
  NOR2_X2 U397 ( .A1(n544), .A2(n543), .ZN(n677) );
  XNOR2_X1 U398 ( .A(n409), .B(n493), .ZN(n439) );
  XNOR2_X1 U399 ( .A(n448), .B(G134), .ZN(n493) );
  XNOR2_X1 U400 ( .A(n426), .B(n410), .ZN(n409) );
  INV_X1 U401 ( .A(KEYINPUT71), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n442), .B(n441), .ZN(n348) );
  NAND2_X1 U403 ( .A1(n745), .A2(KEYINPUT71), .ZN(n351) );
  NAND2_X1 U404 ( .A1(n349), .A2(n350), .ZN(n352) );
  NAND2_X1 U405 ( .A1(n352), .A2(n351), .ZN(n372) );
  INV_X1 U406 ( .A(n745), .ZN(n349) );
  BUF_X1 U407 ( .A(n354), .Z(n353) );
  AND2_X2 U408 ( .A1(n354), .A2(n690), .ZN(n371) );
  NAND2_X1 U409 ( .A1(n622), .A2(n621), .ZN(n354) );
  NAND2_X1 U410 ( .A1(n353), .A2(n355), .ZN(n629) );
  AND2_X1 U411 ( .A1(G469), .A2(n690), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n565), .B(KEYINPUT19), .ZN(n593) );
  XOR2_X1 U413 ( .A(G131), .B(G140), .Z(n471) );
  INV_X1 U414 ( .A(G224), .ZN(n361) );
  INV_X1 U415 ( .A(G128), .ZN(n408) );
  INV_X1 U416 ( .A(KEYINPUT22), .ZN(n416) );
  XNOR2_X1 U417 ( .A(G119), .B(G137), .ZN(n503) );
  XNOR2_X1 U418 ( .A(n492), .B(n491), .ZN(n378) );
  XOR2_X1 U419 ( .A(KEYINPUT97), .B(KEYINPUT7), .Z(n491) );
  INV_X1 U420 ( .A(G237), .ZN(n458) );
  AND2_X1 U421 ( .A1(n677), .A2(n584), .ZN(n562) );
  INV_X1 U422 ( .A(KEYINPUT0), .ZN(n373) );
  XNOR2_X1 U423 ( .A(KEYINPUT16), .B(G122), .ZN(n453) );
  XNOR2_X1 U424 ( .A(n380), .B(n379), .ZN(n509) );
  INV_X1 U425 ( .A(KEYINPUT8), .ZN(n379) );
  XNOR2_X1 U426 ( .A(n443), .B(n444), .ZN(n397) );
  AND2_X1 U427 ( .A1(n396), .A2(n606), .ZN(n395) );
  INV_X1 U428 ( .A(KEYINPUT15), .ZN(n456) );
  XNOR2_X1 U429 ( .A(G902), .B(KEYINPUT85), .ZN(n457) );
  XOR2_X1 U430 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n474) );
  XNOR2_X1 U431 ( .A(G113), .B(G143), .ZN(n472) );
  INV_X1 U432 ( .A(G146), .ZN(n444) );
  XNOR2_X1 U433 ( .A(n362), .B(n360), .ZN(n447) );
  XNOR2_X2 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n362) );
  NOR2_X2 U435 ( .A1(n361), .A2(G953), .ZN(n360) );
  AND2_X1 U436 ( .A1(G953), .A2(G902), .ZN(n466) );
  XNOR2_X1 U437 ( .A(n359), .B(KEYINPUT83), .ZN(n565) );
  NOR2_X1 U438 ( .A1(n500), .A2(n416), .ZN(n411) );
  NAND2_X1 U439 ( .A1(n500), .A2(n416), .ZN(n414) );
  INV_X1 U440 ( .A(G902), .ZN(n514) );
  INV_X1 U441 ( .A(G101), .ZN(n429) );
  XNOR2_X1 U442 ( .A(G113), .B(KEYINPUT70), .ZN(n434) );
  XNOR2_X1 U443 ( .A(G119), .B(G116), .ZN(n433) );
  XNOR2_X1 U444 ( .A(G110), .B(KEYINPUT76), .ZN(n505) );
  XNOR2_X1 U445 ( .A(n378), .B(n490), .ZN(n495) );
  INV_X1 U446 ( .A(n705), .ZN(n609) );
  NAND2_X1 U447 ( .A1(n461), .A2(G214), .ZN(n695) );
  OR2_X1 U448 ( .A1(n501), .A2(KEYINPUT65), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U450 ( .A(n581), .B(n580), .ZN(n767) );
  NAND2_X1 U451 ( .A1(n406), .A2(n405), .ZN(n403) );
  XNOR2_X1 U452 ( .A(n377), .B(n376), .ZN(n680) );
  INV_X1 U453 ( .A(KEYINPUT31), .ZN(n376) );
  AND2_X1 U454 ( .A1(n402), .A2(KEYINPUT100), .ZN(n356) );
  XOR2_X1 U455 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n357) );
  AND2_X1 U456 ( .A1(n404), .A2(n599), .ZN(n358) );
  NAND2_X1 U457 ( .A1(n575), .A2(n695), .ZN(n359) );
  XNOR2_X2 U458 ( .A(n460), .B(n459), .ZN(n575) );
  BUF_X1 U459 ( .A(n348), .Z(n363) );
  NAND2_X1 U460 ( .A1(n412), .A2(n411), .ZN(n375) );
  NAND2_X1 U461 ( .A1(n622), .A2(n621), .ZN(n364) );
  AND2_X2 U462 ( .A1(n367), .A2(n368), .ZN(n622) );
  NAND2_X2 U463 ( .A1(n624), .A2(KEYINPUT2), .ZN(n690) );
  BUF_X1 U464 ( .A(n387), .Z(n365) );
  NAND2_X1 U465 ( .A1(n365), .A2(n384), .ZN(n366) );
  NAND2_X1 U466 ( .A1(n387), .A2(n384), .ZN(n641) );
  NAND2_X1 U467 ( .A1(n623), .A2(n370), .ZN(n367) );
  OR2_X1 U468 ( .A1(n369), .A2(n687), .ZN(n368) );
  INV_X1 U469 ( .A(n618), .ZN(n369) );
  AND2_X1 U470 ( .A1(KEYINPUT78), .A2(n618), .ZN(n370) );
  AND2_X2 U471 ( .A1(n364), .A2(n690), .ZN(n734) );
  NAND2_X1 U472 ( .A1(n763), .A2(KEYINPUT44), .ZN(n417) );
  AND2_X1 U473 ( .A1(n401), .A2(n342), .ZN(n400) );
  XNOR2_X2 U474 ( .A(n374), .B(n373), .ZN(n528) );
  NOR2_X2 U475 ( .A1(n593), .A2(n470), .ZN(n374) );
  NAND2_X1 U476 ( .A1(n413), .A2(n375), .ZN(n534) );
  NOR2_X1 U477 ( .A1(n529), .A2(n717), .ZN(n377) );
  XNOR2_X1 U478 ( .A(n393), .B(KEYINPUT48), .ZN(n615) );
  NAND2_X1 U479 ( .A1(n347), .A2(G234), .ZN(n380) );
  XNOR2_X2 U480 ( .A(n525), .B(n524), .ZN(n769) );
  NAND2_X1 U481 ( .A1(n419), .A2(KEYINPUT44), .ZN(n418) );
  AND2_X2 U482 ( .A1(n382), .A2(n381), .ZN(n387) );
  NAND2_X1 U483 ( .A1(n534), .A2(n402), .ZN(n389) );
  NAND2_X1 U484 ( .A1(n534), .A2(n356), .ZN(n381) );
  NAND2_X1 U485 ( .A1(n383), .A2(KEYINPUT100), .ZN(n382) );
  NAND2_X1 U486 ( .A1(n398), .A2(n400), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n389), .A2(n385), .ZN(n384) );
  AND2_X1 U488 ( .A1(n398), .A2(n386), .ZN(n385) );
  INV_X1 U489 ( .A(KEYINPUT100), .ZN(n388) );
  NAND2_X1 U490 ( .A1(n641), .A2(n769), .ZN(n526) );
  INV_X1 U491 ( .A(n391), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n358), .A2(n392), .ZN(n391) );
  NAND2_X1 U493 ( .A1(n529), .A2(n530), .ZN(n392) );
  NAND2_X1 U494 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U495 ( .A(n592), .B(KEYINPUT46), .ZN(n394) );
  INV_X1 U496 ( .A(n683), .ZN(n396) );
  NAND2_X1 U497 ( .A1(n399), .A2(n413), .ZN(n398) );
  AND2_X1 U498 ( .A1(n501), .A2(KEYINPUT65), .ZN(n402) );
  NAND2_X1 U499 ( .A1(n730), .A2(n530), .ZN(n404) );
  NOR2_X1 U500 ( .A1(n529), .A2(n530), .ZN(n405) );
  INV_X1 U501 ( .A(n730), .ZN(n406) );
  XNOR2_X2 U502 ( .A(n527), .B(n425), .ZN(n730) );
  XNOR2_X2 U503 ( .A(n589), .B(n357), .ZN(n705) );
  XNOR2_X2 U504 ( .A(n407), .B(G469), .ZN(n589) );
  INV_X1 U505 ( .A(n528), .ZN(n412) );
  NAND2_X1 U506 ( .A1(n528), .A2(n416), .ZN(n415) );
  XNOR2_X1 U507 ( .A(n526), .B(KEYINPUT81), .ZN(n424) );
  AND2_X1 U508 ( .A1(n550), .A2(n417), .ZN(n421) );
  INV_X1 U509 ( .A(n424), .ZN(n419) );
  NAND2_X1 U510 ( .A1(n420), .A2(n418), .ZN(n552) );
  NAND2_X1 U511 ( .A1(n424), .A2(n423), .ZN(n422) );
  AND2_X1 U512 ( .A1(n532), .A2(n533), .ZN(n423) );
  XNOR2_X2 U513 ( .A(n440), .B(G110), .ZN(n442) );
  XNOR2_X1 U514 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n425) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n617) );
  XNOR2_X1 U516 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U517 ( .A(KEYINPUT77), .ZN(n688) );
  XNOR2_X1 U518 ( .A(n432), .B(n431), .ZN(n436) );
  INV_X1 U519 ( .A(KEYINPUT65), .ZN(n502) );
  INV_X1 U520 ( .A(n493), .ZN(n494) );
  NAND2_X1 U521 ( .A1(n691), .A2(n690), .ZN(n694) );
  BUF_X1 U522 ( .A(n692), .Z(n754) );
  XNOR2_X1 U523 ( .A(KEYINPUT36), .B(KEYINPUT82), .ZN(n568) );
  XNOR2_X1 U524 ( .A(n569), .B(n568), .ZN(n570) );
  INV_X1 U525 ( .A(KEYINPUT40), .ZN(n580) );
  INV_X1 U526 ( .A(KEYINPUT123), .ZN(n638) );
  XOR2_X1 U527 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n446) );
  INV_X1 U528 ( .A(n446), .ZN(n426) );
  XOR2_X1 U529 ( .A(KEYINPUT93), .B(G131), .Z(n428) );
  NAND2_X1 U530 ( .A1(n477), .A2(G210), .ZN(n427) );
  XNOR2_X1 U531 ( .A(n428), .B(n427), .ZN(n432) );
  XNOR2_X1 U532 ( .A(G146), .B(KEYINPUT5), .ZN(n430) );
  XNOR2_X1 U533 ( .A(n433), .B(KEYINPUT3), .ZN(n435) );
  XNOR2_X1 U534 ( .A(n435), .B(n434), .ZN(n454) );
  XNOR2_X1 U535 ( .A(n436), .B(n454), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n439), .B(n437), .ZN(n642) );
  NAND2_X1 U537 ( .A1(n642), .A2(n514), .ZN(n438) );
  XNOR2_X2 U538 ( .A(n438), .B(G472), .ZN(n712) );
  INV_X1 U539 ( .A(n712), .ZN(n540) );
  XNOR2_X1 U540 ( .A(n439), .B(n471), .ZN(n752) );
  XNOR2_X2 U541 ( .A(G107), .B(G104), .ZN(n440) );
  XNOR2_X1 U542 ( .A(G101), .B(KEYINPUT86), .ZN(n441) );
  NAND2_X1 U543 ( .A1(G227), .A2(n347), .ZN(n443) );
  XNOR2_X1 U544 ( .A(n752), .B(n445), .ZN(n625) );
  AND2_X1 U545 ( .A1(n540), .A2(n705), .ZN(n501) );
  XNOR2_X1 U546 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n448), .B(n482), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n372), .B(n451), .ZN(n455) );
  XNOR2_X1 U549 ( .A(n454), .B(n453), .ZN(n746) );
  XNOR2_X1 U550 ( .A(n455), .B(n746), .ZN(n654) );
  NAND2_X1 U551 ( .A1(n654), .A2(n617), .ZN(n460) );
  NAND2_X1 U552 ( .A1(n514), .A2(n458), .ZN(n461) );
  AND2_X1 U553 ( .A1(n461), .A2(G210), .ZN(n459) );
  NAND2_X1 U554 ( .A1(G234), .A2(G237), .ZN(n462) );
  XNOR2_X1 U555 ( .A(n462), .B(KEYINPUT14), .ZN(n467) );
  NAND2_X1 U556 ( .A1(n467), .A2(G952), .ZN(n463) );
  XOR2_X1 U557 ( .A(KEYINPUT87), .B(n463), .Z(n726) );
  NOR2_X1 U558 ( .A1(n726), .A2(G953), .ZN(n465) );
  INV_X1 U559 ( .A(KEYINPUT88), .ZN(n464) );
  XNOR2_X1 U560 ( .A(n465), .B(n464), .ZN(n557) );
  NAND2_X1 U561 ( .A1(n467), .A2(n466), .ZN(n553) );
  NOR2_X1 U562 ( .A1(G898), .A2(n553), .ZN(n468) );
  XNOR2_X1 U563 ( .A(n468), .B(KEYINPUT89), .ZN(n469) );
  AND2_X1 U564 ( .A1(n557), .A2(n469), .ZN(n470) );
  XNOR2_X1 U565 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U566 ( .A(n663), .B(G122), .ZN(n473) );
  XNOR2_X1 U567 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U568 ( .A(n476), .B(n475), .ZN(n481) );
  XOR2_X1 U569 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n479) );
  NAND2_X1 U570 ( .A1(G214), .A2(n477), .ZN(n478) );
  XNOR2_X1 U571 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n481), .B(n480), .ZN(n484) );
  XNOR2_X1 U573 ( .A(n482), .B(KEYINPUT10), .ZN(n483) );
  XNOR2_X1 U574 ( .A(n483), .B(KEYINPUT68), .ZN(n751) );
  XNOR2_X1 U575 ( .A(n484), .B(n751), .ZN(n647) );
  NOR2_X1 U576 ( .A1(G902), .A2(n647), .ZN(n486) );
  XNOR2_X1 U577 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n487), .B(G475), .ZN(n545) );
  XOR2_X1 U580 ( .A(KEYINPUT9), .B(G122), .Z(n489) );
  XNOR2_X1 U581 ( .A(n489), .B(n488), .ZN(n492) );
  NAND2_X1 U582 ( .A1(G217), .A2(n509), .ZN(n490) );
  XOR2_X1 U583 ( .A(n495), .B(n494), .Z(n634) );
  NOR2_X1 U584 ( .A1(n634), .A2(G902), .ZN(n496) );
  XNOR2_X1 U585 ( .A(n496), .B(G478), .ZN(n546) );
  INV_X1 U586 ( .A(n546), .ZN(n543) );
  OR2_X1 U587 ( .A1(n545), .A2(n543), .ZN(n698) );
  NAND2_X1 U588 ( .A1(n617), .A2(G234), .ZN(n497) );
  XNOR2_X1 U589 ( .A(n497), .B(KEYINPUT20), .ZN(n515) );
  AND2_X1 U590 ( .A1(n515), .A2(G221), .ZN(n499) );
  XNOR2_X1 U591 ( .A(KEYINPUT92), .B(KEYINPUT21), .ZN(n498) );
  XNOR2_X1 U592 ( .A(n499), .B(n498), .ZN(n558) );
  INV_X1 U593 ( .A(n558), .ZN(n709) );
  OR2_X1 U594 ( .A1(n698), .A2(n709), .ZN(n500) );
  INV_X1 U595 ( .A(n751), .ZN(n513) );
  XOR2_X1 U596 ( .A(G140), .B(G128), .Z(n504) );
  XNOR2_X1 U597 ( .A(n504), .B(n503), .ZN(n508) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n506) );
  XNOR2_X1 U599 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U600 ( .A(n508), .B(n507), .Z(n511) );
  NAND2_X1 U601 ( .A1(G221), .A2(n509), .ZN(n510) );
  XNOR2_X1 U602 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U603 ( .A(n512), .B(n513), .ZN(n736) );
  NAND2_X1 U604 ( .A1(n736), .A2(n514), .ZN(n520) );
  XOR2_X1 U605 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n517) );
  NAND2_X1 U606 ( .A1(n515), .A2(G217), .ZN(n516) );
  XNOR2_X1 U607 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n518), .B(KEYINPUT90), .ZN(n519) );
  XOR2_X1 U609 ( .A(n712), .B(KEYINPUT6), .Z(n563) );
  XOR2_X1 U610 ( .A(KEYINPUT74), .B(n563), .Z(n521) );
  NAND2_X1 U611 ( .A1(n521), .A2(n342), .ZN(n522) );
  NOR2_X1 U612 ( .A1(n705), .A2(n522), .ZN(n523) );
  NAND2_X1 U613 ( .A1(n534), .A2(n523), .ZN(n525) );
  XOR2_X1 U614 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n524) );
  INV_X1 U615 ( .A(n708), .ZN(n561) );
  BUF_X1 U616 ( .A(n528), .Z(n529) );
  XNOR2_X1 U617 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n530) );
  AND2_X1 U618 ( .A1(n545), .A2(n543), .ZN(n599) );
  INV_X1 U619 ( .A(n763), .ZN(n532) );
  INV_X1 U620 ( .A(KEYINPUT44), .ZN(n533) );
  AND2_X1 U621 ( .A1(n534), .A2(n705), .ZN(n536) );
  NOR2_X1 U622 ( .A1(n563), .A2(n342), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U624 ( .A(n537), .B(KEYINPUT99), .ZN(n764) );
  NAND2_X1 U625 ( .A1(n712), .A2(n538), .ZN(n717) );
  INV_X1 U626 ( .A(n706), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n571), .A2(n540), .ZN(n541) );
  OR2_X1 U628 ( .A1(n529), .A2(n541), .ZN(n542) );
  INV_X1 U629 ( .A(n542), .ZN(n665) );
  NOR2_X1 U630 ( .A1(n680), .A2(n665), .ZN(n548) );
  INV_X1 U631 ( .A(n545), .ZN(n544) );
  NOR2_X1 U632 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U633 ( .A(KEYINPUT98), .B(n547), .ZN(n681) );
  NOR2_X1 U634 ( .A1(n677), .A2(n681), .ZN(n701) );
  NOR2_X1 U635 ( .A1(n548), .A2(n701), .ZN(n549) );
  NOR2_X1 U636 ( .A1(n764), .A2(n549), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n552), .B(n551), .ZN(n686) );
  XNOR2_X1 U638 ( .A(n553), .B(KEYINPUT102), .ZN(n554) );
  NOR2_X1 U639 ( .A1(G900), .A2(n554), .ZN(n555) );
  XNOR2_X1 U640 ( .A(KEYINPUT103), .B(n555), .ZN(n556) );
  NAND2_X1 U641 ( .A1(n557), .A2(n556), .ZN(n598) );
  NAND2_X1 U642 ( .A1(n558), .A2(n598), .ZN(n559) );
  XOR2_X1 U643 ( .A(KEYINPUT69), .B(n559), .Z(n560) );
  NOR2_X1 U644 ( .A1(n561), .A2(n560), .ZN(n584) );
  NAND2_X1 U645 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U646 ( .A(KEYINPUT104), .B(n564), .ZN(n608) );
  INV_X1 U647 ( .A(n608), .ZN(n567) );
  BUF_X1 U648 ( .A(n565), .Z(n566) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n569) );
  NOR2_X1 U650 ( .A1(n705), .A2(n570), .ZN(n683) );
  XNOR2_X1 U651 ( .A(KEYINPUT105), .B(n571), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n695), .A2(n712), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n572), .B(KEYINPUT30), .ZN(n573) );
  BUF_X1 U654 ( .A(n575), .Z(n576) );
  XNOR2_X1 U655 ( .A(n576), .B(KEYINPUT38), .ZN(n582) );
  INV_X1 U656 ( .A(n598), .ZN(n577) );
  NOR2_X1 U657 ( .A1(n582), .A2(n577), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n602), .A2(n578), .ZN(n579) );
  NAND2_X1 U659 ( .A1(n677), .A2(n607), .ZN(n581) );
  INV_X1 U660 ( .A(n582), .ZN(n696) );
  NAND2_X1 U661 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U662 ( .A1(n698), .A2(n700), .ZN(n583) );
  XNOR2_X1 U663 ( .A(KEYINPUT41), .B(n583), .ZN(n729) );
  AND2_X1 U664 ( .A1(n712), .A2(n584), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n585) );
  XNOR2_X1 U666 ( .A(KEYINPUT28), .B(n585), .ZN(n586) );
  XNOR2_X1 U667 ( .A(n587), .B(n586), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U669 ( .A(KEYINPUT109), .B(n590), .Z(n595) );
  NOR2_X1 U670 ( .A1(n729), .A2(n595), .ZN(n591) );
  XNOR2_X1 U671 ( .A(n591), .B(KEYINPUT42), .ZN(n765) );
  BUF_X1 U672 ( .A(n593), .Z(n594) );
  NOR2_X1 U673 ( .A1(KEYINPUT67), .A2(n701), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n673), .A2(n596), .ZN(n597) );
  XNOR2_X1 U675 ( .A(KEYINPUT47), .B(n597), .ZN(n605) );
  AND2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  AND2_X1 U677 ( .A1(n576), .A2(n600), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT106), .B(n603), .ZN(n768) );
  XNOR2_X1 U680 ( .A(KEYINPUT75), .B(n768), .ZN(n604) );
  NOR2_X1 U681 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n681), .ZN(n685) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n610), .A2(n695), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(KEYINPUT43), .ZN(n613) );
  INV_X1 U686 ( .A(n576), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n640) );
  NAND2_X1 U688 ( .A1(n685), .A2(n640), .ZN(n614) );
  NOR2_X2 U689 ( .A1(n615), .A2(n614), .ZN(n692) );
  INV_X1 U690 ( .A(n692), .ZN(n616) );
  NOR2_X2 U691 ( .A1(n686), .A2(n616), .ZN(n623) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n687) );
  INV_X1 U693 ( .A(n617), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n623), .A2(n618), .ZN(n620) );
  INV_X1 U695 ( .A(KEYINPUT78), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  BUF_X1 U697 ( .A(n623), .Z(n624) );
  XOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n627) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT120), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U701 ( .A(G952), .ZN(n630) );
  AND2_X1 U702 ( .A1(n630), .A2(G953), .ZN(n738) );
  NOR2_X2 U703 ( .A1(n631), .A2(n738), .ZN(n633) );
  INV_X1 U704 ( .A(KEYINPUT121), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n633), .B(n632), .ZN(G54) );
  NAND2_X1 U706 ( .A1(n734), .A2(G478), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X2 U708 ( .A1(n637), .A2(n738), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(G63) );
  XNOR2_X1 U710 ( .A(n640), .B(G140), .ZN(G42) );
  XNOR2_X1 U711 ( .A(n366), .B(G110), .ZN(G12) );
  NAND2_X1 U712 ( .A1(n371), .A2(G472), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n642), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(n645) );
  INV_X1 U715 ( .A(n738), .ZN(n650) );
  NAND2_X1 U716 ( .A1(n645), .A2(n650), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U718 ( .A1(n371), .A2(G475), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT59), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n653) );
  INV_X1 U722 ( .A(KEYINPUT60), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G60) );
  NAND2_X1 U724 ( .A1(n734), .A2(G210), .ZN(n659) );
  BUF_X1 U725 ( .A(n654), .Z(n655) );
  XNOR2_X1 U726 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(KEYINPUT55), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X2 U729 ( .A1(n660), .A2(n738), .ZN(n662) );
  XNOR2_X1 U730 ( .A(KEYINPUT80), .B(KEYINPUT56), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n662), .B(n661), .ZN(G51) );
  NAND2_X1 U732 ( .A1(n665), .A2(n677), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(G6) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT110), .ZN(n669) );
  XOR2_X1 U735 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n667) );
  NAND2_X1 U736 ( .A1(n665), .A2(n681), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(G9) );
  XOR2_X1 U739 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n671) );
  NAND2_X1 U740 ( .A1(n673), .A2(n681), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U742 ( .A(G128), .B(n672), .Z(G30) );
  XOR2_X1 U743 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n675) );
  NAND2_X1 U744 ( .A1(n673), .A2(n677), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U746 ( .A(G146), .B(n676), .ZN(G48) );
  NAND2_X1 U747 ( .A1(n680), .A2(n677), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n678), .B(KEYINPUT114), .ZN(n679) );
  XNOR2_X1 U749 ( .A(G113), .B(n679), .ZN(G15) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U751 ( .A(n682), .B(G116), .ZN(G18) );
  XNOR2_X1 U752 ( .A(G125), .B(n683), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n684), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U754 ( .A(G134), .B(n685), .ZN(G36) );
  BUF_X1 U755 ( .A(n686), .Z(n739) );
  NAND2_X1 U756 ( .A1(n739), .A2(n687), .ZN(n689) );
  NOR2_X1 U757 ( .A1(KEYINPUT2), .A2(n754), .ZN(n693) );
  NOR2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n728) );
  NOR2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT117), .B(n699), .Z(n703) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U763 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n730), .A2(n704), .ZN(n722) );
  XNOR2_X1 U765 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n719) );
  NAND2_X1 U766 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U767 ( .A(KEYINPUT50), .B(n707), .ZN(n715) );
  XOR2_X1 U768 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n711) );
  NAND2_X1 U769 ( .A1(n709), .A2(n342), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U772 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U775 ( .A1(n720), .A2(n729), .ZN(n721) );
  NOR2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(KEYINPUT118), .ZN(n724) );
  XNOR2_X1 U778 ( .A(KEYINPUT52), .B(n724), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT119), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n345), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U783 ( .A1(n371), .A2(G217), .ZN(n735) );
  XOR2_X1 U784 ( .A(n736), .B(n735), .Z(n737) );
  NOR2_X1 U785 ( .A1(n738), .A2(n737), .ZN(G66) );
  INV_X1 U786 ( .A(n739), .ZN(n740) );
  NAND2_X1 U787 ( .A1(n740), .A2(n347), .ZN(n744) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n741) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n741), .ZN(n742) );
  NAND2_X1 U790 ( .A1(n742), .A2(G898), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n744), .A2(n743), .ZN(n750) );
  XNOR2_X1 U792 ( .A(n363), .B(n746), .ZN(n748) );
  NOR2_X1 U793 ( .A1(G898), .A2(n347), .ZN(n747) );
  NOR2_X1 U794 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U795 ( .A(n750), .B(n749), .ZN(G69) );
  XNOR2_X1 U796 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U797 ( .A(n753), .B(KEYINPUT124), .Z(n756) );
  XOR2_X1 U798 ( .A(n756), .B(n754), .Z(n755) );
  NOR2_X1 U799 ( .A1(G953), .A2(n755), .ZN(n761) );
  XNOR2_X1 U800 ( .A(KEYINPUT125), .B(n756), .ZN(n757) );
  XNOR2_X1 U801 ( .A(G227), .B(n757), .ZN(n759) );
  NAND2_X1 U802 ( .A1(G900), .A2(G953), .ZN(n758) );
  NOR2_X1 U803 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U804 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U805 ( .A(KEYINPUT126), .B(n762), .ZN(G72) );
  XOR2_X1 U806 ( .A(n763), .B(G122), .Z(G24) );
  XOR2_X1 U807 ( .A(G101), .B(n764), .Z(G3) );
  XNOR2_X1 U808 ( .A(G137), .B(KEYINPUT127), .ZN(n766) );
  XNOR2_X1 U809 ( .A(n766), .B(n765), .ZN(G39) );
  XOR2_X1 U810 ( .A(n767), .B(G131), .Z(G33) );
  XNOR2_X1 U811 ( .A(G143), .B(n768), .ZN(G45) );
  XNOR2_X1 U812 ( .A(n769), .B(G119), .ZN(G21) );
endmodule

