//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(G2104), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR3_X1   g038(.A1(new_n463), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n464));
  OAI21_X1  g039(.A(G101), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n461), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n461), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n477), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G138), .B(new_n461), .C1(new_n470), .C2(new_n471), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n466), .A2(new_n488), .A3(G138), .A4(new_n461), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n461), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n480), .A2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n490), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT68), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n505), .B2(new_n507), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(KEYINPUT69), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n518), .B1(new_n516), .B2(KEYINPUT69), .ZN(new_n519));
  OAI21_X1  g094(.A(G651), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g097(.A(KEYINPUT70), .B(G651), .C1(new_n517), .C2(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n526), .B(new_n530), .C1(new_n531), .C2(new_n512), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n508), .A2(G89), .A3(new_n509), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n510), .A2(new_n538), .B1(new_n512), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(new_n510), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT71), .B(G81), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n509), .A2(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n536), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n505), .B2(new_n507), .ZN(new_n557));
  AND2_X1   g132(.A1(G78), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g136(.A(KEYINPUT73), .B(G651), .C1(new_n557), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n512), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n508), .A2(G91), .A3(new_n509), .ZN(new_n567));
  XOR2_X1   g142(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n568));
  NAND4_X1  g143(.A1(new_n568), .A2(G53), .A3(G543), .A4(new_n509), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n563), .A2(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(new_n542), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n545), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n510), .A2(new_n578), .B1(new_n512), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n508), .A2(G61), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT74), .B1(new_n584), .B2(G651), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n505), .B2(new_n507), .ZN(new_n587));
  INV_X1    g162(.A(new_n583), .ZN(new_n588));
  OAI211_X1 g163(.A(KEYINPUT74), .B(G651), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n581), .B1(new_n585), .B2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n536), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n545), .A2(G47), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n508), .A2(G85), .A3(new_n509), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT75), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n594), .B1(new_n597), .B2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n542), .A2(new_n601), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT76), .B1(new_n510), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n604), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n508), .A2(G66), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT77), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(KEYINPUT77), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(G54), .B2(new_n545), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G286), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G299), .B(KEYINPUT78), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G297));
  AOI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g204(.A1(new_n462), .A2(new_n464), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n466), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(KEYINPUT79), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(KEYINPUT79), .B2(new_n637), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n480), .A2(G123), .ZN(new_n641));
  INV_X1    g216(.A(G135), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n467), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n635), .A2(new_n636), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(G14), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(G401));
  XOR2_X1   g236(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n662), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(new_n684), .B(new_n683), .S(new_n676), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT82), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  NAND2_X1  g268(.A1(G160), .A2(G29), .ZN(new_n694));
  INV_X1    g269(.A(G34), .ZN(new_n695));
  AOI21_X1  g270(.A(G29), .B1(new_n695), .B2(KEYINPUT24), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(KEYINPUT24), .B2(new_n695), .ZN(new_n697));
  AOI21_X1  g272(.A(G2084), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G33), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT25), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n476), .A2(G139), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n466), .A2(G127), .ZN(new_n706));
  NAND2_X1  g281(.A1(G115), .A2(G2104), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(G2105), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n700), .B1(new_n711), .B2(new_n699), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n698), .B1(G2072), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n694), .A2(G2084), .A3(new_n697), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n713), .B(new_n714), .C1(G2072), .C2(new_n712), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n699), .A2(G32), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n476), .A2(G141), .B1(G129), .B2(new_n480), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n630), .A2(G105), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n699), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT27), .B(G1996), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G29), .A2(G35), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G162), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT29), .B(G2090), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n715), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n732), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n732), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n735), .B1(G1961), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT30), .B(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n699), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n699), .B2(new_n643), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n734), .B2(G1966), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT94), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G16), .A2(G19), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n550), .B2(G16), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1341), .Z(new_n750));
  AND3_X1   g325(.A1(new_n731), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n616), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G4), .B2(G16), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT90), .B(G1348), .Z(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT89), .Z(new_n755));
  AND2_X1   g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n745), .A2(new_n746), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n753), .A2(new_n755), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n732), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  INV_X1    g336(.A(G299), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n732), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT95), .B(G1956), .Z(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n480), .A2(G128), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n461), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G140), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n769), .B2(new_n770), .C1(new_n771), .C2(new_n467), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n767), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(G164), .A2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G27), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n737), .A2(G1961), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n763), .A2(new_n764), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n765), .A2(new_n776), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n751), .A2(new_n759), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G290), .A2(new_n732), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G24), .ZN(new_n788));
  INV_X1    g363(.A(G1986), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g365(.A1(G95), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT83), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n476), .A2(G131), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n480), .A2(G119), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G29), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G25), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT84), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n801), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n798), .B(new_n803), .C1(G25), .C2(G29), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n787), .B(G1986), .C1(G16), .C2(G24), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n790), .A2(new_n805), .A3(KEYINPUT88), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(G16), .A2(G22), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G303), .B2(new_n732), .ZN(new_n809));
  INV_X1    g384(.A(G1971), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n732), .A2(G23), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G288), .B2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT33), .B(G1976), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n732), .A2(G6), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT74), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n587), .A2(new_n588), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n536), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n580), .B1(new_n820), .B2(new_n589), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n817), .B1(new_n821), .B2(new_n732), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT32), .B(G1981), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT86), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT85), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n816), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n809), .A2(new_n810), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n812), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT34), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n807), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n816), .A2(new_n826), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n809), .A2(new_n810), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n834), .A3(new_n811), .A4(new_n827), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n835), .A2(KEYINPUT87), .A3(KEYINPUT34), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT87), .B1(new_n835), .B2(KEYINPUT34), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(new_n832), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n786), .B1(new_n839), .B2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n786), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT96), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n846));
  AOI211_X1 g421(.A(new_n846), .B(new_n786), .C1(new_n839), .C2(new_n841), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n845), .A2(new_n847), .ZN(G150));
  NAND2_X1  g423(.A1(new_n542), .A2(G93), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT97), .B(G55), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n545), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n536), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT98), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n856), .A2(new_n857), .A3(new_n849), .A4(new_n851), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n544), .B(new_n546), .C1(new_n536), .C2(new_n548), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n852), .A2(new_n854), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n550), .A2(new_n861), .A3(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT38), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n615), .A2(new_n624), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AOI21_X1  g442(.A(G860), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n867), .B2(new_n866), .ZN(new_n869));
  INV_X1    g444(.A(new_n861), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(G145));
  XOR2_X1   g448(.A(KEYINPUT101), .B(G37), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G164), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n774), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n772), .B(KEYINPUT91), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(G164), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n877), .A2(new_n879), .A3(new_n722), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n722), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n710), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n877), .A2(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n723), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n879), .A3(new_n722), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n711), .A3(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n797), .A2(new_n632), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n480), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n461), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G142), .ZN(new_n892));
  OR3_X1    g467(.A1(new_n467), .A2(KEYINPUT99), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT99), .B1(new_n467), .B2(new_n892), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n797), .A2(new_n632), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n887), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n887), .B2(new_n896), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n882), .A2(new_n886), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n882), .A2(new_n886), .ZN(new_n902));
  INV_X1    g477(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g479(.A(KEYINPUT100), .B(new_n899), .C1(new_n882), .C2(new_n886), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n484), .B(G160), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(new_n643), .Z(new_n908));
  AOI21_X1  g483(.A(new_n875), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n900), .B2(new_n910), .ZN(new_n911));
  OAI221_X1 g486(.A(new_n911), .B1(new_n910), .B2(new_n900), .C1(new_n904), .C2(new_n905), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT40), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(new_n870), .A2(new_n619), .ZN(new_n916));
  NOR2_X1   g491(.A1(G303), .A2(new_n821), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G290), .B(G288), .ZN(new_n919));
  AOI21_X1  g494(.A(G305), .B1(new_n522), .B2(new_n523), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G288), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n917), .B2(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT103), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  MUX2_X1   g505(.A(new_n926), .B(new_n930), .S(KEYINPUT42), .Z(new_n931));
  XNOR2_X1  g506(.A(new_n626), .B(new_n863), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n615), .A2(G299), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n615), .A2(G299), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT41), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n616), .A2(new_n762), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n615), .A2(G299), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n935), .B1(new_n932), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n931), .B(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n916), .B1(new_n943), .B2(new_n619), .ZN(G295));
  OAI21_X1  g519(.A(new_n916), .B1(new_n943), .B2(new_n619), .ZN(G331));
  OAI21_X1  g520(.A(KEYINPUT104), .B1(new_n532), .B2(new_n533), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n545), .A2(G51), .B1(new_n529), .B2(new_n528), .ZN(new_n947));
  INV_X1    g522(.A(new_n533), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .A4(new_n526), .ZN(new_n950));
  NAND3_X1  g525(.A1(G301), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(G168), .A2(G171), .A3(new_n949), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n863), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n860), .A2(new_n862), .A3(new_n952), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n937), .A3(new_n940), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n939), .A3(new_n938), .A4(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT103), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n922), .B2(new_n925), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n928), .A2(new_n929), .A3(new_n957), .A4(new_n958), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n957), .A2(new_n958), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n875), .B1(new_n930), .B2(new_n959), .ZN(new_n969));
  AOI22_X1  g544(.A1(KEYINPUT43), .A2(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n970), .B2(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n968), .A2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n930), .B2(new_n959), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n963), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n968), .B2(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n962), .A2(new_n963), .A3(new_n874), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n979), .A2(KEYINPUT106), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT106), .B1(new_n979), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n971), .B(new_n978), .C1(new_n982), .C2(new_n983), .ZN(G397));
  INV_X1    g559(.A(G1384), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n490), .B2(new_n501), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  INV_X1    g562(.A(G40), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n469), .A2(new_n988), .A3(new_n474), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n774), .A2(G2067), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n878), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT108), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n796), .B(new_n800), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n991), .A2(new_n722), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n990), .A2(G1996), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n1000), .A2(new_n1001), .B1(G1996), .B2(new_n723), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT127), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT127), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n997), .A2(new_n1005), .A3(new_n999), .A4(new_n1002), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n990), .A2(G290), .A3(G1986), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n997), .A2(new_n1002), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n797), .A2(new_n800), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n994), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n991), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n996), .A2(new_n1000), .A3(KEYINPUT125), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT125), .B1(new_n996), .B2(new_n1000), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT124), .B(KEYINPUT46), .Z(new_n1016));
  NOR2_X1   g591(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1017));
  MUX2_X1   g592(.A(new_n1016), .B(new_n1017), .S(new_n1001), .Z(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1020), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1009), .A2(new_n1013), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n494), .A2(new_n498), .B1(new_n480), .B2(G126), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n487), .A2(new_n489), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n989), .A2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT111), .B(G8), .Z(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1030), .B(new_n1032), .C1(new_n1033), .C2(G288), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1035), .A2(KEYINPUT112), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G288), .A2(new_n1035), .A3(new_n1033), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n821), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(KEYINPUT49), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .A4(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n476), .A2(G137), .ZN(new_n1048));
  INV_X1    g623(.A(new_n474), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(G40), .A4(new_n465), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n986), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n1031), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1047), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n821), .A2(new_n1042), .ZN(new_n1054));
  AOI211_X1 g629(.A(G1981), .B(new_n580), .C1(new_n820), .C2(new_n589), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT113), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1041), .A2(new_n1057), .A3(new_n1043), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1040), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n522), .B2(new_n523), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT110), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n986), .A2(new_n987), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n989), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n810), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1050), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1029), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1029), .B2(new_n1075), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1073), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1072), .B1(new_n1079), .B2(G2090), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1068), .B1(G8), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1026), .B1(new_n1061), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1068), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(new_n1047), .A3(new_n1045), .A4(new_n1052), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1085), .A2(KEYINPUT117), .A3(new_n1087), .A4(new_n1040), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1073), .B(new_n1089), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1090));
  INV_X1    g665(.A(G1966), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1071), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1032), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(G286), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1082), .A2(new_n1088), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT63), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1029), .A2(new_n1075), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1073), .A2(KEYINPUT115), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n989), .B1(new_n1029), .B2(new_n1075), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT50), .B(G1384), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G2090), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1031), .B1(new_n1106), .B2(new_n1072), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(new_n1068), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1094), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1109), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1087), .A2(new_n1033), .A3(new_n923), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1043), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1061), .A2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1052), .B1(new_n1117), .B2(new_n1098), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1097), .A2(new_n1113), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G168), .A2(new_n1031), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1094), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1062), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT51), .B1(new_n1123), .B2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1093), .A2(G286), .A3(new_n1032), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1122), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n989), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n987), .B(G1384), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1131), .A2(G2078), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1069), .A2(new_n779), .A3(new_n989), .A4(new_n1070), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT121), .ZN(new_n1137));
  INV_X1    g712(.A(G1961), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1135), .A2(new_n1137), .B1(new_n1138), .B2(new_n1079), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1136), .B2(new_n1130), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1136), .A2(new_n1140), .A3(new_n1130), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(G301), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(KEYINPUT62), .B(new_n1122), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1129), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1079), .A2(new_n1138), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1133), .A2(KEYINPUT53), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1136), .A2(new_n1140), .A3(new_n1130), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1149), .B(new_n1150), .C1(new_n1151), .C2(new_n1141), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1148), .B1(new_n1152), .B2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1139), .A2(new_n1144), .A3(G301), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1153), .A2(KEYINPUT123), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT123), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G1956), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT56), .B(G2072), .Z(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1069), .A2(new_n989), .A3(new_n1070), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n1163));
  NAND3_X1  g738(.A1(G299), .A2(new_n1163), .A3(KEYINPUT57), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1163), .A2(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(KEYINPUT57), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n563), .A2(new_n570), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1159), .A2(new_n1162), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  AND4_X1   g743(.A1(new_n1159), .A2(new_n1162), .A3(new_n1167), .A4(new_n1164), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n615), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1079), .A2(new_n754), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1051), .A2(new_n993), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1168), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1131), .A2(G1996), .A3(new_n1132), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT58), .B(G1341), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1051), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n550), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n550), .B(new_n1179), .C1(new_n1175), .C2(new_n1177), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1159), .A2(new_n1162), .A3(new_n1167), .A4(new_n1164), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1188), .A2(KEYINPUT61), .A3(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1183), .A2(new_n1185), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT60), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1099), .A2(KEYINPUT109), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1102), .B1(new_n1193), .B2(new_n1076), .ZN(new_n1194));
  INV_X1    g769(.A(new_n754), .ZN(new_n1195));
  OAI211_X1 g770(.A(KEYINPUT60), .B(new_n1172), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n616), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n615), .A4(new_n1172), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1192), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1174), .B1(new_n1191), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(G301), .B1(new_n1151), .B2(new_n1141), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1148), .B1(new_n1145), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1127), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1200), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1147), .B1(new_n1157), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1208), .A2(new_n1098), .A3(new_n1108), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1119), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(G290), .B(new_n789), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1211), .A2(new_n990), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n1003), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1025), .B1(new_n1210), .B2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n909), .A2(new_n912), .ZN(new_n1216));
  NOR4_X1   g790(.A1(G229), .A2(G401), .A3(new_n458), .A4(G227), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1218), .A2(new_n970), .ZN(G308));
  OAI211_X1 g793(.A(new_n1216), .B(new_n1217), .C1(new_n977), .C2(new_n974), .ZN(G225));
endmodule


