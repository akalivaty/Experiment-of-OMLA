//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT66), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G20), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n211), .A2(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n222), .B1(new_n203), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n221), .B(new_n226), .C1(G58), .C2(G232), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G1), .B2(G20), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT1), .Z(new_n229));
  AOI211_X1 g0029(.A(new_n217), .B(new_n229), .C1(new_n212), .C2(new_n211), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n220), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n201), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n202), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n219), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  INV_X1    g0049(.A(KEYINPUT90), .ZN(new_n250));
  OR2_X1    g0050(.A1(KEYINPUT88), .A2(G294), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT88), .A2(G294), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G33), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(G257), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n255), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G250), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n253), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n262), .B1(G33), .B2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT5), .A2(G41), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT5), .A2(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n266), .B(G274), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT5), .B(G41), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n263), .B1(new_n271), .B2(new_n266), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n272), .B2(G264), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(KEYINPUT89), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT89), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n264), .A2(new_n273), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n276), .B1(new_n280), .B2(G169), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n262), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n208), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT71), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(new_n208), .A3(G13), .A4(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(G33), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n287), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n290), .A2(new_n292), .ZN(new_n296));
  INV_X1    g0096(.A(G107), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT25), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n293), .B2(G107), .ZN(new_n300));
  AOI22_X1  g0100(.A1(G107), .A2(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT23), .A2(G107), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT65), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT23), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n297), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G116), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n307), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n209), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT22), .ZN(new_n314));
  OR2_X1    g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n304), .A2(new_n306), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(G87), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n316), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n304), .A2(new_n306), .ZN(new_n320));
  AND4_X1   g0120(.A1(new_n314), .A2(new_n319), .A3(new_n320), .A4(G87), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n303), .B(new_n313), .C1(new_n318), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT24), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(G87), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT22), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n319), .A2(new_n320), .A3(new_n314), .A4(G87), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n312), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT24), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n303), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n302), .B1(new_n330), .B2(new_n286), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n250), .B1(new_n281), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n322), .A2(KEYINPUT24), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n327), .B2(new_n303), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n286), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n301), .ZN(new_n336));
  INV_X1    g0136(.A(new_n279), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n278), .B1(new_n264), .B2(new_n273), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n276), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n336), .A2(new_n341), .A3(KEYINPUT90), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(new_n343), .A3(new_n279), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT91), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n274), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n277), .A2(KEYINPUT91), .A3(new_n343), .A4(new_n279), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n332), .A2(new_n342), .B1(new_n331), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G20), .A2(G33), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n205), .A2(G20), .B1(G150), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n320), .A2(G33), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT8), .B(G58), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n286), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n296), .A2(G50), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n296), .A2(new_n286), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n288), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n360), .B2(G50), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(KEYINPUT72), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n363), .B(new_n358), .C1(new_n360), .C2(G50), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n357), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT9), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT69), .B(G1698), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n319), .A2(new_n368), .A3(G222), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  INV_X1    g0170(.A(G1698), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n315), .B2(new_n316), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G223), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n369), .B1(new_n370), .B2(new_n319), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n263), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G41), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(G1), .A3(G13), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G226), .ZN(new_n381));
  INV_X1    g0181(.A(G274), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n376), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G190), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT9), .B(new_n357), .C1(new_n362), .C2(new_n364), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n385), .B2(G200), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n367), .A2(new_n387), .A3(new_n388), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT10), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n388), .A2(new_n390), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT10), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n387), .A4(new_n367), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n385), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n365), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n275), .B2(new_n386), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  OAI211_X1 g0204(.A(G232), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n259), .C2(new_n235), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n383), .B1(new_n406), .B2(new_n263), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n380), .A2(G238), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n403), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n403), .A3(new_n408), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(G190), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n296), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n287), .A2(new_n293), .A3(G68), .A4(new_n288), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT12), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n293), .B2(G68), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT76), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n352), .A2(G50), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n209), .B2(G68), .C1(new_n354), .C2(new_n370), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n286), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT11), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n425), .A3(new_n286), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n419), .A2(new_n420), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n407), .A2(new_n403), .A3(new_n408), .ZN(new_n428));
  OAI21_X1  g0228(.A(G200), .B1(new_n428), .B2(new_n409), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n412), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n428), .B2(new_n409), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n410), .A2(G179), .A3(new_n411), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(G169), .C1(new_n428), .C2(new_n409), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n427), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT16), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G58), .A2(G68), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT77), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G58), .A3(G68), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n444), .C1(G58), .C2(G68), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(G20), .B1(G159), .B2(new_n352), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n254), .A2(new_n255), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n320), .A2(new_n448), .A3(KEYINPUT7), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n315), .A2(new_n209), .A3(new_n316), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT7), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n203), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n440), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n320), .A2(new_n448), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(KEYINPUT7), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(G68), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n446), .A3(KEYINPUT16), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n286), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n355), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n287), .A2(new_n293), .A3(new_n288), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n296), .A2(new_n355), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT78), .B1(new_n259), .B2(new_n374), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n372), .A2(G226), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n319), .A2(new_n368), .A3(new_n468), .A4(G223), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G87), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n466), .A2(new_n467), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n383), .B1(new_n471), .B2(new_n263), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n380), .A2(G232), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(G179), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n397), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT18), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n472), .A2(new_n473), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G169), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n474), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT18), .A3(new_n465), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(G200), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n458), .A2(new_n286), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n463), .B1(new_n486), .B2(new_n454), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n472), .A2(G190), .A3(new_n473), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT17), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT17), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n485), .A2(new_n487), .A3(new_n491), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n293), .A2(G77), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT73), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n359), .A2(G77), .A3(new_n288), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n215), .A2(G77), .ZN(new_n498));
  INV_X1    g0298(.A(new_n352), .ZN(new_n499));
  XOR2_X1   g0299(.A(KEYINPUT15), .B(G87), .Z(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI221_X1 g0301(.A(new_n498), .B1(new_n499), .B2(new_n355), .C1(new_n501), .C2(new_n354), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n286), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n496), .A2(KEYINPUT74), .A3(new_n497), .A4(new_n503), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n373), .A2(new_n223), .B1(new_n259), .B2(new_n232), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n319), .A2(new_n297), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n263), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n380), .A2(G244), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n384), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n506), .A2(new_n507), .B1(new_n397), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n512), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n275), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n439), .A2(new_n484), .A3(new_n493), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n514), .A2(G190), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(G200), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n506), .A2(new_n518), .A3(new_n519), .A4(new_n507), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n402), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n372), .A2(G244), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n309), .C1(new_n223), .C2(new_n259), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n263), .A2(new_n266), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n263), .B1(G250), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n266), .A2(G274), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(G190), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n526), .A2(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n317), .A2(G68), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n215), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n354), .A2(new_n224), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n533), .B(new_n538), .C1(new_n539), .C2(KEYINPUT19), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n286), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n296), .A2(new_n501), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n295), .A2(G87), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT84), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n526), .A2(new_n545), .A3(G190), .A4(new_n528), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n530), .A2(new_n532), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n531), .A2(new_n397), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n526), .A2(new_n275), .A3(new_n528), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n541), .A2(new_n542), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n287), .A2(new_n293), .A3(new_n294), .A4(new_n500), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT83), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n449), .A2(new_n452), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT79), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT6), .ZN(new_n558));
  AND2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(new_n534), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n297), .A2(KEYINPUT6), .A3(G97), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n320), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n499), .A2(new_n370), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n557), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n563), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n297), .A2(KEYINPUT6), .A3(G97), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n558), .ZN(new_n568));
  OAI211_X1 g0368(.A(KEYINPUT79), .B(new_n565), .C1(new_n568), .C2(new_n320), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n556), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n286), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n287), .A2(new_n293), .A3(G97), .A4(new_n294), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n296), .A2(new_n224), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  INV_X1    g0377(.A(G244), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n259), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n372), .B2(G250), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n319), .A2(new_n368), .A3(KEYINPUT4), .A4(G244), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n263), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n266), .B1(new_n268), .B2(new_n267), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G257), .A3(new_n378), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(KEYINPUT80), .A3(G257), .A4(new_n378), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n270), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(new_n275), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n397), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n576), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n574), .B1(new_n570), .B2(new_n286), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n585), .A2(new_n343), .A3(new_n591), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n585), .B2(new_n591), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT81), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n554), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n219), .A2(G20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n286), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n224), .A2(G33), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n215), .A2(new_n581), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n605), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT86), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n224), .A2(G33), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n320), .A2(new_n580), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(new_n286), .A3(new_n606), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(new_n605), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n616), .A3(new_n605), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(G264), .B(G1698), .C1(new_n254), .C2(new_n255), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n315), .A2(G303), .A3(new_n316), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n619), .B(new_n620), .C1(new_n259), .C2(new_n225), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n263), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n586), .A2(G270), .A3(new_n378), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n269), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G200), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n296), .A2(new_n627), .A3(new_n219), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT85), .B1(new_n293), .B2(G116), .ZN(new_n629));
  AOI22_X1  g0429(.A1(G116), .A2(new_n295), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n623), .B1(new_n621), .B2(new_n263), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(G190), .A3(new_n269), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n618), .A2(new_n626), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n618), .A2(new_n630), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n397), .B1(new_n631), .B2(new_n269), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT21), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n270), .B(new_n623), .C1(new_n263), .C2(new_n621), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n635), .A2(KEYINPUT21), .B1(new_n638), .B2(G179), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n628), .A2(new_n629), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n287), .A2(new_n293), .A3(G116), .A4(new_n294), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n614), .A2(new_n616), .A3(new_n605), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n616), .B1(new_n614), .B2(new_n605), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n645), .B2(new_n615), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n637), .B1(new_n639), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n631), .A2(G179), .A3(new_n269), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n625), .A2(G169), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n651), .A2(KEYINPUT87), .A3(new_n634), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n633), .B(new_n636), .C1(new_n647), .C2(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n351), .A2(new_n522), .A3(new_n604), .A4(new_n653), .ZN(G372));
  AND2_X1   g0454(.A1(new_n490), .A2(new_n492), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n513), .A2(new_n430), .A3(new_n515), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n437), .A2(new_n438), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n484), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n396), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n401), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT92), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n554), .B2(new_n595), .ZN(new_n665));
  INV_X1    g0465(.A(new_n595), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n547), .A3(new_n553), .A4(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n554), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n350), .A2(new_n331), .ZN(new_n670));
  INV_X1    g0470(.A(new_n600), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n636), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n646), .B2(new_n639), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n281), .A2(new_n331), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n668), .B(new_n553), .C1(new_n672), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n522), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n663), .A2(new_n678), .ZN(G369));
  NOR2_X1   g0479(.A1(new_n215), .A2(new_n289), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n208), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n351), .B1(new_n331), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n675), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n687), .A2(new_n646), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n674), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n633), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n639), .A2(new_n646), .A3(new_n637), .ZN(new_n695));
  AOI21_X1  g0495(.A(KEYINPUT87), .B1(new_n651), .B2(new_n634), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n673), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n693), .B1(new_n697), .B2(new_n692), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n673), .B1(new_n695), .B2(new_n696), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n687), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(KEYINPUT93), .A3(new_n687), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n690), .A2(new_n707), .B1(new_n675), .B2(new_n687), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n210), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G1), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n534), .A2(new_n535), .A3(new_n219), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n214), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n604), .A2(new_n351), .A3(new_n653), .A4(new_n687), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n531), .A2(new_n275), .A3(new_n625), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n531), .A2(new_n721), .A3(new_n275), .A4(new_n625), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n720), .A2(new_n274), .A3(new_n593), .A4(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n526), .A2(new_n528), .A3(new_n631), .ZN(new_n724));
  INV_X1    g0524(.A(new_n593), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n276), .A4(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n276), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n526), .A2(new_n528), .A3(new_n631), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n724), .A2(new_n276), .A3(new_n725), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n728), .B1(new_n734), .B2(new_n729), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n687), .B1(new_n727), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n718), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n734), .A2(new_n729), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n727), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n665), .A2(KEYINPUT96), .A3(new_n667), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n702), .B1(new_n332), .B2(new_n342), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n553), .B(new_n745), .C1(new_n746), .C2(new_n672), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n667), .A2(KEYINPUT96), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT29), .B(new_n687), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n677), .A2(new_n687), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n744), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n716), .B1(new_n754), .B2(G1), .ZN(G364));
  NAND2_X1  g0555(.A1(new_n245), .A2(G45), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n710), .A2(new_n319), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n756), .B(new_n757), .C1(G45), .C2(new_n214), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n319), .A2(new_n210), .A3(G355), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n758), .B(new_n759), .C1(G116), .C2(new_n210), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n262), .B1(G20), .B2(new_n397), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n764), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n320), .A2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(G179), .A3(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT32), .Z(new_n772));
  NOR2_X1   g0572(.A1(new_n275), .A2(new_n347), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n215), .A2(G190), .A3(new_n773), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(G68), .B1(new_n777), .B2(G50), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n347), .A2(G179), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n768), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n275), .A2(G200), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n215), .A2(G190), .A3(new_n781), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n780), .A2(new_n297), .B1(new_n202), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n779), .A2(G20), .A3(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(G87), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n768), .A2(new_n781), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n343), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n320), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n370), .B1(new_n224), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n448), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n772), .A2(new_n778), .A3(new_n786), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n780), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n251), .A2(new_n252), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n448), .B1(new_n795), .B2(new_n789), .C1(new_n787), .C2(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n797), .C1(G329), .C2(new_n770), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n785), .A2(G303), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n774), .A2(new_n800), .B1(new_n801), .B2(new_n782), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT98), .Z(new_n803));
  XOR2_X1   g0603(.A(new_n776), .B(KEYINPUT97), .Z(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G326), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n798), .A2(new_n799), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n792), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n763), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n766), .B1(new_n767), .B2(new_n808), .C1(new_n698), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n713), .B1(G45), .B2(new_n680), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G330), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n698), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT99), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n506), .A2(new_n507), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n686), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(new_n520), .B1(new_n513), .B2(new_n515), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n513), .A2(new_n515), .A3(new_n687), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT100), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n520), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n516), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n821), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n750), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(new_n744), .ZN(new_n830));
  INV_X1    g0630(.A(new_n811), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n787), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G159), .B1(new_n777), .B2(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n782), .C1(new_n836), .C2(new_n774), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n319), .B1(new_n789), .B2(new_n202), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n780), .A2(new_n203), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(G132), .C2(new_n770), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n838), .B(new_n841), .C1(new_n201), .C2(new_n784), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n782), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n448), .B1(new_n784), .B2(new_n297), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n780), .A2(new_n535), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n845), .B(new_n846), .C1(G303), .C2(new_n777), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n770), .A2(G311), .B1(G116), .B2(new_n833), .ZN(new_n848));
  INV_X1    g0648(.A(new_n789), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n775), .A2(G283), .B1(G97), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n764), .A2(new_n761), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n852), .A2(new_n764), .B1(new_n370), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n811), .C1(new_n828), .C2(new_n762), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n832), .A2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n828), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n739), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n458), .A2(new_n286), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT16), .B1(new_n457), .B2(new_n446), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n464), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n475), .B2(new_n476), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT103), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n489), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n684), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n864), .B1(new_n863), .B2(new_n489), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n465), .A2(new_n866), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n477), .A2(new_n489), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n465), .B1(new_n482), .B2(new_n866), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(new_n871), .A4(new_n489), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n870), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n867), .B1(new_n484), .B2(new_n493), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n871), .B1(new_n875), .B2(new_n489), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n877), .B2(new_n874), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n872), .B1(new_n484), .B2(new_n493), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n437), .A2(new_n438), .A3(new_n686), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n438), .A2(new_n686), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n657), .A2(new_n430), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT102), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n439), .B2(new_n890), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n859), .A2(KEYINPUT40), .A3(new_n888), .A4(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n737), .B1(new_n717), .B2(KEYINPUT31), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n895), .B(new_n828), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(KEYINPUT105), .A3(KEYINPUT40), .A4(new_n888), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  INV_X1    g0705(.A(new_n882), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n879), .B2(new_n881), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n908), .B2(new_n901), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n739), .A2(new_n858), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n522), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n910), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(G330), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n882), .A2(new_n887), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT39), .B1(new_n906), .B2(new_n907), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n657), .A2(new_n686), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n821), .B1(new_n750), .B2(new_n857), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n895), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(new_n908), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n659), .A2(new_n684), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n749), .A2(new_n752), .A3(new_n522), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n663), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n927), .B(new_n929), .Z(new_n930));
  XNOR2_X1  g0730(.A(new_n915), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n208), .B2(new_n680), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT35), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n216), .B1(new_n568), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(G116), .C1(new_n933), .C2(new_n568), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n203), .A2(G50), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT101), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n442), .A2(new_n444), .A3(G77), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n214), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(G1), .A3(new_n289), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n932), .A2(new_n936), .A3(new_n941), .ZN(G367));
  NAND2_X1  g0742(.A1(new_n849), .A2(G68), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n836), .B2(new_n782), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT111), .Z(new_n945));
  INV_X1    g0745(.A(G159), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n774), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n780), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(G77), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n201), .B2(new_n787), .ZN(new_n950));
  INV_X1    g0750(.A(new_n770), .ZN(new_n951));
  INV_X1    g0751(.A(G137), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n319), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n945), .A2(new_n947), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n202), .B2(new_n784), .C1(new_n835), .C2(new_n804), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G97), .A2(new_n948), .B1(new_n833), .B2(G283), .ZN(new_n956));
  INV_X1    g0756(.A(G317), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n957), .B2(new_n951), .ZN(new_n958));
  INV_X1    g0758(.A(new_n782), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(G303), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n784), .A2(new_n219), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n805), .A2(G311), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n448), .B1(new_n789), .B2(new_n297), .C1(new_n961), .C2(KEYINPUT46), .ZN(new_n964));
  INV_X1    g0764(.A(new_n795), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n964), .B1(new_n965), .B2(new_n775), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n960), .A2(new_n962), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n955), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n764), .ZN(new_n970));
  INV_X1    g0770(.A(new_n757), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n765), .B1(new_n210), .B2(new_n501), .C1(new_n239), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n687), .A2(new_n544), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n669), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n553), .B2(new_n973), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(new_n809), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n811), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n671), .B1(new_n596), .B2(new_n687), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n666), .A2(new_n686), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n707), .A2(new_n690), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT42), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n332), .A2(new_n342), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n595), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n687), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n707), .A2(new_n690), .A3(new_n987), .A4(new_n981), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT106), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT106), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n983), .A2(new_n991), .A3(new_n986), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n993), .A2(new_n994), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n993), .A2(KEYINPUT107), .A3(new_n994), .A4(new_n995), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n981), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n701), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n998), .A2(new_n1003), .A3(new_n999), .A4(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n208), .B1(new_n680), .B2(G45), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n708), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT108), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1002), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n708), .C2(new_n981), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT45), .B1(new_n708), .B2(new_n981), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1013), .B(new_n1016), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n700), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n1017), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1023), .A2(new_n701), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n691), .A2(new_n699), .A3(new_n705), .A4(new_n706), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT109), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n707), .B2(new_n690), .ZN(new_n1027));
  OAI211_X1 g0827(.A(G330), .B(new_n698), .C1(new_n690), .C2(new_n707), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n744), .B(new_n753), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1021), .A2(new_n1024), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n754), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n711), .B(KEYINPUT41), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1009), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT110), .B1(new_n1007), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n1008), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT110), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n978), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(G387));
  INV_X1    g0843(.A(G303), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n787), .A2(new_n1044), .B1(new_n957), .B2(new_n782), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT112), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n796), .B2(new_n774), .C1(new_n801), .C2(new_n804), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n793), .B2(new_n789), .C1(new_n795), .C2(new_n784), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n948), .A2(G116), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n319), .B1(new_n770), .B2(G326), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n951), .A2(new_n836), .B1(new_n201), .B2(new_n782), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n787), .A2(new_n203), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n224), .A2(new_n780), .B1(new_n774), .B2(new_n355), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n849), .A2(new_n500), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n784), .A2(new_n370), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1058), .A2(new_n448), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n946), .C2(new_n776), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n764), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n691), .A2(new_n763), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n460), .A2(new_n201), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n714), .B1(new_n1064), .B2(KEYINPUT50), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1065), .B(new_n265), .C1(KEYINPUT50), .C2(new_n1064), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G68), .B2(G77), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n757), .B1(new_n236), .B2(new_n265), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n319), .A2(new_n210), .A3(new_n714), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n210), .A2(G107), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n765), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1062), .A2(new_n1063), .A3(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1073), .A2(new_n811), .B1(new_n1009), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n711), .B1(new_n1074), .B2(new_n754), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1075), .B1(new_n1032), .B2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n1008), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n789), .A2(new_n370), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n951), .A2(new_n835), .B1(new_n355), .B2(new_n787), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G50), .C2(new_n775), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n836), .A2(new_n776), .B1(new_n782), .B2(new_n946), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n448), .B(new_n846), .C1(G68), .C2(new_n785), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT113), .Z(new_n1087));
  NOR2_X1   g0887(.A1(new_n774), .A2(new_n1044), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n948), .A2(G107), .B1(G116), .B2(new_n849), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n319), .B1(new_n785), .B2(G283), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(new_n843), .C2(new_n787), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT52), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n796), .A2(new_n782), .B1(new_n776), .B2(new_n957), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1088), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n1092), .B2(new_n1093), .C1(new_n801), .C2(new_n951), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n831), .B1(new_n1096), .B2(new_n764), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n765), .B1(new_n224), .B2(new_n210), .C1(new_n248), .C2(new_n971), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n809), .C2(new_n981), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1078), .A2(new_n1031), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n711), .A3(new_n1033), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT114), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT114), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1104), .A3(new_n711), .A4(new_n1033), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1079), .B(new_n1100), .C1(new_n1103), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  AND2_X1   g0907(.A1(new_n918), .A2(new_n919), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n921), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n924), .A2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n687), .B(new_n828), .C1(new_n747), .C2(new_n748), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n821), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n895), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n916), .A2(new_n921), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1108), .A2(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n743), .A2(G330), .A3(new_n828), .A4(new_n895), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n859), .A2(KEYINPUT116), .A3(G330), .A4(new_n895), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT116), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n901), .B2(new_n813), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1116), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1115), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n1115), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n742), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n828), .C1(new_n899), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n895), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1117), .A2(new_n1119), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n923), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1112), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n828), .C1(new_n899), .C2(new_n900), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1129), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1116), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n663), .B(new_n928), .C1(new_n813), .C2(new_n912), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1126), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(KEYINPUT117), .B(new_n1138), .C1(new_n1132), .C2(new_n1136), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1125), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1116), .A2(new_n1135), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n923), .A2(new_n1131), .B1(new_n1143), .B2(new_n1133), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT117), .B1(new_n1144), .B2(new_n1138), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1137), .A2(new_n1126), .A3(new_n1139), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1115), .A2(new_n1124), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .A4(new_n1123), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1148), .A3(new_n711), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1125), .A2(new_n1009), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n951), .A2(new_n843), .B1(new_n219), .B2(new_n782), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n840), .B(new_n1151), .C1(G97), .C2(new_n833), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n448), .B1(new_n370), .B2(new_n789), .C1(new_n774), .C2(new_n297), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G283), .B2(new_n777), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n535), .C2(new_n784), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n319), .B1(new_n776), .B2(new_n1156), .C1(new_n946), .C2(new_n789), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(G137), .B2(new_n775), .ZN(new_n1158));
  INV_X1    g0958(.A(G132), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n780), .A2(new_n201), .B1(new_n1159), .B2(new_n782), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT54), .B(G143), .Z(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n833), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n770), .A2(G125), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n784), .A2(new_n836), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT53), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1158), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n767), .B1(new_n1155), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n355), .B2(new_n853), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n811), .B(new_n1168), .C1(new_n920), .C2(new_n762), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1149), .A2(new_n1150), .A3(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n396), .A2(new_n1171), .A3(new_n401), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n396), .B2(new_n401), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n365), .B(new_n866), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1174), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n365), .A2(new_n866), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(new_n1172), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1180), .A3(new_n1178), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n761), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n853), .A2(new_n201), .ZN(new_n1186));
  INV_X1    g0986(.A(G125), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n774), .A2(new_n1159), .B1(new_n1187), .B2(new_n776), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G150), .A2(new_n849), .B1(new_n959), .B2(G128), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n952), .B2(new_n787), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(new_n785), .C2(new_n1161), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT59), .ZN(new_n1192));
  AOI21_X1  g0992(.A(G41), .B1(new_n770), .B2(G124), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G33), .B1(new_n948), .B2(G159), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n201), .B1(new_n254), .B2(G41), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n319), .B(new_n1058), .C1(new_n959), .C2(G107), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n224), .B2(new_n774), .C1(new_n219), .C2(new_n776), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n770), .A2(G283), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n833), .A2(new_n500), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n948), .A2(G58), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n943), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n1198), .A2(G41), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT58), .Z(new_n1204));
  NAND3_X1  g1004(.A1(new_n1195), .A2(new_n1196), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n831), .B1(new_n1205), .B2(new_n764), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1185), .A2(new_n1186), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT119), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n898), .A2(new_n903), .A3(G330), .A4(new_n909), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1208), .B(new_n927), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n904), .A2(new_n1184), .A3(G330), .A4(new_n909), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n927), .A2(new_n1208), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1207), .B1(new_n1218), .B2(new_n1008), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1214), .A2(new_n1216), .A3(new_n927), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n927), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1138), .B1(new_n1225), .B2(new_n1125), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n711), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1142), .A2(new_n1139), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1215), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1220), .B1(new_n1227), .B2(new_n1232), .ZN(G375));
  AOI22_X1  g1033(.A1(new_n770), .A2(G303), .B1(new_n959), .B2(G283), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n1057), .C1(new_n297), .C2(new_n787), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n775), .A2(G116), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n777), .A2(G294), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n319), .B1(new_n785), .B2(G97), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n949), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1235), .A2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT120), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1201), .B1(new_n201), .B2(new_n789), .C1(new_n1159), .C2(new_n776), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n951), .A2(new_n1156), .B1(new_n952), .B2(new_n782), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1161), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n319), .B1(new_n946), .B2(new_n784), .C1(new_n774), .C2(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n836), .B2(new_n787), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1241), .A2(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT121), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n831), .B1(new_n1249), .B2(new_n764), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n853), .A2(new_n203), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n762), .C2(new_n895), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1144), .B2(new_n1008), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1132), .A2(new_n1138), .A3(new_n1136), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1145), .A2(new_n1146), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1253), .B1(new_n1256), .B2(new_n1035), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G381));
  INV_X1    g1058(.A(KEYINPUT57), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n927), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1259), .B1(new_n1261), .B2(new_n1221), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n712), .B1(new_n1228), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1259), .B1(new_n1226), .B2(new_n1218), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1219), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1150), .A2(new_n1169), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n712), .B1(new_n1225), .B2(new_n1125), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1148), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1075), .B(new_n816), .C1(new_n1032), .C2(new_n1076), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1270), .A2(G384), .ZN(new_n1271));
  AND4_X1   g1071(.A1(new_n1042), .A2(new_n1106), .A3(new_n1257), .A4(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1269), .B1(new_n1272), .B2(KEYINPUT122), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1042), .A2(new_n1106), .A3(new_n1257), .A4(new_n1271), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT122), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1274), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1278), .A2(new_n1279), .ZN(G407));
  NAND3_X1  g1080(.A1(new_n1265), .A2(new_n685), .A3(new_n1268), .ZN(new_n1281));
  OAI211_X1 g1081(.A(G213), .B(new_n1281), .C1(new_n1278), .C2(new_n1279), .ZN(G409));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1228), .A2(new_n1035), .A3(new_n1231), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1008), .B1(new_n1261), .B2(new_n1221), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1268), .A2(new_n1287), .A3(new_n1207), .A4(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1286), .B(new_n1290), .C1(new_n1265), .C2(new_n1268), .ZN(new_n1291));
  INV_X1    g1091(.A(G384), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1254), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n711), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1255), .B2(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1296), .B2(new_n1253), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT124), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1296), .A2(new_n1292), .A3(new_n1253), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT124), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1300), .B(new_n1292), .C1(new_n1296), .C2(new_n1253), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(KEYINPUT62), .B1(new_n1291), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1285), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1298), .A2(new_n1299), .A3(new_n1304), .A4(new_n1301), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1291), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1302), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G375), .A2(G378), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1207), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(G378), .A2(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1226), .A2(new_n1218), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1288), .B1(new_n1313), .B2(new_n1035), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1285), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1309), .A2(new_n1310), .A3(new_n1315), .A4(new_n1316), .ZN(new_n1317));
  AND4_X1   g1117(.A1(new_n1283), .A2(new_n1303), .A3(new_n1308), .A4(new_n1317), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1042), .A2(new_n1106), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1042), .A2(new_n1106), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G393), .A2(G396), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1270), .ZN(new_n1322));
  OAI22_X1  g1122(.A1(new_n1319), .A2(new_n1320), .B1(KEYINPUT125), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(G390), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1042), .A2(new_n1106), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1322), .B(KEYINPUT125), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1323), .A2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1291), .A2(new_n1302), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1329), .B1(new_n1308), .B2(KEYINPUT63), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1309), .A2(new_n1310), .A3(new_n1315), .A4(KEYINPUT63), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1283), .A3(new_n1331), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1318), .A2(new_n1328), .B1(new_n1330), .B2(new_n1332), .ZN(G405));
  AND2_X1   g1133(.A1(new_n1310), .A2(new_n1269), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1309), .A2(KEYINPUT126), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1328), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1328), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1341), .A3(new_n1336), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1342), .ZN(G402));
endmodule


