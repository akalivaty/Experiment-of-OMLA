

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  NOR2_X1 U324 ( .A1(n587), .A2(n453), .ZN(n455) );
  NOR2_X1 U325 ( .A1(n423), .A2(n422), .ZN(n424) );
  XOR2_X1 U326 ( .A(KEYINPUT38), .B(n456), .Z(n504) );
  XOR2_X1 U327 ( .A(n373), .B(KEYINPUT21), .Z(n292) );
  XOR2_X1 U328 ( .A(KEYINPUT101), .B(n417), .Z(n293) );
  AND2_X1 U329 ( .A1(n548), .A2(n550), .ZN(n461) );
  XNOR2_X1 U330 ( .A(G211GAT), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U331 ( .A(n375), .B(n320), .ZN(n321) );
  XNOR2_X1 U332 ( .A(n439), .B(n321), .ZN(n322) );
  XNOR2_X1 U333 ( .A(n326), .B(n325), .ZN(n327) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n406) );
  NAND2_X1 U335 ( .A1(n432), .A2(n431), .ZN(n487) );
  XNOR2_X1 U336 ( .A(n328), .B(n327), .ZN(n330) );
  XNOR2_X1 U337 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U338 ( .A(n409), .B(n408), .ZN(n416) );
  XOR2_X1 U339 ( .A(KEYINPUT41), .B(n579), .Z(n550) );
  INV_X1 U340 ( .A(G29GAT), .ZN(n457) );
  XNOR2_X1 U341 ( .A(n481), .B(n406), .ZN(n482) );
  XNOR2_X1 U342 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U343 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n396) );
  XOR2_X1 U348 ( .A(G162GAT), .B(n396), .Z(n297) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U351 ( .A(G29GAT), .B(n298), .ZN(n315) );
  XOR2_X1 U352 ( .A(KEYINPUT98), .B(KEYINPUT6), .Z(n300) );
  XNOR2_X1 U353 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U355 ( .A(G57GAT), .B(G120GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(G1GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U359 ( .A(G85GAT), .B(G148GAT), .Z(n306) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(G155GAT), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(n309), .B(KEYINPUT1), .Z(n313) );
  XOR2_X1 U364 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n311) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT95), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n382) );
  XNOR2_X1 U367 ( .A(n382), .B(KEYINPUT97), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n315), .B(n314), .Z(n570) );
  INV_X1 U370 ( .A(n570), .ZN(n509) );
  XOR2_X1 U371 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n317) );
  XNOR2_X1 U372 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n332) );
  XOR2_X1 U374 ( .A(G57GAT), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U375 ( .A(KEYINPUT13), .B(KEYINPUT74), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n439) );
  XOR2_X1 U377 ( .A(G148GAT), .B(G78GAT), .Z(n375) );
  AND2_X1 U378 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n322), .B(KEYINPUT76), .ZN(n328) );
  XOR2_X1 U380 ( .A(G85GAT), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n361) );
  XOR2_X1 U383 ( .A(n361), .B(KEYINPUT31), .Z(n326) );
  INV_X1 U384 ( .A(G204GAT), .ZN(n325) );
  XOR2_X1 U385 ( .A(G120GAT), .B(G71GAT), .Z(n393) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(n393), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n579) );
  XOR2_X1 U389 ( .A(G141GAT), .B(G22GAT), .Z(n334) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G197GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n336) );
  XOR2_X1 U392 ( .A(G50GAT), .B(G36GAT), .Z(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n352) );
  XOR2_X1 U394 ( .A(G1GAT), .B(G15GAT), .Z(n338) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G113GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U397 ( .A(G8GAT), .B(KEYINPUT69), .Z(n340) );
  XNOR2_X1 U398 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n350) );
  XOR2_X1 U401 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n344) );
  XNOR2_X1 U402 ( .A(KEYINPUT8), .B(G29GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(KEYINPUT7), .B(n345), .Z(n371) );
  XOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n371), .B(n348), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n354) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U412 ( .A(n354), .B(n353), .Z(n548) );
  INV_X1 U413 ( .A(n548), .ZN(n575) );
  NOR2_X1 U414 ( .A1(n579), .A2(n575), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n355), .B(KEYINPUT78), .ZN(n488) );
  XOR2_X1 U416 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n357) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT11), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U419 ( .A(n358), .B(KEYINPUT10), .Z(n360) );
  XOR2_X1 U420 ( .A(G50GAT), .B(G162GAT), .Z(n378) );
  XNOR2_X1 U421 ( .A(n378), .B(KEYINPUT80), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n365) );
  XOR2_X1 U423 ( .A(n361), .B(KEYINPUT79), .Z(n363) );
  NAND2_X1 U424 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U426 ( .A(n365), .B(n364), .Z(n369) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G190GAT), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n366), .B(G134GAT), .ZN(n403) );
  XNOR2_X1 U429 ( .A(G36GAT), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n367), .B(KEYINPUT81), .ZN(n410) );
  XNOR2_X1 U431 ( .A(n403), .B(n410), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n557) );
  XNOR2_X1 U434 ( .A(KEYINPUT82), .B(n557), .ZN(n543) );
  XOR2_X1 U435 ( .A(KEYINPUT36), .B(n543), .Z(n587) );
  XNOR2_X1 U436 ( .A(n372), .B(KEYINPUT93), .ZN(n373) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n292), .B(n374), .ZN(n409) );
  XOR2_X1 U439 ( .A(G106GAT), .B(G218GAT), .Z(n377) );
  XOR2_X1 U440 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XNOR2_X1 U441 ( .A(n436), .B(n375), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U443 ( .A(n379), .B(n378), .Z(n388) );
  XOR2_X1 U444 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n381) );
  XNOR2_X1 U445 ( .A(KEYINPUT22), .B(KEYINPUT96), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U447 ( .A(n382), .B(KEYINPUT24), .Z(n384) );
  NAND2_X1 U448 ( .A1(G228GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U450 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n409), .B(n389), .ZN(n475) );
  XOR2_X1 U453 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n391) );
  NAND2_X1 U454 ( .A1(G227GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U456 ( .A(n392), .B(G99GAT), .Z(n395) );
  XOR2_X1 U457 ( .A(G15GAT), .B(G127GAT), .Z(n447) );
  XNOR2_X1 U458 ( .A(n447), .B(n393), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U460 ( .A(n397), .B(n396), .Z(n405) );
  XOR2_X1 U461 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n399) );
  XNOR2_X1 U462 ( .A(KEYINPUT90), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U464 ( .A(n400), .B(G183GAT), .Z(n402) );
  XNOR2_X1 U465 ( .A(G169GAT), .B(G176GAT), .ZN(n401) );
  XNOR2_X1 U466 ( .A(n402), .B(n401), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n414), .B(n403), .ZN(n404) );
  XOR2_X1 U468 ( .A(n405), .B(n404), .Z(n514) );
  XOR2_X1 U469 ( .A(G8GAT), .B(KEYINPUT83), .Z(n435) );
  XOR2_X1 U470 ( .A(n435), .B(G92GAT), .Z(n407) );
  XOR2_X1 U471 ( .A(n410), .B(G64GAT), .Z(n412) );
  NAND2_X1 U472 ( .A1(G226GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(n414), .B(n413), .Z(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n524) );
  INV_X1 U476 ( .A(n524), .ZN(n512) );
  NAND2_X1 U477 ( .A1(n514), .A2(n512), .ZN(n417) );
  NAND2_X1 U478 ( .A1(n475), .A2(n293), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n418), .B(KEYINPUT102), .ZN(n419) );
  XNOR2_X1 U480 ( .A(KEYINPUT25), .B(n419), .ZN(n423) );
  NOR2_X1 U481 ( .A1(n514), .A2(n475), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT26), .B(n420), .Z(n572) );
  XOR2_X1 U483 ( .A(KEYINPUT27), .B(n512), .Z(n426) );
  NOR2_X1 U484 ( .A1(n572), .A2(n426), .ZN(n421) );
  XNOR2_X1 U485 ( .A(KEYINPUT100), .B(n421), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n424), .B(KEYINPUT103), .ZN(n425) );
  NAND2_X1 U487 ( .A1(n425), .A2(n570), .ZN(n432) );
  NOR2_X1 U488 ( .A1(n570), .A2(n426), .ZN(n531) );
  INV_X1 U489 ( .A(n531), .ZN(n429) );
  XOR2_X1 U490 ( .A(KEYINPUT28), .B(n475), .Z(n517) );
  INV_X1 U491 ( .A(n517), .ZN(n534) );
  XNOR2_X1 U492 ( .A(n514), .B(KEYINPUT91), .ZN(n427) );
  NAND2_X1 U493 ( .A1(n534), .A2(n427), .ZN(n428) );
  NOR2_X1 U494 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n430), .B(KEYINPUT99), .ZN(n431) );
  XOR2_X1 U496 ( .A(KEYINPUT85), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G1GAT), .B(G183GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n451) );
  XOR2_X1 U499 ( .A(n435), .B(G78GAT), .Z(n438) );
  XNOR2_X1 U500 ( .A(G211GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n443) );
  XOR2_X1 U502 ( .A(KEYINPUT86), .B(n439), .Z(n441) );
  NAND2_X1 U503 ( .A1(G231GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U505 ( .A(n443), .B(n442), .Z(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT84), .B(KEYINPUT14), .Z(n445) );
  XNOR2_X1 U507 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n451), .B(n450), .ZN(n582) );
  INV_X1 U512 ( .A(n582), .ZN(n568) );
  NAND2_X1 U513 ( .A1(n487), .A2(n568), .ZN(n452) );
  XNOR2_X1 U514 ( .A(KEYINPUT108), .B(n452), .ZN(n453) );
  XNOR2_X1 U515 ( .A(KEYINPUT37), .B(KEYINPUT109), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n522) );
  NAND2_X1 U517 ( .A1(n488), .A2(n522), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n509), .A2(n504), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n458) );
  INV_X1 U520 ( .A(n543), .ZN(n484) );
  XOR2_X1 U521 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n478) );
  XNOR2_X1 U522 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n472) );
  XNOR2_X1 U523 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n582), .A2(n557), .ZN(n463) );
  AND2_X1 U526 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT47), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n587), .A2(n568), .ZN(n466) );
  XNOR2_X1 U529 ( .A(KEYINPUT45), .B(n466), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n575), .ZN(n468) );
  OR2_X1 U531 ( .A1(n579), .A2(n468), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(n530) );
  NAND2_X1 U534 ( .A1(n512), .A2(n530), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(n571) );
  AND2_X1 U537 ( .A1(n475), .A2(n570), .ZN(n476) );
  NAND2_X1 U538 ( .A1(n571), .A2(n476), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  INV_X1 U540 ( .A(n514), .ZN(n532) );
  NOR2_X1 U541 ( .A1(n479), .A2(n532), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(KEYINPUT123), .ZN(n560) );
  NOR2_X1 U543 ( .A1(n484), .A2(n560), .ZN(n483) );
  XNOR2_X1 U544 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n481) );
  NAND2_X1 U545 ( .A1(n484), .A2(n582), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n485), .Z(n486) );
  AND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n507) );
  NAND2_X1 U548 ( .A1(n507), .A2(n488), .ZN(n496) );
  NOR2_X1 U549 ( .A1(n570), .A2(n496), .ZN(n489) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n489), .Z(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT34), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n524), .A2(n496), .ZN(n491) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(n491), .Z(n492) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n492), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n532), .A2(n496), .ZN(n494) );
  XNOR2_X1 U556 ( .A(KEYINPUT105), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n495), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n534), .A2(n496), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(n497), .Z(n498) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n512), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT110), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n502) );
  NAND2_X1 U566 ( .A1(n504), .A2(n514), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT112), .ZN(n506) );
  NAND2_X1 U570 ( .A1(n517), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  INV_X1 U573 ( .A(n550), .ZN(n562) );
  NOR2_X1 U574 ( .A1(n562), .A2(n548), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n521), .A2(n507), .ZN(n508) );
  XNOR2_X1 U576 ( .A(KEYINPUT113), .B(n508), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n509), .A2(n518), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U579 ( .A1(n512), .A2(n518), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n513), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n518), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT114), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n527) );
  NOR2_X1 U588 ( .A1(n570), .A2(n527), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n532), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n534), .A2(n527), .ZN(n528) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n532), .A2(n547), .ZN(n533) );
  XNOR2_X1 U599 ( .A(KEYINPUT116), .B(n533), .ZN(n535) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(KEYINPUT117), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n544), .A2(n548), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT118), .B(n537), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n544), .A2(n550), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n582), .A2(n544), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n572), .A2(n547), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n552) );
  NAND2_X1 U618 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .Z(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n582), .A2(n556), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n575), .ZN(n561) );
  XOR2_X1 U628 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n560), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n560), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  AND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n574) );
  INV_X1 U638 ( .A(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n575), .A2(n586), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  INV_X1 U645 ( .A(n586), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n583), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1354GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(n588), .Z(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

