//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .A3(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n190), .A3(new_n198), .A4(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G137), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n207), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G137), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(new_n207), .A3(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n197), .A2(new_n190), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n193), .A2(new_n218), .B1(new_n219), .B2(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT2), .A2(G113), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n225), .A2(new_n226), .B1(KEYINPUT2), .B2(G113), .ZN(new_n227));
  XNOR2_X1  g041(.A(G116), .B(G119), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT28), .B1(new_n222), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n200), .A2(new_n234), .A3(new_n208), .A4(new_n211), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n233), .A2(new_n231), .A3(new_n221), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n238), .A2(new_n239), .B1(new_n231), .B2(new_n222), .ZN(new_n240));
  XOR2_X1   g054(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n241));
  AOI21_X1  g055(.A(new_n232), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G210), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n243), .A2(G237), .A3(G953), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G101), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT29), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n212), .A2(new_n251), .A3(new_n221), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n233), .A2(new_n221), .A3(new_n235), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(KEYINPUT30), .ZN(new_n254));
  OAI22_X1  g068(.A1(new_n238), .A2(new_n239), .B1(new_n254), .B2(new_n231), .ZN(new_n255));
  INV_X1    g069(.A(new_n249), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G902), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n236), .B(new_n237), .ZN(new_n260));
  INV_X1    g074(.A(new_n231), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n253), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n253), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n232), .B1(new_n266), .B2(KEYINPUT28), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT29), .A3(new_n249), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n259), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G472), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT31), .B1(new_n255), .B2(new_n256), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n254), .A2(new_n231), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n260), .A4(new_n249), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n271), .B(new_n274), .C1(new_n242), .C2(new_n249), .ZN(new_n275));
  INV_X1    g089(.A(G472), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n259), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(KEYINPUT32), .A3(new_n276), .A4(new_n259), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G140), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G125), .ZN(new_n283));
  INV_X1    g097(.A(G125), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G140), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT16), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT72), .B1(new_n283), .B2(KEYINPUT16), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G146), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n283), .A2(new_n285), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n191), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n294));
  INV_X1    g108(.A(G128), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(G119), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(G119), .B2(new_n295), .ZN(new_n297));
  OAI22_X1  g111(.A1(new_n296), .A2(new_n297), .B1(G119), .B2(new_n295), .ZN(new_n298));
  XNOR2_X1  g112(.A(G119), .B(G128), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT24), .B(G110), .Z(new_n300));
  OAI22_X1  g114(.A1(new_n298), .A2(G110), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n291), .A2(new_n293), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n290), .B(new_n191), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n298), .A2(G110), .B1(new_n299), .B2(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT22), .B(G137), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT73), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n311), .B(KEYINPUT74), .Z(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G234), .ZN(new_n315));
  AOI21_X1  g129(.A(G902), .B1(new_n315), .B2(G217), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n316), .B(KEYINPUT76), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(G902), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n319), .A2(KEYINPUT75), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G217), .B1(new_n315), .B2(G902), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT75), .B(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n318), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n281), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G469), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n330));
  INV_X1    g144(.A(G107), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G104), .ZN(new_n332));
  INV_X1    g146(.A(G104), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G107), .ZN(new_n334));
  OAI21_X1  g148(.A(G101), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(KEYINPUT80), .B(G101), .C1(new_n332), .C2(new_n334), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n195), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n199), .B1(new_n340), .B2(new_n219), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT3), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n331), .A4(G104), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n333), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n333), .A2(G107), .B1(KEYINPUT78), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n348), .A2(KEYINPUT79), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(KEYINPUT79), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n339), .B(new_n341), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT4), .B(new_n357), .C1(new_n349), .C2(new_n350), .ZN(new_n358));
  OR2_X1    g172(.A1(new_n357), .A2(KEYINPUT4), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n220), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n344), .A2(new_n346), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n347), .A4(new_n345), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(KEYINPUT79), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n363), .A2(new_n364), .B1(new_n337), .B2(new_n338), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT10), .A3(new_n200), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n351), .A2(KEYINPUT81), .A3(new_n352), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n355), .A2(new_n360), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n215), .B(KEYINPUT82), .Z(new_n369));
  OAI21_X1  g183(.A(new_n351), .B1(new_n365), .B2(new_n200), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n370), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT12), .B1(new_n370), .B2(new_n215), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n368), .A2(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n309), .A2(G227), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n282), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT77), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(G110), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n330), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n371), .A2(new_n372), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n360), .A2(new_n366), .ZN(new_n381));
  INV_X1    g195(.A(new_n369), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(new_n355), .A3(new_n367), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n380), .A2(KEYINPUT84), .A3(new_n377), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n368), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n381), .A2(KEYINPUT83), .A3(new_n355), .A4(new_n367), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n215), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n377), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n329), .B(new_n259), .C1(new_n385), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n380), .A2(new_n378), .A3(new_n383), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n368), .A2(new_n369), .ZN(new_n393));
  INV_X1    g207(.A(new_n215), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n368), .B2(new_n386), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n395), .B2(new_n388), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n392), .B1(new_n396), .B2(new_n378), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G469), .ZN(new_n398));
  NAND2_X1  g212(.A1(G469), .A2(G902), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n391), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  MUX2_X1   g216(.A(new_n220), .B(new_n200), .S(new_n284), .Z(new_n403));
  NAND2_X1  g217(.A1(new_n309), .A2(G224), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT7), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n403), .B(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n261), .A2(new_n358), .A3(new_n359), .ZN(new_n407));
  INV_X1    g221(.A(G116), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n408), .A2(KEYINPUT5), .A3(G119), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n228), .B2(KEYINPUT5), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n229), .B1(G113), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n365), .ZN(new_n412));
  XOR2_X1   g226(.A(G110), .B(G122), .Z(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n411), .B(new_n365), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n413), .B(KEYINPUT8), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n406), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(new_n259), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n407), .A2(new_n412), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n403), .B(new_n404), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n424), .A3(new_n413), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G210), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n426), .A3(new_n428), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n402), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(KEYINPUT9), .B(G234), .Z(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n400), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G237), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n309), .A3(G214), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(new_n188), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(KEYINPUT18), .A3(G131), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n292), .B(new_n191), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n206), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n440), .B(new_n441), .C1(new_n439), .C2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT85), .ZN(new_n445));
  OR3_X1    g259(.A1(new_n439), .A2(KEYINPUT86), .A3(G131), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(G131), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(new_n439), .B2(G131), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n292), .B(KEYINPUT19), .Z(new_n450));
  OAI211_X1 g264(.A(new_n449), .B(new_n291), .C1(G146), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G113), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n333), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n439), .A2(KEYINPUT17), .A3(G131), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n303), .B(new_n457), .C1(KEYINPUT17), .C2(new_n449), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n445), .A3(new_n454), .ZN(new_n459));
  AOI21_X1  g273(.A(G475), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n259), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n463), .A3(new_n259), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n459), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n454), .B1(new_n458), .B2(new_n445), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n259), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G475), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G952), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n315), .B2(new_n437), .ZN(new_n474));
  AOI211_X1 g288(.A(new_n259), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n188), .A2(G128), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n188), .A2(G128), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT88), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n480), .A2(new_n202), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n483), .B(KEYINPUT90), .Z(new_n484));
  INV_X1    g298(.A(G122), .ZN(new_n485));
  OR3_X1    g299(.A1(new_n485), .A2(KEYINPUT87), .A3(G116), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT87), .B1(new_n485), .B2(G116), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n486), .A2(new_n487), .B1(G116), .B2(new_n485), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(new_n331), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n480), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n482), .A2(new_n490), .ZN(new_n493));
  OAI21_X1  g307(.A(G134), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n484), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n202), .B1(new_n480), .B2(new_n482), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n483), .A2(new_n496), .A3(KEYINPUT91), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n485), .A2(G116), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n331), .B1(new_n498), .B2(KEYINPUT14), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n488), .B(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT91), .B1(new_n483), .B2(new_n496), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n497), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n433), .A2(G217), .A3(new_n309), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n495), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n259), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n510), .A2(KEYINPUT92), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(KEYINPUT92), .ZN(new_n512));
  OAI21_X1  g326(.A(G478), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n509), .B(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n471), .A2(new_n478), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n328), .A2(new_n436), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(G101), .ZN(G3));
  AND2_X1   g331(.A1(new_n400), .A2(new_n435), .ZN(new_n518));
  INV_X1    g332(.A(new_n277), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n276), .B1(new_n275), .B2(new_n259), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n326), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n508), .A2(KEYINPUT33), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT33), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n505), .A2(new_n524), .A3(new_n507), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(G478), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n508), .A2(new_n527), .A3(new_n259), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n259), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n470), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n432), .A2(new_n478), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n522), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT34), .B(G104), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT93), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n534), .B(new_n536), .ZN(G6));
  XOR2_X1   g351(.A(new_n509), .B(new_n513), .Z(new_n538));
  INV_X1    g352(.A(new_n464), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n539), .A2(new_n462), .A3(KEYINPUT94), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(KEYINPUT94), .B2(new_n462), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n538), .B(new_n469), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n522), .A2(new_n533), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G107), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(G9));
  NAND2_X1  g359(.A1(new_n323), .A2(new_n325), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n313), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n306), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n546), .B1(new_n317), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n515), .A2(new_n436), .A3(new_n521), .A4(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT37), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G110), .ZN(G12));
  OAI21_X1  g368(.A(new_n474), .B1(new_n476), .B2(G900), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n542), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(new_n436), .A3(new_n281), .A4(new_n551), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G128), .ZN(G30));
  XNOR2_X1  g373(.A(new_n555), .B(KEYINPUT39), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n518), .A2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT40), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT40), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n551), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n430), .A2(new_n431), .ZN(new_n565));
  XOR2_X1   g379(.A(new_n565), .B(KEYINPUT95), .Z(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT38), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n259), .B1(new_n266), .B2(new_n249), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n256), .B1(new_n272), .B2(new_n260), .ZN(new_n569));
  OAI21_X1  g383(.A(G472), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n279), .A2(new_n280), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n538), .A2(new_n470), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n572), .A2(new_n402), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n564), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT97), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n188), .ZN(G45));
  NAND3_X1  g391(.A1(new_n531), .A2(new_n470), .A3(new_n555), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n281), .A2(new_n579), .A3(new_n436), .A4(new_n551), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G146), .ZN(G48));
  NOR2_X1   g395(.A1(new_n532), .A2(new_n533), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n379), .B(new_n384), .C1(new_n396), .C2(new_n377), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n259), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(G469), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n583), .B(new_n259), .C1(KEYINPUT98), .C2(new_n329), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n586), .A2(new_n435), .A3(new_n587), .ZN(new_n588));
  AND4_X1   g402(.A1(new_n326), .A2(new_n582), .A3(new_n281), .A4(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT41), .B(G113), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G15));
  INV_X1    g405(.A(new_n588), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n327), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n542), .A2(new_n533), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G116), .ZN(G18));
  NAND4_X1  g410(.A1(new_n586), .A2(new_n432), .A3(new_n435), .A4(new_n587), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n515), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n281), .A2(new_n551), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G119), .ZN(G21));
  NOR2_X1   g416(.A1(G472), .A2(G902), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT99), .B(new_n271), .C1(new_n267), .C2(new_n249), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n274), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT28), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n263), .A2(new_n265), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(new_n260), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n256), .B1(new_n608), .B2(new_n232), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT99), .B1(new_n609), .B2(new_n271), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n603), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n520), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n533), .ZN(new_n614));
  OAI211_X1 g428(.A(KEYINPUT100), .B(new_n603), .C1(new_n605), .C2(new_n610), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n326), .A2(new_n613), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n592), .A2(new_n573), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G122), .ZN(G24));
  NOR2_X1   g433(.A1(new_n597), .A2(new_n578), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(new_n551), .A3(new_n615), .A4(new_n613), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G125), .ZN(G27));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT42), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n430), .A2(new_n401), .A3(new_n431), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n435), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n399), .B(KEYINPUT101), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n397), .B2(G469), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n628), .B1(new_n631), .B2(new_n391), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI211_X1 g448(.A(KEYINPUT102), .B(new_n628), .C1(new_n631), .C2(new_n391), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n391), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n435), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n632), .A2(new_n633), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n640), .A4(new_n627), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n624), .B(new_n578), .C1(new_n636), .C2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n326), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n279), .A2(KEYINPUT105), .A3(new_n280), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n277), .A2(new_n645), .A3(new_n278), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n644), .B2(new_n646), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n643), .B1(new_n649), .B2(new_n270), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n623), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n626), .B1(new_n638), .B2(KEYINPUT102), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT103), .B1(new_n652), .B2(new_n640), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n634), .A2(new_n625), .A3(new_n635), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT42), .B(new_n579), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n644), .A2(new_n646), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n270), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n326), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n655), .A2(new_n661), .A3(KEYINPUT107), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n327), .B1(new_n636), .B2(new_n641), .ZN(new_n663));
  AOI211_X1 g477(.A(KEYINPUT104), .B(KEYINPUT42), .C1(new_n663), .C2(new_n579), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n328), .B(new_n579), .C1(new_n653), .C2(new_n654), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(new_n666), .B2(new_n624), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n651), .A2(new_n662), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT108), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n206), .ZN(G33));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n557), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G134), .ZN(G36));
  INV_X1    g486(.A(new_n391), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n397), .B(KEYINPUT45), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT109), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n629), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n679), .B1(new_n678), .B2(new_n677), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n435), .A3(new_n560), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n531), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n470), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT43), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n685), .B(new_n551), .C1(new_n519), .C2(new_n520), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n626), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n682), .B(new_n688), .C1(new_n687), .C2(new_n686), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT110), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G137), .ZN(G39));
  NOR2_X1   g505(.A1(new_n326), .A2(new_n626), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n281), .A2(new_n578), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n680), .A2(KEYINPUT47), .A3(new_n435), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT47), .B1(new_n680), .B2(new_n435), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n692), .B(new_n693), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G140), .ZN(G42));
  NOR3_X1   g512(.A1(new_n592), .A2(new_n474), .A3(new_n626), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n685), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n650), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT48), .ZN(new_n703));
  INV_X1    g517(.A(new_n474), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n685), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n613), .A2(new_n615), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n706), .A2(new_n326), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n598), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n699), .A2(new_n326), .A3(new_n572), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n470), .A3(new_n531), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n703), .A2(new_n473), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n713), .B(KEYINPUT115), .Z(new_n714));
  INV_X1    g528(.A(new_n696), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n586), .A2(new_n587), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n628), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n694), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n627), .A3(new_n709), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n701), .A2(new_n551), .A3(new_n706), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n711), .A2(new_n471), .A3(new_n683), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OR3_X1    g536(.A1(new_n567), .A2(new_n401), .A3(new_n592), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT113), .B1(new_n708), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT50), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(KEYINPUT50), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n722), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT51), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(KEYINPUT51), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n729), .A2(KEYINPUT51), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n719), .A2(new_n727), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n714), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n532), .B1(new_n514), .B2(new_n470), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n614), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n516), .B(new_n552), .C1(new_n522), .C2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n579), .B(new_n706), .C1(new_n653), .C2(new_n654), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n469), .B1(new_n541), .B2(new_n540), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n518), .A2(new_n627), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n281), .A3(new_n514), .A4(new_n555), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n739), .B1(new_n744), .B2(new_n551), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n589), .B1(new_n616), .B2(new_n617), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n593), .A2(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n538), .A2(new_n432), .A3(new_n470), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n550), .A2(new_n317), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n556), .B(new_n749), .C1(new_n323), .C2(new_n325), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n748), .A2(new_n750), .A3(new_n571), .A4(new_n632), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n558), .A2(new_n621), .A3(new_n580), .A4(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n746), .B(new_n747), .C1(new_n752), .C2(KEYINPUT52), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(KEYINPUT52), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n668), .A2(new_n745), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n671), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n668), .A2(new_n759), .A3(new_n754), .A4(new_n755), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT53), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n755), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n327), .B(new_n578), .C1(new_n636), .C2(new_n641), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT104), .B1(new_n764), .B2(KEYINPUT42), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n666), .A2(new_n665), .A3(new_n624), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n642), .A2(new_n623), .A3(new_n650), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT107), .B1(new_n655), .B2(new_n661), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n763), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n671), .A3(new_n745), .A4(new_n754), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(KEYINPUT53), .B2(new_n760), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n736), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n753), .B(new_n763), .C1(new_n767), .C2(new_n770), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n671), .A4(new_n745), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT53), .B1(new_n756), .B2(new_n757), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n735), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n758), .A2(new_n761), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n772), .A2(KEYINPUT53), .A3(new_n760), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT54), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT54), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT112), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n734), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n472), .A2(new_n309), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n734), .B(KEYINPUT116), .C1(new_n780), .C2(new_n785), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n716), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n567), .A2(new_n643), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n716), .A2(new_n792), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n572), .A2(new_n684), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n401), .A3(new_n435), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n791), .A2(new_n797), .ZN(G75));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n762), .A2(new_n773), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(G902), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT118), .B(new_n799), .C1(new_n801), .C2(new_n243), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n422), .A2(new_n425), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n423), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n309), .A2(G952), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT119), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n799), .B1(new_n801), .B2(new_n243), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n802), .A2(new_n806), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n807), .A2(new_n812), .A3(new_n813), .ZN(G51));
  NAND2_X1  g628(.A1(new_n781), .A2(new_n782), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(KEYINPUT120), .A3(new_n736), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT120), .B1(new_n815), .B2(new_n736), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n774), .A3(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n629), .B(KEYINPUT57), .Z(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n583), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n801), .A2(new_n676), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n808), .B1(new_n821), .B2(new_n822), .ZN(G54));
  NAND4_X1  g637(.A1(new_n800), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n456), .A2(new_n459), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n824), .A2(new_n826), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n827), .A2(new_n828), .A3(new_n808), .ZN(G60));
  NAND3_X1  g643(.A1(new_n774), .A2(new_n735), .A3(new_n779), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT112), .B1(new_n783), .B2(new_n784), .ZN(new_n831));
  XNOR2_X1  g645(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n530), .B(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n523), .A2(new_n525), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n809), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n836), .A2(new_n833), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n818), .B2(new_n840), .ZN(G63));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n842));
  NAND2_X1  g656(.A1(G217), .A2(G902), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT60), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n800), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n809), .B1(new_n845), .B2(new_n314), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n846), .A2(new_n847), .B1(new_n550), .B2(new_n845), .ZN(new_n848));
  AOI211_X1 g662(.A(KEYINPUT122), .B(new_n809), .C1(new_n845), .C2(new_n314), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n845), .A2(new_n314), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n842), .B1(new_n851), .B2(KEYINPUT123), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n845), .A2(new_n550), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n314), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n856), .A3(new_n838), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n850), .A2(new_n857), .ZN(G66));
  AOI21_X1  g672(.A(new_n309), .B1(new_n477), .B2(G224), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n746), .A2(new_n747), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n739), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n309), .ZN(new_n863));
  INV_X1    g677(.A(G898), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n803), .B1(new_n864), .B2(G953), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n863), .B(new_n865), .ZN(G69));
  AND3_X1   g680(.A1(new_n558), .A2(new_n621), .A3(new_n580), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n575), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT62), .Z(new_n869));
  NAND4_X1  g683(.A1(new_n328), .A2(new_n561), .A3(new_n627), .A4(new_n737), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT124), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n697), .A3(new_n689), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n309), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n254), .B(new_n450), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n309), .A2(G900), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n680), .A2(new_n435), .A3(new_n560), .A4(new_n748), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n877), .B1(new_n878), .B2(new_n661), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n697), .A2(new_n689), .A3(new_n867), .A4(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n877), .A3(new_n661), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n668), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n757), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT127), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n876), .B1(new_n887), .B2(new_n309), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n875), .B1(new_n888), .B2(new_n874), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT125), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n889), .B(new_n891), .ZN(G72));
  NAND3_X1  g706(.A1(new_n882), .A2(new_n861), .A3(new_n886), .ZN(new_n893));
  NAND2_X1  g707(.A1(G472), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT63), .Z(new_n895));
  AOI211_X1 g709(.A(new_n255), .B(new_n249), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n872), .B2(new_n862), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n808), .B1(new_n897), .B2(new_n569), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n255), .B(new_n256), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n777), .A2(new_n778), .A3(new_n895), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n896), .A2(new_n901), .ZN(G57));
endmodule


