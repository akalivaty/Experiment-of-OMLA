//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G137), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n190), .A2(G137), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(G143), .B2(new_n201), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(G128), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n191), .A2(new_n195), .A3(new_n193), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n196), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n202), .A2(new_n204), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  OR2_X1    g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(KEYINPUT64), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n220), .A2(new_n223), .B1(new_n210), .B2(new_n221), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n217), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT65), .B1(new_n217), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n214), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G119), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT66), .A3(G116), .ZN(new_n229));
  INV_X1    g043(.A(G116), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G119), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n230), .B2(G119), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n232), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n231), .A3(new_n229), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n239), .B2(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n233), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n227), .A2(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n217), .A2(new_n224), .B1(new_n200), .B2(new_n213), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n238), .A2(new_n240), .B1(new_n233), .B2(new_n239), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(KEYINPUT28), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n246), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G237), .A2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(KEYINPUT27), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT26), .B(G101), .Z(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n217), .A2(new_n224), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n214), .A3(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n243), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT30), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(new_n227), .ZN(new_n262));
  INV_X1    g076(.A(new_n256), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n257), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n246), .B1(new_n245), .B2(KEYINPUT30), .ZN(new_n266));
  INV_X1    g080(.A(new_n214), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n217), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n271), .B2(KEYINPUT30), .ZN(new_n272));
  INV_X1    g086(.A(new_n264), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(KEYINPUT31), .A3(new_n273), .ZN(new_n274));
  AOI221_X4 g088(.A(new_n188), .B1(new_n251), .B2(new_n256), .C1(new_n265), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n265), .A2(new_n274), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n251), .A2(new_n256), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT68), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n187), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n262), .A2(new_n257), .A3(new_n264), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT31), .B1(new_n272), .B2(new_n273), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n188), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(KEYINPUT68), .A3(new_n277), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n187), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n281), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n187), .A2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT74), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n291), .C1(new_n286), .C2(new_n287), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n244), .A2(new_n263), .A3(new_n247), .A4(new_n250), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n258), .A2(new_n214), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(new_n243), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n227), .A2(new_n261), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n266), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT70), .B1(new_n303), .B2(new_n263), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n272), .A2(new_n248), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n256), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n299), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n256), .A2(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n250), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n248), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n243), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n246), .A2(KEYINPUT71), .A3(new_n258), .A4(new_n214), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n310), .B1(new_n315), .B2(KEYINPUT28), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT72), .B1(new_n316), .B2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n314), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT71), .B1(new_n245), .B2(new_n246), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT28), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n250), .A3(new_n309), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G472), .B1(new_n308), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n299), .A2(new_n304), .A3(new_n307), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n317), .A3(new_n324), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT73), .A3(G472), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n290), .A2(new_n296), .A3(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n334));
  INV_X1    g148(.A(G107), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G104), .ZN(new_n336));
  AND2_X1   g150(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  INV_X1    g153(.A(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G107), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(G107), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n338), .A2(new_n339), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n335), .B2(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n336), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n341), .A2(new_n346), .ZN(new_n349));
  OAI21_X1  g163(.A(G101), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n213), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT82), .B1(new_n351), .B2(KEYINPUT10), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n213), .A2(new_n345), .A3(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n217), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n345), .A2(new_n350), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(KEYINPUT83), .A3(KEYINPUT10), .A4(new_n213), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n213), .A2(KEYINPUT10), .A3(new_n345), .A4(new_n350), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n344), .A2(new_n341), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n343), .B1(new_n342), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G101), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT4), .A3(new_n345), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(G101), .C1(new_n365), .C2(new_n367), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n224), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n357), .A2(new_n358), .A3(new_n364), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G953), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G227), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT79), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n361), .A2(new_n362), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n361), .A2(new_n362), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n372), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n217), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT84), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT84), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n217), .C1(new_n382), .C2(new_n385), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n379), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n359), .A2(new_n213), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n217), .B1(new_n391), .B2(new_n351), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT12), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT12), .B(new_n217), .C1(new_n391), .C2(new_n351), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n378), .B1(new_n396), .B2(new_n373), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT85), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n373), .A2(new_n378), .ZN(new_n399));
  INV_X1    g213(.A(new_n389), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n364), .B(new_n372), .C1(new_n384), .C2(new_n383), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n388), .B1(new_n401), .B2(new_n217), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n399), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n404));
  INV_X1    g218(.A(new_n397), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n406), .A3(G469), .ZN(new_n407));
  INV_X1    g221(.A(G469), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n387), .A2(new_n389), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n378), .B1(new_n409), .B2(new_n373), .ZN(new_n410));
  INV_X1    g224(.A(new_n396), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n379), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n408), .B(new_n323), .C1(new_n410), .C2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(G469), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G214), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n232), .A2(KEYINPUT5), .A3(new_n237), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n228), .A2(G116), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n418), .B(G113), .C1(KEYINPUT5), .C2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n359), .A3(new_n241), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n369), .A2(new_n371), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n246), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n421), .B(new_n424), .C1(new_n422), .C2(new_n246), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n213), .A2(G125), .ZN(new_n429));
  INV_X1    g243(.A(G125), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n224), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n374), .A2(G224), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n423), .A2(new_n435), .A3(new_n425), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n428), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n433), .A2(KEYINPUT7), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n431), .B1(new_n440), .B2(new_n429), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT86), .B1(new_n213), .B2(G125), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n439), .B1(new_n443), .B2(KEYINPUT87), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n424), .B(KEYINPUT8), .ZN(new_n445));
  INV_X1    g259(.A(new_n421), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n359), .B1(new_n241), .B2(new_n420), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n439), .A2(KEYINPUT87), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n444), .A2(new_n427), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n437), .A2(new_n450), .A3(new_n323), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n437), .A2(new_n450), .A3(new_n323), .A4(new_n452), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n417), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT9), .B(G234), .ZN(new_n457));
  OAI21_X1  g271(.A(G221), .B1(new_n457), .B2(G902), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n415), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI211_X1 g273(.A(KEYINPUT13), .B(new_n190), .C1(new_n208), .C2(G143), .ZN(new_n460));
  XNOR2_X1  g274(.A(G128), .B(G143), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n461), .A2(G134), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(G134), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR4_X1   g278(.A1(new_n208), .A2(new_n190), .A3(KEYINPUT13), .A4(G143), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n466));
  INV_X1    g280(.A(G122), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G116), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n230), .A2(G122), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n335), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n469), .A3(new_n335), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(KEYINPUT94), .A3(new_n470), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n464), .A2(new_n465), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n462), .A2(new_n463), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n469), .A2(KEYINPUT14), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n468), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G107), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n474), .A2(KEYINPUT95), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n474), .A2(KEYINPUT95), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G217), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n457), .A2(new_n486), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n488), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(KEYINPUT96), .A3(new_n323), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G478), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n491), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT93), .A2(KEYINPUT20), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(KEYINPUT93), .A2(KEYINPUT20), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G140), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G125), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n430), .A2(G140), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT88), .ZN(new_n504));
  XNOR2_X1  g318(.A(G125), .B(G140), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n507), .A3(G146), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n201), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n374), .A3(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n203), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n252), .A2(G143), .A3(G214), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n515), .B(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n505), .A2(KEYINPUT16), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n521));
  AOI21_X1  g335(.A(G146), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n520), .A2(G146), .A3(new_n521), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(KEYINPUT77), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n194), .B1(new_n513), .B2(new_n514), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n513), .A2(new_n194), .A3(new_n514), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(KEYINPUT17), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n524), .A2(new_n525), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(G113), .B(G122), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(G104), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT92), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n519), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n534), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n510), .A2(new_n518), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT19), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n505), .B2(new_n541), .ZN(new_n542));
  AND4_X1   g356(.A1(new_n540), .A2(new_n501), .A3(new_n502), .A4(new_n541), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT19), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT89), .A4(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n201), .ZN(new_n550));
  INV_X1    g364(.A(new_n529), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n523), .B1(new_n551), .B2(new_n526), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n539), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n538), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n552), .B1(new_n549), .B2(new_n201), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT91), .B1(new_n557), .B2(new_n539), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n537), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(G475), .A2(G902), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n499), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(G146), .B(new_n544), .C1(new_n547), .C2(new_n548), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n519), .B(new_n555), .C1(new_n562), .C2(new_n552), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(new_n534), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n564), .B2(new_n536), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n497), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n538), .B1(new_n519), .B2(new_n532), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n323), .B1(new_n537), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G475), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n495), .A2(new_n561), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(G234), .A2(G237), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(G902), .A3(G953), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(KEYINPUT97), .Z(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT21), .B(G898), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G952), .ZN(new_n576));
  AOI211_X1 g390(.A(G953), .B(new_n576), .C1(G234), .C2(G237), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT98), .B1(new_n570), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n499), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n569), .B1(new_n565), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n496), .B(new_n560), .C1(new_n564), .C2(new_n536), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n579), .A4(new_n495), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n486), .B1(G234), .B2(new_n323), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n524), .A2(new_n525), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT24), .B(G110), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT75), .ZN(new_n593));
  XNOR2_X1  g407(.A(G119), .B(G128), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT23), .B1(new_n208), .B2(G119), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT76), .B1(new_n208), .B2(G119), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n593), .A2(new_n594), .B1(new_n597), .B2(G110), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n593), .A2(new_n594), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n597), .A2(G110), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n523), .B(new_n509), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT22), .B(G137), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n374), .A2(G221), .A3(G234), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n599), .B2(new_n602), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT25), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n599), .A2(new_n602), .ZN(new_n612));
  INV_X1    g426(.A(new_n605), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n606), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n611), .B1(new_n615), .B2(G902), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n590), .B1(new_n610), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n589), .A2(G902), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT78), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n609), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n333), .A2(new_n459), .A3(new_n588), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  OAI21_X1  g436(.A(new_n323), .B1(new_n275), .B2(new_n278), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G472), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n281), .A2(new_n624), .A3(new_n289), .A4(new_n620), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n415), .A2(new_n458), .ZN(new_n626));
  INV_X1    g440(.A(new_n456), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n476), .B2(new_n484), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n488), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT33), .B1(new_n629), .B2(new_n488), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n489), .A2(new_n634), .A3(new_n490), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n487), .B1(new_n485), .B2(new_n628), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT33), .A4(new_n630), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n492), .A2(G902), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n633), .A2(new_n635), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n489), .A2(new_n323), .A3(new_n490), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n492), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n583), .B2(new_n584), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n579), .ZN(new_n646));
  NOR4_X1   g460(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  XOR2_X1   g464(.A(new_n579), .B(KEYINPUT102), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n417), .B(new_n652), .C1(new_n454), .C2(new_n455), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n491), .B(new_n493), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n654), .A3(new_n585), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n625), .A2(new_n626), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G107), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT103), .B(KEYINPUT35), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  AND2_X1   g473(.A1(new_n281), .A2(new_n289), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n613), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n612), .B(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n619), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n617), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n660), .A2(KEYINPUT104), .A3(new_n624), .A4(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n281), .A2(new_n624), .A3(new_n289), .A4(new_n664), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n668), .A3(new_n588), .A4(new_n459), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n669), .B(new_n671), .ZN(G12));
  NAND3_X1  g486(.A1(new_n561), .A2(new_n566), .A3(new_n569), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n573), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n578), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n673), .A2(new_n495), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n333), .A2(new_n459), .A3(new_n664), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  AND2_X1   g494(.A1(new_n415), .A2(new_n458), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n676), .B(KEYINPUT39), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT40), .Z(new_n684));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n281), .A2(new_n282), .A3(new_n289), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n292), .B1(new_n275), .B2(new_n278), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n294), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n262), .A2(new_n264), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n315), .A2(new_n256), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n315), .A2(KEYINPUT106), .A3(new_n256), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n323), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(KEYINPUT107), .B(new_n689), .C1(new_n692), .C2(new_n693), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n288), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n688), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n685), .B1(new_n686), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n688), .A2(new_n698), .A3(new_n699), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT108), .A3(new_n290), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n454), .A2(new_n455), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT38), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n673), .A2(new_n654), .ZN(new_n707));
  NOR4_X1   g521(.A1(new_n706), .A2(new_n417), .A3(new_n664), .A4(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n684), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n203), .ZN(G45));
  OAI211_X1 g524(.A(new_n643), .B(new_n676), .C1(new_n583), .C2(new_n584), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n333), .A2(new_n459), .A3(new_n664), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  INV_X1    g528(.A(new_n620), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n330), .A2(KEYINPUT73), .A3(G472), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT73), .B1(new_n330), .B2(G472), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n688), .A2(new_n699), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n715), .B1(new_n720), .B2(new_n290), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n373), .B1(new_n400), .B2(new_n402), .ZN(new_n722));
  INV_X1    g536(.A(new_n378), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n412), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(G469), .B1(new_n724), .B2(G902), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n456), .A3(new_n413), .A4(new_n458), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n646), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND3_X1  g544(.A1(new_n725), .A2(new_n458), .A3(new_n413), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n655), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  AOI21_X1  g548(.A(new_n726), .B1(new_n587), .B2(new_n581), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n333), .A3(new_n664), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  XOR2_X1   g551(.A(KEYINPUT109), .B(G472), .Z(new_n738));
  NAND2_X1  g552(.A1(new_n623), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n320), .A2(new_n250), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n276), .B1(new_n263), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n187), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n620), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n456), .A2(new_n654), .A3(new_n673), .A4(new_n651), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n743), .A2(new_n731), .A3(new_n744), .A4(KEYINPUT110), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n731), .A2(new_n744), .ZN(new_n747));
  INV_X1    g561(.A(new_n743), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n467), .ZN(G24));
  AOI22_X1  g565(.A1(new_n623), .A2(new_n738), .B1(new_n187), .B2(new_n741), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n752), .A2(new_n664), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n711), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n673), .A2(KEYINPUT111), .A3(new_n643), .A4(new_n676), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n726), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n753), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  AOI22_X1  g574(.A1(new_n279), .A2(new_n282), .B1(new_n288), .B2(new_n292), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n717), .B2(new_n716), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(new_n762), .A3(new_n620), .ZN(new_n763));
  INV_X1    g577(.A(new_n458), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n705), .A2(new_n417), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n414), .B(KEYINPUT112), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n397), .B1(new_n409), .B2(new_n399), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(G469), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n413), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n766), .B1(new_n413), .B2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n765), .ZN(new_n775));
  INV_X1    g589(.A(new_n772), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n413), .A2(new_n766), .A3(new_n770), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n755), .A2(new_n756), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(KEYINPUT42), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n778), .A2(new_n333), .A3(new_n780), .A4(new_n620), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT114), .B(G131), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G33));
  NAND4_X1  g598(.A1(new_n778), .A2(new_n333), .A3(new_n620), .A4(new_n678), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  NOR2_X1   g600(.A1(new_n705), .A2(new_n417), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n643), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n673), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n281), .A2(new_n624), .A3(new_n289), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n664), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT44), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  INV_X1    g610(.A(new_n413), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n398), .B2(new_n406), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(G469), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n767), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n458), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n682), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT115), .B(G137), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G39));
  NOR2_X1   g623(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n458), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n333), .A2(new_n620), .A3(new_n711), .A4(new_n788), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G140), .ZN(G42));
  NAND2_X1  g629(.A1(new_n725), .A2(new_n413), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT49), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n764), .A2(new_n417), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n706), .A2(new_n620), .A3(new_n818), .A4(new_n790), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n704), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n791), .A2(new_n577), .ZN(new_n821));
  INV_X1    g635(.A(new_n731), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n787), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n715), .B1(new_n332), .B2(new_n761), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT48), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n704), .A2(new_n715), .A3(new_n578), .A4(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n645), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n743), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n576), .B(G953), .C1(new_n830), .C2(new_n758), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n706), .A2(new_n417), .A3(new_n822), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(KEYINPUT50), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(KEYINPUT50), .B1(new_n753), .B2(new_n824), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n585), .A3(new_n789), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n816), .A2(new_n458), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n812), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n830), .A2(new_n787), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n839), .B(new_n840), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n810), .A2(new_n811), .ZN(new_n845));
  INV_X1    g659(.A(new_n841), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT51), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n832), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n627), .A2(new_n707), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n617), .A2(new_n663), .A3(new_n764), .A4(new_n677), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n851), .B(new_n852), .C1(new_n771), .C2(new_n772), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n686), .A2(new_n700), .A3(new_n685), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT108), .B1(new_n702), .B2(new_n290), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n679), .A3(new_n713), .A4(new_n759), .ZN(new_n858));
  XNOR2_X1  g672(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n679), .A2(new_n759), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n713), .A4(new_n857), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n459), .A2(new_n588), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n666), .B(KEYINPUT104), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n868), .B2(new_n721), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n743), .A2(new_n731), .A3(new_n744), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n746), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n644), .B1(new_n495), .B2(new_n673), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n653), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n625), .A2(new_n626), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n617), .A2(new_n663), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n720), .B2(new_n290), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n735), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n333), .B(new_n620), .C1(new_n732), .C2(new_n727), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n869), .A2(new_n871), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n752), .A2(new_n755), .A3(new_n664), .A4(new_n756), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n773), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n454), .A2(new_n416), .A3(new_n455), .A4(new_n676), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT116), .B1(new_n570), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n570), .A2(new_n882), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n626), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n881), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n888), .A2(new_n774), .A3(new_n781), .A4(new_n785), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n866), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n669), .B(new_n621), .C1(new_n745), .C2(new_n749), .ZN(new_n893));
  INV_X1    g707(.A(new_n874), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n878), .A3(new_n736), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n886), .A2(new_n883), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n333), .A3(new_n681), .A4(new_n664), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n778), .A2(new_n753), .A3(new_n757), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n785), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n782), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n892), .A2(new_n896), .A3(new_n901), .A4(new_n864), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT53), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n891), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n890), .A2(KEYINPUT53), .A3(new_n864), .A4(new_n861), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n850), .A2(new_n905), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n576), .A2(new_n374), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(KEYINPUT119), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n820), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n374), .A2(G952), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n323), .B1(new_n906), .B2(new_n907), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n918), .B2(G210), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n428), .A2(new_n436), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n434), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n917), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n919), .A2(new_n922), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n919), .A2(KEYINPUT120), .A3(new_n922), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n908), .B(KEYINPUT54), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n767), .B(KEYINPUT121), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT57), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n410), .B2(new_n412), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n798), .A2(new_n800), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n916), .B1(new_n933), .B2(new_n935), .ZN(G54));
  AND3_X1   g750(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  INV_X1    g751(.A(new_n559), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n917), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n938), .B2(new_n937), .ZN(G60));
  AND3_X1   g754(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n941));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n929), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n909), .A2(new_n905), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n945), .B2(new_n943), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n946), .A3(new_n916), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n908), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(KEYINPUT122), .A3(new_n615), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n906), .B2(new_n907), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n609), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n916), .B1(new_n954), .B2(new_n662), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n952), .A2(new_n955), .A3(new_n956), .A4(KEYINPUT61), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n853), .B1(new_n701), .B2(new_n703), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n333), .A2(new_n459), .A3(new_n664), .A4(new_n712), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n863), .B1(new_n962), .B2(new_n862), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT53), .B1(new_n964), .B2(new_n890), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n669), .A2(new_n621), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n750), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n774), .A2(new_n781), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n894), .A2(new_n878), .A3(new_n736), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n785), .A2(new_n898), .A3(new_n899), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n967), .A2(new_n968), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n865), .A2(new_n971), .A3(new_n903), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n662), .B(new_n950), .C1(new_n965), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n917), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n954), .A2(new_n609), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n958), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n957), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n957), .A2(new_n976), .A3(KEYINPUT123), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G66));
  INV_X1    g795(.A(G224), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n574), .A2(new_n982), .A3(new_n374), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n896), .B2(new_n374), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n920), .B1(G898), .B2(new_n374), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(G69));
  NAND2_X1  g800(.A1(new_n862), .A2(new_n713), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n709), .A2(KEYINPUT62), .A3(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n683), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n721), .A2(new_n989), .A3(new_n787), .A4(new_n872), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(new_n807), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT62), .B1(new_n709), .B2(new_n987), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n988), .A2(new_n992), .A3(new_n814), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n549), .B(KEYINPUT124), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n302), .A2(new_n259), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n999), .B(new_n1000), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n374), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n806), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n825), .A2(new_n851), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n812), .A2(new_n813), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n807), .A2(new_n987), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1007), .A2(KEYINPUT127), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(KEYINPUT127), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n968), .A2(new_n785), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n374), .ZN(new_n1012));
  INV_X1    g826(.A(G227), .ZN(new_n1013));
  OAI22_X1  g827(.A1(new_n1010), .A2(new_n1012), .B1(new_n1013), .B2(new_n374), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n1001), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n674), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1003), .B(new_n1015), .C1(new_n374), .C2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(new_n305), .A2(new_n263), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n996), .A2(new_n997), .A3(new_n896), .ZN(new_n1019));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  AOI21_X1  g835(.A(new_n1018), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1011), .A2(new_n896), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1021), .B1(new_n1010), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n256), .A3(new_n303), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n304), .A2(new_n307), .ZN(new_n1026));
  OAI221_X1 g840(.A(new_n1021), .B1(new_n689), .B2(new_n1026), .C1(new_n891), .C2(new_n904), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1025), .A2(new_n917), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1022), .A2(new_n1028), .ZN(G57));
endmodule


