//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AND2_X1   g0003(.A1(KEYINPUT64), .A2(G77), .ZN(new_n204));
  NOR2_X1   g0004(.A1(KEYINPUT64), .A2(G77), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G58), .A2(G232), .ZN(new_n212));
  NAND4_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n203), .B1(new_n208), .B2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT65), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n214), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT67), .Z(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n203), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT0), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n223), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n218), .A2(new_n220), .A3(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT68), .Z(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT70), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT71), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n251), .A2(new_n253), .A3(new_n225), .A4(G87), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT22), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT22), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(new_n225), .A4(G87), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT23), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(new_n225), .B2(G107), .ZN(new_n261));
  INV_X1    g0061(.A(G107), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(KEYINPUT23), .A3(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G116), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n250), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n225), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n259), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n203), .B2(new_n250), .ZN(new_n274));
  NAND4_X1  g0074(.A1(KEYINPUT72), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(new_n224), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n259), .A2(KEYINPUT24), .A3(new_n269), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n272), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n275), .A2(new_n224), .ZN(new_n279));
  INV_X1    g0079(.A(G1), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G13), .A3(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n250), .A2(G1), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n279), .A2(new_n281), .A3(new_n274), .A4(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n262), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n281), .A2(G107), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT25), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT96), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n286), .B(KEYINPUT25), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT96), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n290), .B(new_n291), .C1(new_n262), .C2(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n278), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT97), .ZN(new_n295));
  MUX2_X1   g0095(.A(G250), .B(G257), .S(G1698), .Z(new_n296));
  AOI22_X1  g0096(.A1(new_n296), .A2(new_n256), .B1(G33), .B2(G294), .ZN(new_n297));
  AND2_X1   g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  NAND2_X1  g0103(.A1(KEYINPUT5), .A2(G41), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT5), .A2(G41), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(G33), .A2(G41), .ZN(new_n308));
  OAI21_X1  g0108(.A(G274), .B1(new_n308), .B2(new_n224), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT90), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n280), .A2(G45), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT5), .ZN(new_n312));
  INV_X1    g0112(.A(G41), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n304), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT90), .ZN(new_n316));
  INV_X1    g0116(.A(G274), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n298), .B2(new_n299), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n307), .A2(G264), .A3(new_n300), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n301), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n301), .A2(G179), .A3(new_n320), .A4(new_n321), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT97), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n278), .A2(new_n293), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n295), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(G200), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n301), .A2(G190), .A3(new_n320), .A4(new_n321), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n329), .A2(new_n278), .A3(new_n293), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n280), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n274), .A2(new_n224), .A3(new_n281), .A4(new_n275), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(new_n281), .B2(new_n335), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n251), .A2(new_n253), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n340), .B2(new_n225), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n342), .B(G20), .C1(new_n251), .C2(new_n253), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT81), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n225), .A2(new_n250), .ZN(new_n346));
  INV_X1    g0146(.A(G159), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(G20), .A2(G33), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT81), .A3(G159), .ZN(new_n350));
  XNOR2_X1  g0150(.A(G58), .B(G68), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n348), .A2(new_n350), .B1(G20), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT16), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT82), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n342), .B1(new_n256), .B2(G20), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(new_n350), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(G20), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT82), .B(new_n354), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n355), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n276), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n358), .A2(KEYINPUT80), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT80), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n340), .A2(new_n368), .A3(KEYINPUT7), .A4(new_n225), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n357), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n362), .B1(new_n370), .B2(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n339), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  INV_X1    g0174(.A(G1698), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n251), .A2(new_n253), .A3(G223), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT83), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n256), .A2(KEYINPUT83), .A3(G223), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G33), .A2(G87), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n256), .A2(G226), .A3(G1698), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n308), .A2(new_n224), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n280), .B1(G41), .B2(G45), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n318), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n300), .A2(G232), .A3(new_n385), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n374), .B1(new_n384), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT73), .B(G179), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n392), .B(new_n389), .C1(new_n382), .C2(new_n383), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT84), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n392), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n384), .A2(new_n395), .A3(new_n390), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT84), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n382), .B2(new_n383), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n397), .C1(new_n374), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n373), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n343), .A2(new_n368), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n369), .A2(new_n357), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n352), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n354), .B1(new_n359), .B2(new_n362), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT82), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n405), .A2(new_n408), .A3(new_n276), .A4(new_n363), .ZN(new_n409));
  INV_X1    g0209(.A(new_n339), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n394), .A4(new_n399), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT85), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT85), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n401), .A2(new_n416), .A3(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n398), .A2(G190), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n398), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n409), .A2(new_n418), .A3(new_n410), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n420), .A2(new_n418), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n424), .A2(new_n409), .A3(KEYINPUT17), .A4(new_n410), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n415), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n300), .A2(new_n385), .ZN(new_n429));
  INV_X1    g0229(.A(G238), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n387), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n256), .A2(G226), .A3(new_n375), .ZN(new_n432));
  INV_X1    g0232(.A(G97), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n256), .A2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G232), .ZN(new_n435));
  OAI221_X1 g0235(.A(new_n432), .B1(new_n250), .B2(new_n433), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n431), .B1(new_n436), .B2(new_n383), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  OAI21_X1  g0241(.A(G169), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT78), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT13), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n437), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n437), .B2(new_n447), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(G179), .A4(new_n439), .ZN(new_n450));
  OAI211_X1 g0250(.A(G169), .B(new_n443), .C1(new_n440), .C2(new_n441), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n281), .A2(G68), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT12), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT11), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n349), .A2(G50), .B1(G20), .B2(new_n356), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n250), .A2(G20), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G77), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n276), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n463));
  INV_X1    g0263(.A(new_n338), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G68), .A3(new_n336), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n452), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n448), .A2(new_n449), .A3(G190), .A4(new_n439), .ZN(new_n469));
  OAI21_X1  g0269(.A(G200), .B1(new_n440), .B2(new_n441), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n256), .A2(G222), .A3(new_n375), .ZN(new_n473));
  INV_X1    g0273(.A(G223), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n473), .B1(new_n206), .B2(new_n256), .C1(new_n434), .C2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(new_n383), .ZN(new_n476));
  INV_X1    g0276(.A(G226), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n387), .B1(new_n429), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT9), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n464), .A2(G50), .A3(new_n336), .ZN(new_n481));
  INV_X1    g0281(.A(G150), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n334), .A2(new_n458), .B1(new_n482), .B2(new_n346), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G58), .A2(G68), .ZN(new_n484));
  INV_X1    g0284(.A(G50), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n225), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n276), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n281), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n485), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n479), .A2(G190), .B1(new_n480), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n479), .A2(new_n419), .B1(new_n490), .B2(new_n480), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT10), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n493), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT10), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT15), .B(G87), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(KEYINPUT75), .A3(new_n457), .ZN(new_n501));
  INV_X1    g0301(.A(new_n206), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n335), .A2(new_n349), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT75), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n499), .B2(new_n458), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n276), .B1(new_n206), .B2(new_n488), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n464), .A2(G77), .A3(new_n336), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n340), .A2(G107), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n434), .B2(new_n430), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n340), .A2(new_n435), .A3(G1698), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n383), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT74), .ZN(new_n515));
  INV_X1    g0315(.A(new_n429), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G244), .B1(new_n318), .B2(new_n386), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n514), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n510), .B1(new_n520), .B2(new_n374), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT76), .ZN(new_n522));
  INV_X1    g0322(.A(new_n519), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n525), .B2(new_n392), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n522), .B(new_n392), .C1(new_n518), .C2(new_n519), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n521), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(G190), .B1(new_n518), .B2(new_n519), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n510), .C1(new_n525), .C2(new_n419), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n490), .B1(new_n479), .B2(G169), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n476), .A2(new_n395), .A3(new_n478), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n498), .A2(new_n529), .A3(new_n531), .A4(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n428), .A2(new_n472), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n284), .A2(new_n433), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n281), .A2(G97), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT86), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n346), .B2(new_n459), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n349), .A2(KEYINPUT86), .A3(G77), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  NOR2_X1   g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT87), .B(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n262), .A2(KEYINPUT6), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n546), .A2(KEYINPUT6), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n543), .B1(new_n549), .B2(G20), .ZN(new_n550));
  OAI21_X1  g0350(.A(G107), .B1(new_n341), .B2(new_n343), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n538), .B(new_n539), .C1(new_n552), .C2(new_n276), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n315), .A2(new_n383), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G257), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n320), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n251), .A2(new_n253), .A3(G244), .A4(new_n375), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT88), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n557), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n251), .A2(new_n253), .A3(G250), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G283), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n556), .B1(new_n383), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G190), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n558), .A2(new_n559), .A3(new_n557), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n570), .A2(new_n560), .A3(new_n565), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT89), .B1(new_n571), .B2(new_n300), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT89), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(new_n573), .A3(new_n383), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n556), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n553), .B(new_n569), .C1(new_n575), .C2(new_n419), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n539), .B1(new_n552), .B2(new_n276), .ZN(new_n577));
  INV_X1    g0377(.A(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G97), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n310), .A2(new_n319), .B1(new_n554), .B2(G257), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n571), .B2(new_n300), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n577), .A2(new_n579), .B1(new_n581), .B2(new_n374), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n571), .A2(KEYINPUT89), .A3(new_n300), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n573), .B1(new_n567), .B2(new_n383), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n392), .B(new_n580), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n281), .A2(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n265), .A2(G20), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n433), .A2(KEYINPUT87), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(G33), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n564), .A2(new_n225), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n276), .B(new_n590), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n225), .B(new_n564), .C1(new_n547), .C2(G33), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n276), .A4(new_n590), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n589), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n338), .A2(new_n265), .A3(new_n282), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n375), .A2(G264), .ZN(new_n606));
  NOR2_X1   g0406(.A1(G257), .A2(G1698), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n340), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n383), .B1(new_n256), .B2(G303), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT95), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G303), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n300), .B1(new_n340), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT95), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n256), .B1(new_n607), .B2(new_n606), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n310), .A2(new_n319), .B1(new_n554), .B2(G270), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n605), .B(new_n374), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n617), .A2(G179), .A3(new_n618), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n604), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n374), .B1(new_n617), .B2(new_n618), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n602), .B(new_n589), .C1(new_n598), .C2(new_n600), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n605), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n617), .A2(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  INV_X1    g0427(.A(G190), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n627), .B(new_n624), .C1(new_n628), .C2(new_n626), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT94), .ZN(new_n631));
  INV_X1    g0431(.A(G250), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n280), .B2(G45), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n318), .A2(new_n303), .B1(new_n300), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(G238), .A2(G1698), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n635), .B1(new_n207), .B2(G1698), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n266), .B1(new_n636), .B2(new_n256), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n300), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT93), .B1(new_n638), .B2(new_n628), .ZN(new_n639));
  INV_X1    g0439(.A(new_n635), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n207), .A2(G1698), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n256), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n266), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n383), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT93), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G190), .A4(new_n634), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n639), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n638), .A2(G200), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n500), .A2(new_n281), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n578), .A2(G87), .ZN(new_n653));
  INV_X1    g0453(.A(G87), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n591), .A2(new_n593), .A3(new_n654), .A4(new_n262), .ZN(new_n655));
  NAND3_X1  g0455(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n225), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n251), .A2(new_n253), .A3(new_n225), .A4(G68), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT91), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n256), .A2(KEYINPUT91), .A3(new_n225), .A4(G68), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n591), .A2(new_n593), .ZN(new_n664));
  AOI211_X1 g0464(.A(KEYINPUT92), .B(KEYINPUT19), .C1(new_n664), .C2(new_n457), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n547), .A2(new_n458), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT92), .B1(new_n667), .B2(KEYINPUT19), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n652), .B(new_n653), .C1(new_n669), .C2(new_n366), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n650), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n300), .A2(new_n633), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n309), .B2(new_n311), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n383), .B2(new_n644), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n392), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n638), .A2(new_n374), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n660), .A2(new_n659), .B1(new_n655), .B2(new_n657), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT19), .B1(new_n664), .B2(new_n457), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n662), .B(new_n678), .C1(new_n681), .C2(new_n665), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n651), .B1(new_n682), .B2(new_n276), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n578), .A2(new_n500), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n677), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n631), .B1(new_n671), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n652), .B(new_n684), .C1(new_n669), .C2(new_n366), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n675), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n683), .A2(new_n648), .A3(new_n653), .A4(new_n649), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT94), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n630), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n333), .A2(new_n537), .A3(new_n588), .A4(new_n692), .ZN(G372));
  INV_X1    g0493(.A(new_n414), .ZN(new_n694));
  INV_X1    g0494(.A(new_n529), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(new_n471), .B1(new_n452), .B2(new_n467), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n694), .B1(new_n696), .B2(new_n426), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n534), .B1(new_n697), .B2(new_n498), .ZN(new_n698));
  INV_X1    g0498(.A(new_n537), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n582), .A2(new_n689), .A3(new_n585), .A4(new_n690), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n689), .B1(new_n700), .B2(KEYINPUT26), .ZN(new_n701));
  INV_X1    g0501(.A(new_n586), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n689), .A2(new_n690), .A3(KEYINPUT94), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT94), .B1(new_n689), .B2(new_n690), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n701), .B1(KEYINPUT26), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n689), .A2(new_n331), .A3(new_n690), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n587), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n325), .A2(new_n294), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT98), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n626), .A2(KEYINPUT21), .A3(G169), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n617), .A2(new_n618), .A3(G179), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n624), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT21), .B1(new_n604), .B2(new_n622), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n621), .A2(new_n625), .A3(KEYINPUT98), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n710), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n708), .B1(new_n718), .B2(KEYINPUT99), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT99), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n720), .B(new_n710), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n706), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n698), .B1(new_n699), .B2(new_n723), .ZN(G369));
  NAND3_X1  g0524(.A1(new_n280), .A2(new_n225), .A3(G13), .ZN(new_n725));
  OAI21_X1  g0525(.A(G213), .B1(new_n725), .B2(KEYINPUT27), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n727), .A2(KEYINPUT100), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(KEYINPUT100), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G343), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n295), .A2(new_n327), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n333), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n328), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n732), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n624), .A2(new_n731), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n630), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n716), .A2(new_n717), .A3(new_n739), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n731), .B1(new_n714), .B2(new_n715), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n731), .B(KEYINPUT101), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n332), .A2(new_n746), .B1(new_n709), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(G399));
  INV_X1    g0550(.A(new_n221), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G41), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n655), .A2(G116), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(G1), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n227), .B2(new_n753), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT28), .ZN(new_n757));
  INV_X1    g0557(.A(new_n747), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n692), .A2(new_n333), .A3(new_n588), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n674), .A2(new_n395), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n761), .A2(new_n322), .A3(new_n626), .A4(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n321), .B1(new_n297), .B2(new_n300), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n638), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(G179), .A3(new_n617), .A4(new_n618), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT30), .B1(new_n766), .B2(new_n581), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT30), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n620), .A2(new_n568), .A3(new_n768), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n760), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n732), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT31), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n738), .B1(new_n759), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n722), .A2(new_n758), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT29), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n714), .A2(new_n715), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT102), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n328), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n328), .B2(new_n780), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n671), .A2(new_n685), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n785), .A2(new_n576), .A3(new_n586), .A4(new_n331), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT26), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n685), .B1(new_n700), .B2(KEYINPUT26), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(KEYINPUT29), .B(new_n731), .C1(new_n787), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n776), .B1(new_n779), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n757), .B1(new_n793), .B2(G1), .ZN(G364));
  AND2_X1   g0594(.A1(new_n225), .A2(G13), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n280), .B1(new_n795), .B2(G45), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n752), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n256), .A2(new_n221), .ZN(new_n799));
  INV_X1    g0599(.A(G355), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(G116), .B2(new_n221), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n751), .A2(new_n256), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT103), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n302), .B2(new_n228), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n244), .A2(new_n302), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G13), .A2(G33), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(G20), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n224), .B1(G20), .B2(new_n374), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n798), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n225), .A2(new_n628), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n419), .A2(G179), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n225), .A2(G190), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G179), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G303), .A2(new_n817), .B1(new_n821), .B2(G329), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n815), .A2(new_n818), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n340), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n395), .A2(G20), .A3(G200), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n628), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(G190), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G326), .A2(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n395), .A2(new_n419), .A3(new_n818), .ZN(new_n832));
  INV_X1    g0632(.A(G322), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n395), .A2(new_n419), .A3(new_n814), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n819), .A2(G190), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G20), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n825), .B(new_n835), .C1(G294), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT104), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(G58), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n842), .A2(new_n834), .B1(new_n832), .B2(new_n206), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G50), .B2(new_n827), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n821), .A2(G159), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n845), .A2(KEYINPUT32), .ZN(new_n846));
  INV_X1    g0646(.A(new_n837), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n433), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(KEYINPUT32), .B2(new_n845), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n256), .B1(new_n824), .B2(new_n262), .C1(new_n654), .C2(new_n816), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G68), .B2(new_n828), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n844), .A2(new_n846), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n840), .A2(new_n841), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n813), .B1(new_n853), .B2(new_n810), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n740), .A2(new_n741), .A3(new_n809), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n740), .A2(new_n738), .A3(new_n741), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n743), .B(new_n857), .C1(new_n752), .C2(new_n797), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G396));
  OR3_X1    g0660(.A1(new_n510), .A2(KEYINPUT107), .A3(new_n731), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n531), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n529), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT76), .B1(new_n520), .B2(new_n395), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n527), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT107), .B1(new_n865), .B2(new_n521), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n510), .A2(new_n731), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n863), .B(new_n758), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n722), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n714), .A2(new_n715), .A3(new_n711), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT98), .B1(new_n621), .B2(new_n625), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n709), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n720), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n718), .A2(KEYINPUT99), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n708), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n747), .B1(new_n876), .B2(new_n706), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n870), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n776), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n798), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n881), .B2(new_n880), .ZN(new_n883));
  INV_X1    g0683(.A(new_n810), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n808), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n798), .B1(G77), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n834), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n827), .A2(G303), .B1(new_n887), .B2(G294), .ZN(new_n888));
  INV_X1    g0688(.A(new_n828), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n888), .B1(new_n265), .B2(new_n832), .C1(new_n823), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n340), .B1(new_n820), .B2(new_n831), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n816), .A2(new_n262), .B1(new_n824), .B2(new_n654), .ZN(new_n892));
  OR4_X1    g0692(.A1(new_n848), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(G137), .A2(new_n827), .B1(new_n828), .B2(G150), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT105), .Z(new_n895));
  INV_X1    g0695(.A(new_n832), .ZN(new_n896));
  AOI22_X1  g0696(.A1(G143), .A2(new_n887), .B1(new_n896), .B2(G159), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(KEYINPUT34), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n256), .B1(new_n816), .B2(new_n485), .ZN(new_n899));
  INV_X1    g0699(.A(new_n824), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G68), .ZN(new_n901));
  INV_X1    g0701(.A(G132), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n820), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n899), .B(new_n903), .C1(G58), .C2(new_n837), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT34), .B1(new_n895), .B2(new_n897), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n884), .B1(new_n907), .B2(KEYINPUT106), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n886), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n808), .B2(new_n879), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n883), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(G384));
  OAI211_X1 g0713(.A(G116), .B(new_n226), .C1(new_n549), .C2(KEYINPUT35), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n549), .A2(KEYINPUT35), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(KEYINPUT108), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT36), .Z(new_n919));
  OAI211_X1 g0719(.A(new_n502), .B(new_n228), .C1(new_n842), .C2(new_n356), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n485), .A2(G68), .ZN(new_n921));
  AOI211_X1 g0721(.A(new_n280), .B(G13), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n467), .A2(new_n732), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n468), .A2(new_n471), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n471), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n467), .B(new_n732), .C1(new_n926), .C2(new_n452), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n695), .A2(new_n731), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n929), .B1(new_n870), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n404), .A2(new_n352), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n354), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n339), .B1(new_n372), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n730), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n426), .B1(new_n414), .B2(KEYINPUT85), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(new_n417), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n421), .B1(new_n400), .B2(new_n935), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT37), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n411), .A2(new_n394), .A3(new_n399), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n411), .A2(new_n730), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT37), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n421), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n932), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n942), .A2(new_n946), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n401), .A2(new_n416), .A3(new_n413), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n416), .B1(new_n401), .B2(new_n413), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n950), .A2(new_n951), .A3(new_n426), .ZN(new_n952));
  OAI211_X1 g0752(.A(KEYINPUT38), .B(new_n949), .C1(new_n952), .C2(new_n938), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n931), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n694), .A2(new_n730), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n955), .A2(KEYINPUT109), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n940), .A2(new_n932), .A3(new_n947), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n411), .B(new_n730), .C1(new_n414), .C2(new_n426), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n943), .A2(new_n421), .A3(new_n944), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT37), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n946), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT38), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n959), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n468), .A2(new_n732), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n948), .A2(new_n953), .A3(KEYINPUT39), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n958), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n956), .B1(new_n931), .B2(new_n954), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT109), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n537), .B(new_n792), .C1(new_n877), .C2(KEYINPUT29), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n975), .A2(new_n698), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n974), .B(new_n976), .Z(new_n977));
  AOI21_X1  g0777(.A(new_n878), .B1(new_n925), .B2(new_n927), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n773), .A2(new_n774), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n732), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n759), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT40), .B1(new_n954), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n965), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n953), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n978), .A2(KEYINPUT40), .A3(new_n981), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n537), .A2(new_n981), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n738), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n988), .B2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n977), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n280), .B2(new_n795), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n977), .A2(new_n991), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n923), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT110), .Z(G367));
  NAND2_X1  g0796(.A1(new_n670), .A2(new_n732), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n785), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n685), .A2(new_n670), .A3(new_n732), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n809), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n811), .B1(new_n221), .B2(new_n499), .C1(new_n240), .C2(new_n803), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n1003), .A2(new_n798), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n828), .A2(G159), .B1(new_n887), .B2(G150), .ZN(new_n1005));
  INV_X1    g0805(.A(G143), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n827), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1005), .B1(new_n485), .B2(new_n832), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n847), .A2(new_n356), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n256), .B1(new_n820), .B2(new_n1010), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n816), .A2(new_n842), .B1(new_n824), .B2(new_n206), .ZN(new_n1012));
  NOR4_X1   g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n828), .A2(G294), .B1(new_n887), .B2(G303), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n831), .B2(new_n1007), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT46), .B1(new_n817), .B2(G116), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n262), .B2(new_n847), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n256), .B1(new_n821), .B2(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n547), .B2(new_n824), .C1(new_n823), .C2(new_n832), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT47), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1002), .B(new_n1004), .C1(new_n1023), .C2(new_n884), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n553), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n747), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n576), .A2(new_n586), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT111), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n582), .A2(new_n585), .A3(new_n747), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1028), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT112), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT112), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n745), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(KEYINPUT113), .B(new_n586), .C1(new_n1038), .C2(new_n328), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT113), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1032), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1035), .A2(KEYINPUT112), .A3(new_n1036), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n328), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1041), .B1(new_n1044), .B2(new_n702), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1040), .A2(new_n1045), .A3(new_n758), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n746), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n333), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT42), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT43), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1001), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1046), .A2(new_n1055), .A3(new_n1001), .A4(new_n1051), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1039), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1039), .A3(new_n1059), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1060), .B1(KEYINPUT114), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT45), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1047), .B2(new_n748), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n749), .B(KEYINPUT45), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1047), .A2(KEYINPUT44), .A3(new_n748), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1035), .A2(new_n748), .A3(new_n1036), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT44), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n744), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n734), .A2(new_n736), .A3(new_n746), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n1049), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n742), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n743), .A2(new_n1074), .A3(new_n1049), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1066), .A2(new_n745), .A3(new_n1071), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n793), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n793), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n752), .B(KEYINPUT41), .Z(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n796), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1039), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1053), .B(new_n1056), .C1(new_n1046), .C2(new_n1051), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1059), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT114), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1024), .B1(new_n1062), .B2(new_n1091), .ZN(G387));
  NAND2_X1  g0892(.A1(new_n737), .A2(new_n809), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n236), .A2(new_n302), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(new_n803), .B1(new_n754), .B2(new_n799), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n334), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1096));
  AOI21_X1  g0896(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT50), .B1(new_n334), .B2(G50), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n754), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1095), .A2(new_n1099), .B1(new_n262), .B2(new_n751), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n798), .B1(new_n1100), .B2(new_n812), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n816), .A2(new_n206), .B1(new_n824), .B2(new_n433), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n340), .B(new_n1102), .C1(G150), .C2(new_n821), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n827), .A2(G159), .B1(new_n896), .B2(G68), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n828), .A2(new_n335), .B1(new_n887), .B2(G50), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n500), .A2(new_n837), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n256), .B1(new_n821), .B2(G326), .ZN(new_n1108));
  INV_X1    g0908(.A(G294), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n847), .A2(new_n823), .B1(new_n816), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G303), .A2(new_n896), .B1(new_n887), .B2(G317), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n889), .B2(new_n831), .C1(new_n833), .C2(new_n1007), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT48), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1113), .B2(new_n1112), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT49), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1108), .B1(new_n265), .B2(new_n824), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1107), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1101), .B1(new_n1119), .B2(new_n810), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1078), .A2(new_n797), .B1(new_n1093), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n779), .A2(new_n792), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n881), .A3(new_n1078), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n752), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n793), .A2(new_n1078), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1121), .B1(new_n1124), .B2(new_n1125), .ZN(G393));
  INV_X1    g0926(.A(new_n1079), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n745), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1123), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1080), .A3(new_n752), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n248), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n811), .B1(new_n221), .B2(new_n547), .C1(new_n803), .C2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n827), .A2(G317), .B1(new_n887), .B2(G311), .ZN(new_n1133));
  XOR2_X1   g0933(.A(new_n1133), .B(KEYINPUT52), .Z(new_n1134));
  OAI21_X1  g0934(.A(new_n340), .B1(new_n824), .B2(new_n262), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n816), .A2(new_n823), .B1(new_n820), .B2(new_n833), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(G116), .C2(new_n837), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n828), .A2(G303), .B1(new_n896), .B2(G294), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n827), .A2(G150), .B1(new_n887), .B2(G159), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT51), .Z(new_n1141));
  OAI21_X1  g0941(.A(new_n256), .B1(new_n824), .B2(new_n654), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n816), .A2(new_n356), .B1(new_n820), .B2(new_n1006), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(G77), .C2(new_n837), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n828), .A2(G50), .B1(new_n896), .B2(new_n335), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1141), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1139), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n798), .B(new_n1132), .C1(new_n1147), .C2(new_n884), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n1038), .B2(new_n809), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n797), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT115), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1130), .A2(new_n1151), .A3(KEYINPUT115), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(G390));
  NAND3_X1  g0956(.A1(new_n978), .A2(G330), .A3(new_n981), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n868), .B1(new_n876), .B2(new_n706), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n930), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n928), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n967), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n966), .A2(new_n968), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n879), .B(new_n731), .C1(new_n787), .C2(new_n791), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n929), .B1(new_n1164), .B2(new_n930), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n947), .B1(new_n428), .B2(new_n937), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n965), .B1(new_n1166), .B2(KEYINPUT38), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1165), .A2(new_n1167), .A3(new_n967), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1158), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1160), .B1(new_n722), .B2(new_n869), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1162), .B1(new_n1170), .B2(new_n929), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n948), .A2(KEYINPUT39), .A3(new_n953), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT39), .B1(new_n953), .B2(new_n985), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1164), .A2(new_n930), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n986), .B(new_n1162), .C1(new_n1175), .C2(new_n929), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n776), .A2(new_n879), .A3(new_n928), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1169), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n537), .A2(G330), .A3(new_n981), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n975), .A2(new_n698), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1170), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n928), .B1(new_n776), .B2(new_n879), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT116), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1157), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(KEYINPUT116), .B(new_n928), .C1(new_n776), .C2(new_n879), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n981), .A2(G330), .A3(new_n879), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1175), .B(new_n1177), .C1(new_n928), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n753), .B1(new_n1179), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1169), .A2(new_n1190), .A3(new_n1178), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n807), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n798), .B1(new_n335), .B2(new_n885), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G107), .A2(new_n828), .B1(new_n827), .B2(G283), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n547), .B2(new_n832), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT118), .Z(new_n1199));
  OAI21_X1  g0999(.A(new_n340), .B1(new_n816), .B2(new_n654), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT119), .Z(new_n1201));
  OAI221_X1 g1001(.A(new_n901), .B1(new_n1109), .B2(new_n820), .C1(new_n459), .C2(new_n847), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G116), .B2(new_n887), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n827), .A2(G128), .B1(new_n887), .B2(G132), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT117), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n340), .B1(new_n821), .B2(G125), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT54), .B(G143), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1207), .B1(new_n485), .B2(new_n824), .C1(new_n832), .C2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G137), .B2(new_n828), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n817), .A2(G150), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1211), .A2(KEYINPUT53), .B1(G159), .B2(new_n837), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(KEYINPUT53), .C2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1204), .B1(new_n1206), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1196), .B1(new_n1214), .B2(new_n810), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1195), .A2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1179), .B2(new_n796), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1194), .A2(new_n1217), .ZN(G378));
  AND2_X1   g1018(.A1(new_n490), .A2(new_n730), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n498), .A2(new_n535), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n498), .B2(new_n535), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n978), .A2(KEYINPUT40), .A3(new_n981), .ZN(new_n1229));
  OAI21_X1  g1029(.A(G330), .B1(new_n1167), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n984), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n738), .B1(new_n986), .B2(new_n987), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n982), .B1(new_n948), .B2(new_n953), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1232), .B(new_n1233), .C1(KEYINPUT40), .C2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1231), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1236), .A2(new_n970), .A3(new_n973), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n958), .A2(new_n969), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1235), .B(new_n1231), .C1(new_n1238), .C2(new_n972), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(KEYINPUT121), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT121), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n974), .A2(new_n1241), .A3(new_n1235), .A4(new_n1231), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1240), .A2(new_n1242), .A3(new_n797), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n798), .B1(G50), .B2(new_n885), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n847), .A2(new_n482), .B1(new_n1208), .B2(new_n816), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n827), .A2(G125), .B1(new_n887), .B2(G128), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1010), .B2(new_n832), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(G132), .C2(new_n828), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT59), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n250), .B(new_n313), .C1(new_n824), .C2(new_n347), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G124), .B2(new_n821), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n827), .A2(G116), .B1(new_n896), .B2(new_n500), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n433), .B2(new_n889), .C1(new_n262), .C2(new_n834), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n816), .A2(new_n206), .B1(new_n820), .B2(new_n823), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n313), .B(new_n340), .C1(new_n824), .C2(new_n842), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1256), .A2(new_n1009), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT58), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1259), .A2(KEYINPUT58), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G50), .B1(new_n250), .B2(new_n313), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n256), .B2(G41), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1254), .A2(new_n1260), .A3(new_n1261), .A4(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1244), .B1(new_n1264), .B2(new_n810), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1228), .B2(new_n808), .ZN(new_n1266));
  XOR2_X1   g1066(.A(new_n1266), .B(KEYINPUT120), .Z(new_n1267));
  AND2_X1   g1067(.A1(new_n1243), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1181), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1193), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1240), .A2(new_n1242), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1237), .A2(KEYINPUT122), .A3(new_n1239), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT122), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n974), .A2(new_n1275), .A3(new_n1235), .A4(new_n1231), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1274), .A2(new_n1276), .A3(KEYINPUT57), .A4(new_n1270), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n752), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1268), .B1(new_n1273), .B2(new_n1278), .ZN(G375));
  NAND2_X1  g1079(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n796), .B(KEYINPUT123), .Z(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n929), .A2(new_n807), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n798), .B1(G68), .B2(new_n885), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(G159), .A2(new_n817), .B1(new_n821), .B2(G128), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n340), .B1(new_n900), .B2(G58), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n485), .C2(new_n847), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n827), .A2(G132), .B1(new_n896), .B2(G150), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n1288), .B1(new_n1010), .B2(new_n834), .C1(new_n889), .C2(new_n1208), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n828), .A2(G116), .B1(new_n896), .B2(G107), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1290), .B1(new_n823), .B2(new_n834), .C1(new_n1109), .C2(new_n1007), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G97), .A2(new_n817), .B1(new_n900), .B2(G77), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n256), .B1(new_n821), .B2(G303), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1106), .A3(new_n1293), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n1287), .A2(new_n1289), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1284), .B1(new_n1295), .B2(new_n810), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1280), .A2(new_n1282), .B1(new_n1283), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1190), .A2(new_n1082), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1181), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1298), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(G381));
  NOR2_X1   g1103(.A1(new_n1194), .A2(new_n1217), .ZN(new_n1304));
  INV_X1    g1104(.A(G390), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1302), .A4(new_n1306), .ZN(new_n1307));
  OR3_X1    g1107(.A1(G375), .A2(new_n1307), .A3(G387), .ZN(G407));
  INV_X1    g1108(.A(G343), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(G213), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(KEYINPUT124), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1304), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G407), .B(G213), .C1(G375), .C2(new_n1312), .ZN(G409));
  XNOR2_X1  g1113(.A(G393), .B(new_n859), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G390), .B(new_n1024), .C1(new_n1062), .C2(new_n1091), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1089), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1060), .A2(KEYINPUT114), .B1(new_n1084), .B2(new_n796), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(G390), .B1(new_n1321), .B2(new_n1024), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G387), .A2(new_n1305), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1323), .A2(new_n1324), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT126), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1327), .B(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1082), .B1(new_n1193), .B2(new_n1269), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1240), .A2(new_n1330), .A3(new_n1242), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT125), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT125), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1240), .A2(new_n1330), .A3(new_n1242), .A4(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1274), .A2(new_n1276), .A3(new_n1282), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1332), .A2(new_n1266), .A3(new_n1334), .A4(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1304), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G378), .B(new_n1268), .C1(new_n1273), .C2(new_n1278), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1310), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1300), .A2(KEYINPUT60), .A3(new_n1181), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n752), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1191), .A2(KEYINPUT60), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1342), .B1(new_n1343), .B2(new_n1301), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n912), .B1(new_n1344), .B2(new_n1298), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1343), .A2(new_n1301), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G384), .B(new_n1297), .C1(new_n1346), .C2(new_n1342), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1309), .A2(G213), .A3(G2897), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  AOI22_X1  g1150(.A1(new_n1345), .A2(new_n1347), .B1(G2897), .B2(new_n1311), .ZN(new_n1351));
  OR2_X1    g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1311), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT63), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1348), .A2(new_n1354), .ZN(new_n1355));
  AOI22_X1  g1155(.A1(new_n1340), .A2(new_n1352), .B1(new_n1353), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1348), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1339), .A2(new_n1357), .A3(new_n1310), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1354), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1329), .A2(new_n1356), .A3(new_n1359), .ZN(new_n1360));
  NOR2_X1   g1160(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1324), .B1(new_n1353), .B2(new_n1361), .ZN(new_n1362));
  XOR2_X1   g1162(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1363));
  NAND2_X1  g1163(.A1(new_n1358), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1353), .A2(KEYINPUT62), .A3(new_n1357), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1362), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1367));
  INV_X1    g1167(.A(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1360), .B1(new_n1366), .B2(new_n1368), .ZN(G405));
  NAND2_X1  g1169(.A1(G375), .A2(new_n1304), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1348), .B1(new_n1370), .B2(new_n1338), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1371), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1370), .A2(new_n1348), .A3(new_n1338), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1367), .ZN(G402));
endmodule


