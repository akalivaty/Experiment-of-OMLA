//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NOR2_X1   g0012(.A1(G58), .A2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G20), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  OR3_X1    g0017(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(KEYINPUT66), .B(G238), .Z(new_n223));
  AOI21_X1  g0023(.A(new_n222), .B1(G68), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(KEYINPUT67), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n227), .B(new_n228), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n220), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n244), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G179), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G226), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G87), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n259), .B(new_n260), .C1(new_n253), .C2(new_n254), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n255), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G45), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n205), .A2(G274), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n278), .C2(new_n270), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G232), .ZN(new_n283));
  AND4_X1   g0083(.A1(new_n252), .A2(new_n265), .A3(new_n277), .A4(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n275), .A2(new_n276), .B1(G232), .B2(new_n282), .ZN(new_n285));
  AOI21_X1  g0085(.A(G169), .B1(new_n285), .B2(new_n265), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT78), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT78), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(new_n252), .A3(new_n265), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n265), .A2(new_n277), .A3(new_n283), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT73), .A2(G58), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT8), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n205), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT77), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n217), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n298), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n294), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n304), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n278), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n312), .A2(new_n313), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT7), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n253), .A2(new_n254), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n206), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(G68), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(G58), .A2(G68), .ZN(new_n323));
  OAI21_X1  g0123(.A(G20), .B1(new_n323), .B2(new_n213), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n310), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n253), .A2(new_n254), .A3(G20), .ZN(new_n332));
  OAI21_X1  g0132(.A(G68), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n319), .A2(new_n216), .A3(new_n320), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n328), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n312), .A2(new_n206), .A3(new_n316), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n246), .B1(new_n337), .B2(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n319), .A2(new_n216), .A3(new_n320), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n327), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n309), .B1(new_n331), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT18), .B1(new_n292), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n331), .ZN(new_n346));
  INV_X1    g0146(.A(new_n309), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n348), .A2(new_n349), .A3(new_n287), .A4(new_n291), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n285), .A2(new_n351), .A3(new_n265), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n290), .B2(G200), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n346), .A2(new_n353), .A3(new_n347), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n353), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n345), .A2(new_n350), .A3(new_n356), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n282), .A2(G244), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n277), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n312), .A2(new_n316), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n362), .A3(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n258), .B1(new_n312), .B2(new_n316), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n362), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n223), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT70), .A2(G1698), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n361), .A2(new_n370), .A3(G232), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT74), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n371), .A2(new_n372), .B1(G107), .B2(new_n319), .ZN(new_n373));
  INV_X1    g0173(.A(new_n261), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT74), .A3(G232), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n367), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n360), .B1(new_n376), .B2(new_n264), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT75), .A3(new_n252), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n313), .A2(new_n315), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n278), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT8), .B(G58), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n206), .A2(new_n278), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n202), .A2(new_n216), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n304), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n305), .A2(G77), .A3(new_n295), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(G77), .C2(new_n301), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n377), .A2(G169), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT75), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n376), .A2(new_n264), .ZN(new_n394));
  INV_X1    g0194(.A(new_n360), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n392), .A2(new_n393), .B1(G179), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n396), .B2(G200), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n377), .A2(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n358), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n277), .B1(new_n221), .B2(new_n281), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n374), .A2(G222), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(KEYINPUT71), .B1(G77), .B2(new_n319), .ZN(new_n406));
  OAI21_X1  g0206(.A(G223), .B1(new_n364), .B2(new_n366), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n374), .A2(new_n408), .A3(G222), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n406), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n404), .B1(new_n410), .B2(new_n264), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n220), .B1(new_n205), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n305), .A2(new_n414), .B1(new_n220), .B2(new_n302), .ZN(new_n415));
  INV_X1    g0215(.A(G150), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n201), .A2(new_n206), .B1(new_n385), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n380), .B2(new_n294), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n418), .B2(new_n310), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT9), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n411), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT10), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n410), .A2(new_n264), .ZN(new_n424));
  INV_X1    g0224(.A(new_n404), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT10), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n412), .A4(new_n420), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n325), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n381), .B2(new_n202), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n304), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT11), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(KEYINPUT11), .A3(new_n304), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT12), .B1(new_n301), .B2(G68), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n246), .B1(new_n205), .B2(G20), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n437), .A2(new_n438), .B1(new_n305), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n275), .A2(new_n276), .B1(G238), .B2(new_n282), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n259), .A2(G226), .A3(new_n260), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G232), .A2(G1698), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n319), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G97), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n278), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n264), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n443), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n444), .B1(new_n443), .B2(new_n450), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n442), .B(G169), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n282), .A2(G238), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n277), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n450), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT13), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n443), .A2(new_n444), .A3(new_n450), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(G179), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n442), .B1(new_n461), .B2(G169), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n441), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(G200), .ZN(new_n464));
  INV_X1    g0264(.A(new_n441), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n351), .C2(new_n461), .ZN(new_n466));
  INV_X1    g0266(.A(new_n419), .ZN(new_n467));
  INV_X1    g0267(.A(G169), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n467), .B1(new_n426), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G179), .B2(new_n426), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n430), .A2(new_n463), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT79), .B1(new_n403), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n471), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n402), .A2(new_n358), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  INV_X1    g0278(.A(G257), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n312), .B2(new_n316), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(new_n370), .B1(new_n319), .B2(G303), .ZN(new_n481));
  OAI211_X1 g0281(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n279), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n266), .A2(G1), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(G270), .A3(new_n279), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n205), .A2(G45), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n485), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G274), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G169), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n278), .A2(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n313), .A2(new_n315), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT20), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n303), .A2(new_n217), .B1(G20), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(KEYINPUT85), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n302), .A2(new_n500), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n205), .A2(G33), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n310), .A2(G116), .A3(new_n301), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n499), .A2(KEYINPUT85), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n507), .B(new_n508), .C1(new_n498), .C2(new_n501), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n478), .B1(new_n495), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n494), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n312), .A2(G303), .A3(new_n316), .ZN(new_n513));
  OAI21_X1  g0313(.A(G257), .B1(new_n253), .B2(new_n254), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n259), .A2(new_n260), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n482), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n264), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n517), .A3(G190), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n494), .B1(new_n264), .B2(new_n516), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n510), .C1(new_n519), .C2(new_n421), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n468), .B1(new_n512), .B2(new_n517), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(KEYINPUT21), .B1(new_n519), .B2(G179), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n511), .B(new_n520), .C1(new_n522), .C2(new_n510), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT86), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n512), .A2(new_n517), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n495), .A2(new_n478), .B1(new_n252), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n510), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n529), .A2(KEYINPUT86), .A3(new_n511), .A4(new_n520), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n313), .B(new_n315), .C1(new_n253), .C2(new_n254), .ZN(new_n532));
  INV_X1    g0332(.A(G87), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(KEYINPUT87), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT22), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n361), .A2(new_n216), .A3(new_n537), .A4(new_n534), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n540), .A2(new_n541), .B1(new_n206), .B2(G107), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(G20), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n216), .A2(KEYINPUT23), .A3(G107), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n539), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n539), .B2(new_n546), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n304), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G13), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(G1), .ZN(new_n552));
  INV_X1    g0352(.A(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(G20), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT25), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n301), .A2(new_n504), .A3(new_n217), .A4(new_n303), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(G107), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT89), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n488), .A2(G264), .A3(new_n279), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n493), .ZN(new_n562));
  OAI211_X1 g0362(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G294), .ZN(new_n564));
  INV_X1    g0364(.A(G250), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n261), .C2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n562), .B1(new_n264), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n560), .B1(new_n567), .B2(new_n468), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT90), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n488), .A2(new_n570), .A3(G264), .A4(new_n279), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n569), .A2(new_n571), .B1(new_n566), .B2(new_n264), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G179), .A3(new_n493), .ZN(new_n573));
  INV_X1    g0373(.A(new_n562), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n566), .A2(new_n264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(KEYINPUT89), .A3(G169), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n568), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n559), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n576), .A2(G190), .ZN(new_n580));
  AOI21_X1  g0380(.A(G200), .B1(new_n572), .B2(new_n493), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n550), .B(new_n558), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  OR3_X1    g0383(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n533), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT84), .B1(new_n556), .B2(new_n533), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n313), .A2(new_n315), .A3(G33), .A4(G97), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n361), .A2(new_n216), .A3(G68), .ZN(new_n590));
  NAND3_X1  g0390(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n313), .A2(new_n315), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n533), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n304), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n382), .A2(new_n302), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n586), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n600));
  INV_X1    g0400(.A(G238), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n543), .B(new_n600), .C1(new_n261), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n264), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n272), .A2(G45), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n490), .A2(G250), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n264), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n421), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n351), .B(new_n606), .C1(new_n602), .C2(new_n264), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n599), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n603), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G169), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n603), .A2(G179), .A3(new_n607), .ZN(new_n613));
  INV_X1    g0413(.A(new_n382), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n557), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n597), .A2(new_n598), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n612), .A2(new_n613), .B1(new_n616), .B2(KEYINPUT83), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n302), .A2(new_n448), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n556), .B2(new_n448), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n318), .A2(G107), .A3(new_n321), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n385), .A2(new_n202), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT6), .ZN(new_n624));
  AND2_X1   g0424(.A1(G97), .A2(G107), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n593), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n553), .A2(KEYINPUT6), .A3(G97), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n623), .B1(new_n628), .B2(new_n379), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n621), .B1(new_n630), .B2(new_n304), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n365), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n632));
  OAI21_X1  g0432(.A(G244), .B1(new_n253), .B2(new_n254), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n260), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT80), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT4), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n368), .A2(new_n369), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G244), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n312), .B2(new_n316), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT80), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n633), .B2(new_n515), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n632), .A2(new_n635), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n264), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n488), .A2(new_n279), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n493), .B1(new_n645), .B2(new_n479), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n631), .B1(new_n648), .B2(new_n468), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n646), .B1(new_n643), .B2(new_n264), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT82), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n650), .A2(new_n651), .A3(new_n252), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n650), .B2(new_n252), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n644), .A2(G190), .A3(new_n647), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT81), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n648), .A2(G200), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT81), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n650), .A2(new_n658), .A3(G190), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n656), .A2(new_n657), .A3(new_n631), .A4(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n619), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n477), .A2(new_n531), .A3(new_n583), .A4(new_n661), .ZN(G372));
  INV_X1    g0462(.A(new_n470), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n345), .A2(new_n350), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n398), .A2(new_n463), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n466), .A2(new_n356), .A3(new_n357), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n663), .B1(new_n668), .B2(new_n430), .ZN(new_n669));
  INV_X1    g0469(.A(new_n477), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n310), .B1(new_n622), .B2(new_n629), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n650), .A2(G169), .B1(new_n671), .B2(new_n621), .ZN(new_n672));
  OAI21_X1  g0472(.A(KEYINPUT82), .B1(new_n648), .B2(G179), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n650), .A2(new_n651), .A3(new_n252), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n619), .A2(new_n675), .A3(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n610), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n612), .A2(new_n613), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n616), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n654), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n676), .B1(new_n681), .B2(KEYINPUT26), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n582), .A2(new_n677), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT21), .B1(new_n528), .B2(new_n521), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n527), .B2(new_n528), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n579), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(new_n686), .A3(new_n654), .A4(new_n660), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n687), .A3(new_n679), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n669), .B1(new_n670), .B2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(new_n685), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n216), .A2(new_n552), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n528), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT91), .ZN(new_n699));
  MUX2_X1   g0499(.A(new_n531), .B(new_n691), .S(new_n699), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n559), .A2(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n583), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n559), .A2(new_n578), .A3(new_n697), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n700), .A2(G330), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n697), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n579), .A2(new_n582), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n691), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n559), .A2(new_n578), .A3(new_n706), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(KEYINPUT92), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT92), .B1(new_n708), .B2(new_n709), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n705), .B1(new_n711), .B2(new_n712), .ZN(G399));
  NOR2_X1   g0513(.A1(new_n594), .A2(G116), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G1), .ZN(new_n715));
  INV_X1    g0515(.A(new_n209), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n716), .A2(KEYINPUT93), .A3(G41), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT93), .B1(new_n716), .B2(G41), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g0519(.A(new_n215), .B(new_n715), .S(new_n719), .Z(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  AOI21_X1  g0521(.A(KEYINPUT26), .B1(new_n619), .B2(new_n675), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n681), .A2(KEYINPUT26), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n687), .A2(new_n679), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n706), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n688), .A2(new_n706), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n252), .B(new_n606), .C1(new_n602), .C2(new_n264), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n650), .A2(new_n519), .A3(new_n572), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n569), .A2(new_n571), .ZN(new_n738));
  AND4_X1   g0538(.A1(new_n517), .A2(new_n738), .A3(new_n512), .A4(new_n575), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .A3(new_n650), .A4(new_n734), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n572), .A2(new_n493), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n512), .B2(new_n517), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n648), .A2(new_n741), .A3(new_n611), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n737), .A2(new_n740), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT31), .B1(new_n744), .B2(new_n697), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n661), .A2(new_n531), .A3(new_n707), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n721), .B1(new_n752), .B2(G1), .ZN(G364));
  INV_X1    g0553(.A(new_n719), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n379), .A2(new_n551), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G45), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G1), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n700), .B2(G330), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n700), .ZN(new_n760));
  INV_X1    g0560(.A(new_n758), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n250), .A2(new_n266), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n716), .A2(new_n361), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n215), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n267), .A2(new_n269), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n762), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n209), .A2(new_n361), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n209), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n767), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n768), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n217), .B1(G20), .B2(new_n468), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n761), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  NOR4_X1   g0579(.A1(new_n216), .A2(G179), .A3(G190), .A4(new_n421), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT96), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G107), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n206), .A2(new_n351), .A3(new_n421), .A4(G179), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n319), .B1(new_n783), .B2(G87), .ZN(new_n784));
  INV_X1    g0584(.A(G58), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n216), .A2(new_n252), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n351), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n786), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n790), .A2(new_n351), .A3(new_n421), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n790), .A2(G190), .A3(new_n421), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n220), .A2(new_n792), .B1(new_n794), .B2(new_n246), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n216), .B1(new_n252), .B2(new_n787), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n448), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G190), .A2(G200), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n379), .A2(new_n252), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  OR3_X1    g0604(.A1(new_n803), .A2(KEYINPUT32), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(KEYINPUT32), .B1(new_n803), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n786), .A2(new_n802), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n805), .B(new_n806), .C1(new_n202), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n807), .A2(new_n810), .B1(new_n797), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G329), .ZN(new_n813));
  INV_X1    g0613(.A(new_n783), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n319), .B1(new_n803), .B2(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n788), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n812), .B(new_n816), .C1(G322), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT33), .B(G317), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n793), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT98), .B(G326), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n792), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G283), .C2(new_n781), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n796), .A2(new_n809), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n777), .ZN(new_n825));
  INV_X1    g0625(.A(new_n776), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n779), .B1(new_n824), .B2(new_n825), .C1(new_n700), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n760), .A2(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n389), .A2(new_n697), .ZN(new_n829));
  AOI211_X1 g0629(.A(G179), .B(new_n360), .C1(new_n376), .C2(new_n264), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n396), .A2(new_n468), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n830), .B1(new_n831), .B2(KEYINPUT75), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n401), .B(new_n829), .C1(new_n832), .C2(new_n390), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n397), .A2(new_n378), .A3(new_n389), .A4(new_n697), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n730), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n688), .A2(new_n706), .A3(new_n835), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n758), .B1(new_n839), .B2(new_n750), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n750), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n777), .A2(new_n774), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n758), .B1(G77), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n319), .B1(new_n814), .B2(new_n553), .ZN(new_n845));
  INV_X1    g0645(.A(new_n803), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(G311), .B2(new_n846), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n500), .B2(new_n807), .C1(new_n811), .C2(new_n788), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n801), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n781), .A2(G87), .B1(G303), .B2(new_n791), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT99), .B(G283), .Z(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n850), .C1(new_n794), .C2(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G137), .A2(new_n791), .B1(new_n793), .B2(G150), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT100), .Z(new_n854));
  INV_X1    g0654(.A(new_n807), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n817), .B1(new_n855), .B2(G159), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n781), .A2(G68), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n361), .B1(new_n814), .B2(new_n220), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G132), .B2(new_n846), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n859), .B(new_n861), .C1(new_n785), .C2(new_n797), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n844), .B1(new_n863), .B2(new_n777), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n775), .B2(new_n835), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n841), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  NOR3_X1   g0667(.A1(new_n216), .A2(new_n500), .A3(new_n217), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n628), .B(KEYINPUT101), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g0673(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n873), .B(new_n874), .ZN(new_n875));
  OR3_X1    g0675(.A1(new_n215), .A2(new_n202), .A3(new_n323), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n205), .B(G13), .C1(new_n876), .C2(new_n245), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n391), .A2(new_n397), .A3(new_n706), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n838), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n838), .A2(KEYINPUT103), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT104), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n310), .B1(new_n886), .B2(new_n330), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n885), .A2(new_n887), .B1(new_n336), .B2(new_n342), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n304), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n309), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n354), .B1(new_n891), .B2(new_n292), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n695), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n348), .A2(new_n287), .A3(new_n291), .ZN(new_n895));
  INV_X1    g0695(.A(new_n695), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n348), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n895), .A2(new_n897), .A3(new_n898), .A4(new_n354), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n894), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n358), .A2(new_n893), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n894), .A2(new_n899), .B1(new_n358), .B2(new_n893), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n465), .A2(new_n706), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n463), .A2(new_n466), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n463), .B2(new_n466), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n884), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n354), .B1(new_n292), .B2(new_n344), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n344), .A2(new_n695), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n899), .A2(new_n918), .B1(new_n358), .B2(new_n917), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n915), .B1(new_n919), .B2(KEYINPUT38), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n899), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n358), .A2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(KEYINPUT106), .A3(new_n903), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n924), .A3(new_n906), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n463), .A2(new_n697), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT105), .Z(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n900), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n665), .A2(new_n896), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n914), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n477), .A2(new_n732), .A3(new_n729), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n669), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(G330), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT107), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n661), .A2(new_n531), .A3(new_n707), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n744), .A2(new_n697), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT31), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n943), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n463), .A2(new_n466), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n908), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n463), .A2(new_n466), .A3(new_n909), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n833), .B2(new_n834), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT107), .ZN(new_n955));
  AND4_X1   g0755(.A1(KEYINPUT40), .A2(new_n950), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n925), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n950), .A2(new_n954), .A3(new_n955), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n933), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT107), .B1(new_n747), .B2(new_n748), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT107), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n670), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n942), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n941), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n205), .B2(new_n755), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n941), .A2(new_n966), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n878), .B1(new_n968), .B2(new_n969), .ZN(G367));
  XNOR2_X1  g0770(.A(new_n719), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n704), .B1(new_n691), .B2(new_n706), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n691), .B2(new_n707), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n700), .A2(G330), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n752), .ZN(new_n977));
  INV_X1    g0777(.A(new_n712), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n654), .B(new_n660), .C1(new_n631), .C2(new_n706), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n675), .A2(new_n697), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n978), .A2(new_n710), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n984));
  INV_X1    g0784(.A(new_n705), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n984), .B1(KEYINPUT110), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n982), .B1(new_n978), .B2(new_n710), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n983), .A2(KEYINPUT44), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n985), .A2(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n991), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n986), .A2(new_n988), .A3(new_n993), .A4(new_n989), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n977), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n752), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n972), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n757), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n982), .A2(new_n708), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(KEYINPUT42), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n654), .B1(new_n979), .B2(new_n579), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1002), .A2(new_n1003), .B1(new_n706), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n599), .A2(new_n697), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n679), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n677), .A2(new_n679), .A3(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  MUX2_X1   g0810(.A(new_n1006), .B(KEYINPUT43), .S(new_n1010), .Z(new_n1011));
  OR2_X1    g0811(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1005), .A2(new_n1009), .A3(new_n1008), .A4(new_n1006), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT109), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(KEYINPUT109), .A3(new_n1013), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1015), .A2(new_n985), .A3(new_n981), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1016), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1018), .A2(new_n1014), .B1(new_n705), .B2(new_n982), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1000), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n814), .B2(new_n500), .ZN(new_n1023));
  INV_X1    g0823(.A(G317), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n780), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n803), .C1(new_n1025), .C2(new_n448), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G311), .B2(new_n791), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n815), .A2(new_n788), .B1(new_n807), .B2(new_n851), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n319), .C1(new_n553), .C2(new_n797), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1027), .B(new_n1031), .C1(new_n811), .C2(new_n794), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n361), .B1(new_n785), .B2(new_n814), .C1(new_n1025), .C2(new_n202), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G137), .B2(new_n846), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n800), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(G68), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G50), .A2(new_n855), .B1(new_n817), .B2(G150), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G143), .A2(new_n791), .B1(new_n793), .B2(G159), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1032), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n777), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n763), .A2(new_n240), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n778), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n716), .B2(new_n614), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n761), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1042), .B(new_n1046), .C1(new_n826), .C2(new_n1010), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1021), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(G387));
  OR2_X1    g0850(.A1(new_n976), .A2(new_n752), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(new_n754), .A3(new_n977), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n702), .A2(new_n703), .A3(new_n776), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n763), .B1(new_n237), .B2(new_n766), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n714), .B2(new_n769), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n384), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1057), .A2(new_n714), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1055), .A2(new_n1059), .B1(new_n553), .B2(new_n716), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n758), .B1(new_n1060), .B2(new_n1044), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n361), .B1(new_n788), .B2(new_n220), .C1(new_n246), .C2(new_n807), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n794), .A2(new_n307), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G97), .C2(new_n781), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n791), .A2(G159), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n783), .A2(G77), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n416), .B2(new_n803), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT111), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n1035), .A2(new_n614), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1064), .A2(new_n1066), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT113), .Z(new_n1072));
  AOI21_X1  g0872(.A(new_n361), .B1(new_n780), .B2(G116), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n797), .A2(new_n851), .B1(new_n814), .B2(new_n811), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G303), .A2(new_n855), .B1(new_n817), .B2(G317), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n791), .A2(G322), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(new_n810), .C2(new_n794), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1073), .B1(new_n803), .B2(new_n821), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1061), .B1(new_n1084), .B2(new_n777), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n976), .A2(new_n757), .B1(new_n1053), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1052), .A2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n992), .A2(new_n994), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n757), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n778), .B1(new_n448), .B2(new_n209), .C1(new_n764), .C2(new_n244), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n758), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n781), .A2(G87), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n361), .B1(new_n814), .B2(new_n246), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G143), .B2(new_n846), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(new_n384), .C2(new_n807), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G50), .B2(new_n793), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n791), .A2(G150), .B1(G159), .B2(new_n817), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n1035), .A2(G77), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n319), .B1(new_n814), .B2(new_n851), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G322), .B2(new_n846), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n782), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT115), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n797), .A2(new_n500), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n793), .B2(G303), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1104), .B1(KEYINPUT116), .B2(new_n1107), .C1(new_n811), .C2(new_n807), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n792), .A2(new_n1024), .B1(new_n788), .B2(new_n810), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1109), .A2(new_n1111), .B1(new_n1107), .B2(KEYINPUT116), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1100), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1091), .B1(new_n1114), .B2(new_n777), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n826), .B2(new_n981), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n995), .A2(new_n719), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1088), .B1(new_n752), .B2(new_n976), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1089), .B(new_n1116), .C1(new_n1117), .C2(new_n1118), .ZN(G390));
  OAI211_X1 g0919(.A(new_n706), .B(new_n835), .C1(new_n727), .C2(new_n728), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n913), .A2(new_n749), .A3(G330), .A4(new_n835), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n879), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n950), .A2(G330), .A3(new_n955), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n912), .B1(new_n1123), .B2(new_n836), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n912), .B1(new_n750), .B2(new_n836), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n950), .A2(new_n954), .A3(G330), .A4(new_n955), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1122), .A2(new_n1124), .B1(new_n884), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n477), .A2(G330), .A3(new_n950), .A4(new_n955), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n939), .A3(new_n669), .ZN(new_n1130));
  OAI21_X1  g0930(.A(KEYINPUT117), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n884), .A2(new_n1127), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n879), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n726), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n724), .A3(new_n723), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n728), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n697), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1133), .B1(new_n1137), .B2(new_n835), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1124), .A2(new_n1138), .A3(new_n1121), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1129), .A2(new_n939), .A3(new_n669), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1131), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n912), .B1(new_n882), .B2(new_n883), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT38), .B1(new_n921), .B2(new_n922), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(KEYINPUT106), .B1(KEYINPUT38), .B2(new_n905), .ZN(new_n1147));
  AOI21_X1  g0947(.A(KEYINPUT39), .B1(new_n1147), .B2(new_n920), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n907), .A2(new_n926), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1145), .A2(new_n930), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n930), .B1(new_n1147), .B2(new_n920), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n912), .B2(new_n1138), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1152), .A3(new_n1121), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n883), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT103), .B1(new_n838), .B2(new_n879), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n913), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n929), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n927), .A2(new_n934), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1138), .A2(new_n912), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1157), .A2(new_n1158), .B1(new_n1159), .B2(new_n1151), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1153), .B1(new_n1160), .B2(new_n1126), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n719), .B1(new_n1144), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1150), .A2(new_n1152), .A3(new_n1121), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1126), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1131), .A2(new_n1143), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1162), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n757), .B(new_n1153), .C1(new_n1160), .C2(new_n1126), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1158), .A2(new_n774), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n758), .B1(new_n294), .B2(new_n843), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n416), .ZN(new_n1172));
  OAI21_X1  g0972(.A(KEYINPUT53), .B1(new_n814), .B2(new_n416), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1025), .B2(new_n220), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G128), .C2(new_n791), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n793), .A2(G137), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n800), .A2(new_n804), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n319), .B1(new_n846), .B2(G125), .ZN(new_n1179));
  INV_X1    g0979(.A(G132), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1179), .B1(new_n788), .B2(new_n1180), .C1(new_n1182), .C2(new_n807), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1177), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n791), .A2(G283), .B1(G97), .B2(new_n855), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n553), .B2(new_n794), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT119), .Z(new_n1187));
  AOI21_X1  g0987(.A(new_n361), .B1(new_n783), .B2(G87), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT120), .Z(new_n1189));
  AOI22_X1  g0989(.A1(new_n817), .A2(G116), .B1(G294), .B2(new_n846), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n859), .A2(new_n1099), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1184), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1171), .B1(new_n1192), .B2(new_n777), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1170), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1169), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1168), .A2(new_n1196), .ZN(G378));
  XNOR2_X1  g0997(.A(new_n1130), .B(KEYINPUT124), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n430), .A2(new_n470), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n467), .A2(new_n695), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n835), .B1(new_n910), .B2(new_n911), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n963), .A2(new_n962), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n907), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n942), .B1(new_n1212), .B2(new_n958), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1209), .B1(new_n1213), .B2(new_n957), .ZN(new_n1214));
  AND4_X1   g1014(.A1(G330), .A2(new_n957), .A3(new_n960), .A4(new_n1209), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n938), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n957), .A2(new_n960), .A3(G330), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1209), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n936), .B1(new_n1145), .B2(new_n907), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n957), .A2(new_n960), .A3(new_n1209), .A4(G330), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1219), .A2(new_n935), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1216), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT57), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n754), .B1(new_n1199), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT57), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT123), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1216), .A2(new_n1222), .A3(KEYINPUT123), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1231), .B2(new_n1199), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n758), .B1(G50), .B2(new_n843), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n780), .A2(G58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n846), .A2(G283), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n361), .A2(G41), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n1067), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G107), .A2(new_n817), .B1(new_n855), .B2(new_n614), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G97), .A2(new_n793), .B1(new_n791), .B2(G116), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1036), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT121), .ZN(new_n1242));
  INV_X1    g1042(.A(G128), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1182), .A2(new_n814), .B1(new_n788), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G137), .B2(new_n855), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G125), .A2(new_n791), .B1(new_n793), .B2(G132), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n416), .C2(new_n800), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n780), .A2(G159), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G33), .B(G41), .C1(new_n846), .C2(G124), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(KEYINPUT58), .A2(new_n1242), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1253), .B1(KEYINPUT58), .B2(new_n1242), .C1(new_n1237), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n777), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT122), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1234), .B(new_n1257), .C1(new_n774), .C2(new_n1218), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1216), .A2(KEYINPUT123), .A3(new_n1222), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1228), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1260), .B2(new_n757), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1233), .A2(new_n1261), .ZN(G375));
  OAI21_X1  g1062(.A(new_n758), .B1(G68), .B2(new_n843), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G137), .A2(new_n817), .B1(new_n855), .B2(G150), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n846), .A2(G128), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n319), .B1(new_n783), .B2(G159), .ZN(new_n1266));
  AND4_X1   g1066(.A1(new_n1235), .A2(new_n1264), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n1180), .B2(new_n792), .C1(new_n794), .C2(new_n1182), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n800), .A2(new_n220), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n781), .A2(G77), .B1(G294), .B2(new_n791), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n500), .B2(new_n794), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n319), .B1(new_n814), .B2(new_n448), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G303), .B2(new_n846), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n817), .A2(G283), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n855), .A2(G107), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1070), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n1268), .A2(new_n1269), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1263), .B1(new_n1277), .B2(new_n777), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n775), .B2(new_n913), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n1128), .B2(new_n998), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1131), .A2(new_n1143), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n971), .ZN(G381));
  NAND4_X1  g1084(.A1(new_n1052), .A2(new_n827), .A3(new_n760), .A4(new_n1086), .ZN(new_n1285));
  OR3_X1    g1085(.A1(G390), .A2(G384), .A3(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(G387), .A2(G381), .A3(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(G375), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1195), .B1(new_n1162), .B2(new_n1167), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1288), .A3(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G213), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(G343), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1288), .A2(new_n1289), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1293), .B(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1096(.A(new_n1198), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1144), .B2(new_n1161), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT57), .B1(new_n1260), .B2(new_n1298), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1261), .C1(new_n1299), .C2(new_n1225), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n972), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1258), .B1(new_n1223), .B2(new_n757), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1289), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1292), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1283), .A2(KEYINPUT60), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n719), .B1(new_n1282), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1311), .B2(new_n1281), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n866), .B(new_n1280), .C1(new_n1308), .C2(new_n1310), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1292), .A2(G2897), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G2897), .B(new_n1292), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1314), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1320), .B1(new_n1307), .B2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G390), .B(new_n1047), .C1(new_n1000), .C2(new_n1020), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G393), .A2(G396), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1285), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(KEYINPUT126), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1324), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(G390), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1021), .B2(new_n1048), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1323), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1330), .A2(new_n1323), .A3(new_n1327), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1292), .B1(new_n1300), .B2(new_n1304), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(KEYINPUT63), .A3(new_n1314), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1319), .A2(new_n1322), .A3(new_n1335), .A4(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1336), .A2(new_n1339), .A3(new_n1314), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1341), .B1(new_n1336), .B2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1339), .B1(new_n1336), .B2(new_n1314), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1340), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1338), .B1(new_n1345), .B2(new_n1335), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1289), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1321), .A3(new_n1300), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G378), .B1(new_n1233), .B2(new_n1261), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1300), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1314), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1348), .A2(new_n1351), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1352), .A2(new_n1335), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1335), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


