//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT92), .ZN(new_n203));
  INV_X1    g002(.A(G227gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT66), .B1(new_n208), .B2(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n208), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217));
  INV_X1    g016(.A(new_n215), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n212), .A2(new_n213), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT24), .B1(new_n209), .B2(new_n210), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n216), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n228));
  AND2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n215), .B1(new_n229), .B2(KEYINPUT24), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n229), .B2(KEYINPUT24), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n232), .A3(new_n208), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT25), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT65), .A4(new_n233), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n222), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n240), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT70), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n241), .A2(new_n224), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(G183gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n245), .B(G190gat), .C1(new_n248), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n251), .A2(new_n253), .ZN(new_n256));
  INV_X1    g055(.A(G190gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT28), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n213), .B(new_n244), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n228), .A2(new_n238), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G120gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  OR3_X1    g064(.A1(new_n265), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n264), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(KEYINPUT1), .B2(new_n261), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n259), .A2(new_n238), .ZN(new_n272));
  INV_X1    g071(.A(new_n270), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n228), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n207), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT32), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT34), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n271), .A2(new_n274), .A3(new_n207), .ZN(new_n278));
  XNOR2_X1  g077(.A(G15gat), .B(G43gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  OAI211_X1 g080(.A(new_n278), .B(new_n281), .C1(new_n275), .C2(KEYINPUT33), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n260), .A2(new_n270), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n273), .B1(new_n272), .B2(new_n228), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  INV_X1    g085(.A(new_n281), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n207), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n206), .B1(new_n283), .B2(new_n284), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT34), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(KEYINPUT32), .A3(new_n290), .ZN(new_n291));
  AND4_X1   g090(.A1(new_n277), .A2(new_n282), .A3(new_n288), .A4(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n288), .A2(new_n282), .B1(new_n291), .B2(new_n277), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT31), .B(G50gat), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT85), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G78gat), .ZN(new_n297));
  INV_X1    g096(.A(G106gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300));
  INV_X1    g099(.A(G155gat), .ZN(new_n301));
  INV_X1    g100(.A(G162gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n302), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT81), .ZN(new_n309));
  XOR2_X1   g108(.A(G141gat), .B(G148gat), .Z(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT82), .B(KEYINPUT2), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n306), .B1(new_n303), .B2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n302), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n307), .B1(new_n317), .B2(KEYINPUT2), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n310), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G218gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT22), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  AND2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G197gat), .A2(G204gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n323), .B(new_n325), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G218gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G197gat), .B(G204gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(new_n328), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n321), .B(new_n330), .C1(new_n334), .C2(new_n329), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n333), .B2(new_n328), .ZN(new_n336));
  INV_X1    g135(.A(new_n330), .ZN(new_n337));
  OAI21_X1  g136(.A(G218gat), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT29), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n320), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n335), .A2(new_n338), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n344), .A3(new_n319), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n340), .A2(new_n342), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n346), .B1(new_n335), .B2(new_n338), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n320), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n348), .A3(KEYINPUT86), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n350), .B1(new_n341), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n299), .B1(new_n357), .B2(KEYINPUT87), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n341), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n350), .ZN(new_n361));
  AND4_X1   g160(.A1(KEYINPUT87), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n357), .B2(KEYINPUT87), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(KEYINPUT87), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G22gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n359), .A2(new_n361), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT87), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n357), .A2(KEYINPUT87), .A3(new_n360), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n299), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n294), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n346), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n227), .A2(KEYINPUT25), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n259), .A2(new_n238), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n228), .A2(KEYINPUT75), .A3(new_n238), .A4(new_n259), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n376), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n343), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n260), .A2(new_n373), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n374), .A3(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n260), .A2(new_n387), .A3(new_n373), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n343), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(new_n384), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n380), .A2(new_n381), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n343), .B(new_n397), .C1(new_n398), .C2(new_n376), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n399), .A3(new_n394), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n395), .B1(KEYINPUT30), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n390), .B2(new_n394), .ZN(new_n406));
  NOR4_X1   g205(.A1(new_n385), .A2(new_n389), .A3(KEYINPUT77), .A4(new_n393), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n404), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n400), .A2(KEYINPUT77), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n396), .A2(new_n399), .A3(new_n405), .A4(new_n394), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n404), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n372), .A2(new_n402), .A3(new_n409), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT91), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n316), .A2(new_n319), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT84), .B1(new_n418), .B2(new_n273), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT84), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n320), .A2(new_n420), .A3(new_n270), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n418), .A2(KEYINPUT4), .A3(new_n273), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n270), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n345), .A3(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(new_n423), .A3(new_n424), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n320), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n419), .B2(new_n421), .ZN(new_n431));
  INV_X1    g230(.A(new_n423), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n433), .A3(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n273), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n420), .ZN(new_n436));
  INV_X1    g235(.A(new_n421), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n417), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n432), .A2(KEYINPUT5), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n438), .A2(new_n428), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(G85gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT0), .B(G57gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  INV_X1    g247(.A(new_n446), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n416), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n203), .B1(new_n415), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n364), .A2(new_n371), .ZN(new_n459));
  INV_X1    g258(.A(new_n294), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT92), .B1(new_n202), .B2(KEYINPUT91), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n413), .B1(new_n412), .B2(new_n404), .ZN(new_n463));
  AOI211_X1 g262(.A(KEYINPUT79), .B(new_n403), .C1(new_n410), .C2(new_n411), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n451), .A2(new_n452), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n462), .A2(new_n465), .A3(new_n402), .A4(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n455), .A2(new_n458), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n409), .A2(new_n402), .A3(new_n414), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n438), .A2(new_n428), .A3(new_n439), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n432), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n449), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n475), .A3(new_n449), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n470), .A2(new_n432), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n478), .B(KEYINPUT39), .C1(new_n432), .C2(new_n431), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT40), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n472), .A2(new_n475), .A3(new_n449), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n475), .B1(new_n472), .B2(new_n449), .ZN(new_n482));
  OAI211_X1 g281(.A(KEYINPUT40), .B(new_n479), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n447), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n459), .ZN(new_n487));
  INV_X1    g286(.A(new_n466), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n394), .B1(new_n390), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n489), .B2(new_n390), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT38), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n386), .A2(new_n388), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n383), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n386), .A2(KEYINPUT90), .A3(new_n343), .A4(new_n388), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT38), .B1(new_n498), .B2(KEYINPUT37), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n490), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n488), .A2(new_n492), .A3(new_n412), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n487), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n409), .A2(new_n402), .A3(new_n414), .A4(new_n466), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n459), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n294), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n510), .C1(new_n292), .C2(new_n293), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n503), .B2(new_n459), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n505), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n468), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G99gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT101), .B1(new_n521), .B2(new_n298), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT101), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(G99gat), .A3(G106gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(KEYINPUT8), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT102), .B(G85gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n525), .B(new_n527), .C1(G92gat), .C2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G99gat), .B(G106gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT103), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G57gat), .B(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G71gat), .B(G78gat), .Z(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT98), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT107), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n529), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(new_n530), .Z(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT10), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n535), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n540), .B(KEYINPUT98), .Z(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT10), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n520), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n519), .B1(new_n542), .B2(new_n546), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT108), .ZN(new_n555));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(KEYINPUT108), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OR3_X1    g362(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n564), .A2(new_n565), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  INV_X1    g365(.A(G50gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(G43gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(G43gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(KEYINPUT15), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT93), .B(G43gat), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(new_n572), .B2(new_n567), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n566), .B(new_n571), .C1(new_n573), .C2(KEYINPUT15), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n575), .B(new_n576), .C1(new_n566), .C2(new_n571), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT16), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n579), .B2(G1gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(G1gat), .B2(new_n578), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G8gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n583), .A2(KEYINPUT95), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(KEYINPUT95), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT13), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n577), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n582), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n588), .A3(new_n585), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n598), .A2(KEYINPUT18), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(KEYINPUT18), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n591), .A2(new_n592), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  INV_X1    g401(.A(G197gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT11), .B(G169gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT12), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  OAI221_X1 g408(.A(new_n609), .B1(new_n599), .B2(new_n600), .C1(new_n591), .C2(new_n592), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT97), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n601), .A2(new_n612), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n518), .A2(new_n563), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n582), .B1(new_n550), .B2(KEYINPUT21), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G183gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n550), .A2(KEYINPUT21), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT99), .B(G211gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n620), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G127gat), .B(G155gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n624), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n594), .A2(new_n535), .A3(new_n596), .ZN(new_n630));
  AND2_X1   g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n549), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n634), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n637), .A2(KEYINPUT106), .A3(new_n640), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT100), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n644), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n616), .A2(new_n629), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n466), .B(KEYINPUT109), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  INV_X1    g457(.A(new_n469), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT16), .B(G8gat), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n653), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n662));
  OAI21_X1  g461(.A(G8gat), .B1(new_n653), .B2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n653), .A2(new_n666), .A3(new_n513), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n654), .A2(new_n294), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n487), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(new_n629), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n650), .A2(new_n651), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n616), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(G29gat), .A3(new_n655), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n676), .B(KEYINPUT45), .Z(new_n677));
  NAND2_X1  g476(.A1(new_n502), .A2(new_n516), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n468), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n674), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n652), .A2(new_n681), .ZN(new_n682));
  AOI22_X1  g481(.A1(new_n680), .A2(new_n681), .B1(new_n518), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n562), .B(KEYINPUT110), .Z(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n614), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n673), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n683), .A2(KEYINPUT111), .A3(new_n673), .A4(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G29gat), .B1(new_n691), .B2(new_n655), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n692), .ZN(G1328gat));
  OAI21_X1  g492(.A(G36gat), .B1(new_n691), .B2(new_n659), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n675), .A2(G36gat), .A3(new_n659), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(G1329gat));
  NOR3_X1   g496(.A1(new_n675), .A2(new_n572), .A3(new_n460), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n572), .B1(new_n686), .B2(new_n513), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n690), .A2(new_n512), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n698), .B1(new_n702), .B2(new_n572), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n703), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g503(.A(KEYINPUT48), .B(G50gat), .C1(new_n686), .C2(new_n487), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n459), .A2(new_n567), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT112), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n675), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT113), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n705), .B(new_n708), .C1(new_n709), .C2(KEYINPUT48), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n690), .A2(new_n459), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(G50gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g513(.A1(new_n465), .A2(new_n372), .A3(new_n402), .A4(new_n453), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n457), .B1(new_n715), .B2(new_n203), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n716), .A2(new_n467), .B1(new_n502), .B2(new_n516), .ZN(new_n717));
  INV_X1    g516(.A(new_n684), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n629), .A2(new_n652), .A3(new_n614), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n655), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT114), .B(G57gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1332gat));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n659), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT49), .B(G64gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n726), .B2(new_n729), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n722), .B2(new_n513), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n719), .A2(new_n294), .A3(new_n721), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(G71gat), .B2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g533(.A1(new_n722), .A2(new_n487), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g535(.A1(new_n615), .A2(new_n629), .A3(new_n563), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT115), .B1(new_n683), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n518), .A2(new_n682), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n681), .B1(new_n717), .B2(new_n652), .ZN(new_n740));
  AND4_X1   g539(.A1(KEYINPUT115), .A2(new_n739), .A3(new_n740), .A4(new_n737), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n528), .B1(new_n742), .B2(new_n655), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n717), .A2(new_n652), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n615), .A2(new_n629), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n562), .A3(new_n749), .ZN(new_n750));
  OR2_X1    g549(.A1(new_n655), .A2(new_n528), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n743), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NOR2_X1   g551(.A1(new_n718), .A2(new_n659), .ZN(new_n753));
  INV_X1    g552(.A(G92gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n747), .A2(new_n749), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n740), .A3(new_n737), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n758), .B2(new_n659), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n469), .B1(new_n738), .B2(new_n741), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n746), .B(new_n763), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n762), .A2(G92gat), .B1(new_n764), .B2(new_n756), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(new_n760), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n742), .B2(new_n513), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n294), .A2(new_n521), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n750), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n758), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n739), .A2(new_n740), .A3(KEYINPUT115), .A4(new_n737), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n487), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT117), .B1(new_n773), .B2(new_n298), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n459), .B1(new_n738), .B2(new_n741), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT117), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n718), .A2(G106gat), .A3(new_n487), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n764), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT53), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n747), .A2(new_n749), .A3(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n758), .B2(new_n487), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT118), .Z(new_n786));
  NAND2_X1  g585(.A1(new_n781), .A2(new_n786), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788));
  INV_X1    g587(.A(new_n552), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n548), .A2(new_n520), .A3(new_n551), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n559), .B1(new_n552), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n554), .A2(new_n558), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n791), .B2(new_n793), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n587), .A2(new_n589), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n588), .B1(new_n597), .B2(new_n585), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n606), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n610), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n674), .A2(new_n799), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n611), .A2(new_n613), .A3(new_n799), .ZN(new_n809));
  INV_X1    g608(.A(new_n803), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n562), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n652), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n629), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n720), .A2(new_n562), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n788), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n807), .A2(new_n799), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n652), .A3(new_n805), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n809), .A2(new_n811), .B1(new_n651), .B2(new_n650), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n673), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n815), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT120), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(new_n656), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n415), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n615), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G113gat), .ZN(G1340gat));
  INV_X1    g625(.A(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n827), .B2(new_n718), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n265), .A3(new_n562), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n629), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(G127gat), .ZN(G1342gat));
  INV_X1    g631(.A(G134gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n824), .A2(new_n833), .A3(new_n674), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n834), .A2(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n827), .B2(new_n652), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(KEYINPUT56), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n816), .A2(new_n822), .A3(new_n839), .A4(new_n656), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n512), .A2(new_n487), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n659), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n823), .A2(KEYINPUT122), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n614), .A2(G141gat), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT123), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n652), .B1(new_n812), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT121), .B1(new_n809), .B2(new_n811), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n808), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n815), .B1(new_n851), .B2(new_n673), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT57), .B1(new_n852), .B2(new_n487), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n816), .A2(new_n822), .A3(new_n854), .A4(new_n459), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n655), .A2(new_n469), .A3(new_n512), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(new_n615), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G141gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT58), .B1(new_n847), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n842), .B1(KEYINPUT122), .B2(new_n823), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n846), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1344gat));
  AOI21_X1  g664(.A(G148gat), .B1(new_n861), .B2(new_n562), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n563), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n816), .A2(new_n459), .A3(new_n822), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n851), .A2(new_n673), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n815), .B(KEYINPUT124), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n854), .B(new_n459), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n856), .A2(KEYINPUT59), .A3(new_n562), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n868), .A2(KEYINPUT59), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI22_X1  g675(.A1(KEYINPUT59), .A2(new_n866), .B1(new_n876), .B2(G148gat), .ZN(G1345gat));
  NAND4_X1  g676(.A1(new_n843), .A2(new_n301), .A3(new_n629), .A4(new_n844), .ZN(new_n878));
  OAI21_X1  g677(.A(G155gat), .B1(new_n867), .B2(new_n673), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT125), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n302), .A3(new_n652), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n861), .A2(new_n674), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n302), .ZN(G1347gat));
  NAND4_X1  g686(.A1(new_n816), .A2(new_n822), .A3(new_n372), .A4(new_n655), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n659), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n615), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(G169gat), .ZN(G1348gat));
  AOI21_X1  g690(.A(G176gat), .B1(new_n889), .B2(new_n562), .ZN(new_n892));
  INV_X1    g691(.A(G176gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n892), .B1(new_n753), .B2(new_n894), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n888), .A2(new_n673), .A3(new_n659), .ZN(new_n896));
  INV_X1    g695(.A(new_n248), .ZN(new_n897));
  INV_X1    g696(.A(new_n254), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n899), .B1(new_n250), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n899), .B(new_n902), .C1(new_n250), .C2(new_n896), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  NAND2_X1  g703(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(KEYINPUT61), .B(G190gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n674), .ZN(new_n907));
  MUX2_X1   g706(.A(new_n905), .B(new_n906), .S(new_n907), .Z(G1351gat));
  NOR3_X1   g707(.A1(new_n656), .A2(new_n659), .A3(new_n512), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT126), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n870), .A2(new_n873), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n614), .ZN(new_n912));
  INV_X1    g711(.A(new_n869), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n909), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n603), .A3(new_n615), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(G1352gat));
  INV_X1    g715(.A(G204gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n917), .A3(new_n562), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n911), .B2(new_n718), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1353gat));
  NAND2_X1  g721(.A1(new_n909), .A2(new_n629), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n870), .A2(new_n873), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(G211gat), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n926), .A2(new_n927), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n329), .A3(new_n924), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n930), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G1354gat));
  INV_X1    g733(.A(new_n331), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n911), .A2(new_n652), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G218gat), .B1(new_n914), .B2(new_n674), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1355gat));
endmodule


