

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794;

  NAND2_X1 U374 ( .A1(n403), .A2(n402), .ZN(n505) );
  AND2_X1 U375 ( .A1(n398), .A2(n404), .ZN(n403) );
  NOR2_X1 U376 ( .A1(n699), .A2(n499), .ZN(n647) );
  BUF_X1 U377 ( .A(n468), .Z(n354) );
  NOR2_X1 U378 ( .A1(n629), .A2(n630), .ZN(n631) );
  BUF_X1 U379 ( .A(n694), .Z(n468) );
  XNOR2_X1 U380 ( .A(n694), .B(n473), .ZN(n624) );
  NAND2_X1 U381 ( .A1(G214), .A2(n540), .ZN(n700) );
  OR2_X1 U382 ( .A1(n657), .A2(G902), .ZN(n482) );
  XNOR2_X1 U383 ( .A(n532), .B(n487), .ZN(n766) );
  XNOR2_X1 U384 ( .A(n546), .B(KEYINPUT16), .ZN(n487) );
  BUF_X1 U385 ( .A(G107), .Z(n353) );
  XOR2_X1 U386 ( .A(G143), .B(G128), .Z(n535) );
  XNOR2_X1 U387 ( .A(n478), .B(G101), .ZN(n534) );
  INV_X4 U388 ( .A(G953), .ZN(n784) );
  INV_X1 U389 ( .A(KEYINPUT4), .ZN(n478) );
  XNOR2_X2 U390 ( .A(n538), .B(KEYINPUT90), .ZN(n514) );
  XNOR2_X2 U391 ( .A(KEYINPUT15), .B(G902), .ZN(n656) );
  INV_X2 U392 ( .A(KEYINPUT0), .ZN(n432) );
  XNOR2_X2 U393 ( .A(n352), .B(n574), .ZN(n476) );
  NAND2_X2 U394 ( .A1(n433), .A2(n573), .ZN(n352) );
  XNOR2_X2 U395 ( .A(n516), .B(KEYINPUT69), .ZN(n367) );
  XNOR2_X1 U396 ( .A(n367), .B(G137), .ZN(n463) );
  XNOR2_X1 U397 ( .A(n535), .B(n462), .ZN(n547) );
  AND2_X1 U398 ( .A1(n387), .A2(n492), .ZN(n725) );
  NOR2_X1 U399 ( .A1(n794), .A2(n442), .ZN(n648) );
  NOR2_X1 U400 ( .A1(n675), .A2(n382), .ZN(n596) );
  OR2_X1 U401 ( .A1(n641), .A2(n355), .ZN(n515) );
  AND2_X1 U402 ( .A1(n505), .A2(n504), .ZN(n782) );
  AND2_X1 U403 ( .A1(n407), .A2(n506), .ZN(n401) );
  OR2_X1 U404 ( .A1(n669), .A2(n791), .ZN(n448) );
  XNOR2_X1 U405 ( .A(n606), .B(KEYINPUT35), .ZN(n788) );
  AND2_X1 U406 ( .A1(n428), .A2(n427), .ZN(n391) );
  AND2_X1 U407 ( .A1(n376), .A2(n500), .ZN(n443) );
  XNOR2_X1 U408 ( .A(n648), .B(KEYINPUT46), .ZN(n428) );
  XNOR2_X1 U409 ( .A(n513), .B(n512), .ZN(n791) );
  AND2_X1 U410 ( .A1(n672), .A2(n363), .ZN(n638) );
  XNOR2_X1 U411 ( .A(n645), .B(KEYINPUT40), .ZN(n794) );
  XNOR2_X1 U412 ( .A(n408), .B(KEYINPUT107), .ZN(n789) );
  AND2_X1 U413 ( .A1(n425), .A2(n675), .ZN(n645) );
  AND2_X1 U414 ( .A1(n637), .A2(n364), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n467), .B(n619), .ZN(n701) );
  INV_X1 U416 ( .A(n685), .ZN(n355) );
  XNOR2_X1 U417 ( .A(G475), .B(n567), .ZN(n603) );
  XNOR2_X1 U418 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U419 ( .A(n501), .B(n587), .ZN(n756) );
  XNOR2_X1 U420 ( .A(n366), .B(n556), .ZN(n559) );
  XNOR2_X1 U421 ( .A(n767), .B(n477), .ZN(n578) );
  XNOR2_X1 U422 ( .A(n534), .B(KEYINPUT73), .ZN(n477) );
  XNOR2_X1 U423 ( .A(n533), .B(G110), .ZN(n767) );
  XNOR2_X1 U424 ( .A(n580), .B(n579), .ZN(n485) );
  XNOR2_X1 U425 ( .A(n497), .B(G146), .ZN(n561) );
  NAND2_X1 U426 ( .A1(n362), .A2(n407), .ZN(n399) );
  NAND2_X1 U427 ( .A1(n391), .A2(n443), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n356), .B(n490), .ZN(n358) );
  XNOR2_X1 U429 ( .A(n531), .B(n530), .ZN(n356) );
  NAND2_X1 U430 ( .A1(n359), .A2(n357), .ZN(n488) );
  NAND2_X1 U431 ( .A1(n358), .A2(n489), .ZN(n357) );
  NAND2_X1 U432 ( .A1(n392), .A2(n360), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n361), .B(n529), .ZN(n360) );
  XNOR2_X1 U434 ( .A(n386), .B(n530), .ZN(n361) );
  AND2_X1 U435 ( .A1(n362), .A2(n405), .ZN(n400) );
  NAND2_X1 U436 ( .A1(n672), .A2(n637), .ZN(n365) );
  INV_X1 U437 ( .A(KEYINPUT47), .ZN(n364) );
  NAND2_X1 U438 ( .A1(n365), .A2(KEYINPUT47), .ZN(n642) );
  INV_X1 U439 ( .A(n367), .ZN(n366) );
  AND2_X1 U440 ( .A1(n650), .A2(n701), .ZN(n368) );
  XNOR2_X1 U441 ( .A(n397), .B(n378), .ZN(n435) );
  NAND2_X1 U442 ( .A1(n632), .A2(n370), .ZN(n371) );
  NAND2_X1 U443 ( .A1(n369), .A2(n485), .ZN(n372) );
  NAND2_X1 U444 ( .A1(n371), .A2(n372), .ZN(n379) );
  INV_X1 U445 ( .A(n632), .ZN(n369) );
  INV_X1 U446 ( .A(n485), .ZN(n370) );
  XNOR2_X1 U447 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n373) );
  XNOR2_X1 U448 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n457) );
  XNOR2_X2 U449 ( .A(n374), .B(n432), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n635), .A2(n541), .ZN(n374) );
  NAND2_X1 U451 ( .A1(n635), .A2(n541), .ZN(n440) );
  AND2_X2 U452 ( .A1(n493), .A2(n491), .ZN(n385) );
  XNOR2_X2 U453 ( .A(n486), .B(n377), .ZN(n632) );
  INV_X1 U454 ( .A(G146), .ZN(n517) );
  INV_X1 U455 ( .A(KEYINPUT22), .ZN(n574) );
  OR2_X1 U456 ( .A1(n644), .A2(n625), .ZN(n639) );
  NOR2_X1 U457 ( .A1(n629), .A2(n475), .ZN(n474) );
  INV_X1 U458 ( .A(n700), .ZN(n475) );
  INV_X1 U459 ( .A(KEYINPUT74), .ZN(n424) );
  XNOR2_X1 U460 ( .A(n561), .B(KEYINPUT87), .ZN(n489) );
  INV_X1 U461 ( .A(n688), .ZN(n419) );
  OR2_X1 U462 ( .A1(G237), .A2(G902), .ZN(n540) );
  XNOR2_X1 U463 ( .A(n591), .B(n590), .ZN(n621) );
  NOR2_X1 U464 ( .A1(G902), .A2(n756), .ZN(n591) );
  INV_X1 U465 ( .A(n682), .ZN(n504) );
  XNOR2_X1 U466 ( .A(n520), .B(n519), .ZN(n532) );
  XNOR2_X2 U467 ( .A(G113), .B(G116), .ZN(n518) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n557) );
  INV_X1 U469 ( .A(n725), .ZN(n491) );
  INV_X1 U470 ( .A(G902), .ZN(n434) );
  BUF_X1 U471 ( .A(n621), .Z(n685) );
  XNOR2_X1 U472 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n473) );
  XNOR2_X1 U473 ( .A(n503), .B(n584), .ZN(n459) );
  XOR2_X1 U474 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n584) );
  XNOR2_X1 U475 ( .A(n586), .B(KEYINPUT23), .ZN(n503) );
  XNOR2_X1 U476 ( .A(G119), .B(G128), .ZN(n586) );
  INV_X1 U477 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U478 ( .A(G113), .B(G143), .ZN(n552) );
  XOR2_X1 U479 ( .A(G104), .B(G122), .Z(n553) );
  XNOR2_X1 U480 ( .A(KEYINPUT11), .B(KEYINPUT97), .ZN(n554) );
  XOR2_X1 U481 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n555) );
  XNOR2_X1 U482 ( .A(n562), .B(KEYINPUT10), .ZN(n774) );
  NAND2_X1 U483 ( .A1(n651), .A2(n422), .ZN(n411) );
  NOR2_X1 U484 ( .A1(G902), .A2(n747), .ZN(n566) );
  OR2_X1 U485 ( .A1(n628), .A2(n422), .ZN(n429) );
  NOR2_X1 U486 ( .A1(n641), .A2(n626), .ZN(n627) );
  NAND2_X1 U487 ( .A1(n430), .A2(n429), .ZN(n406) );
  NAND2_X1 U488 ( .A1(n431), .A2(n655), .ZN(n430) );
  NOR2_X1 U489 ( .A1(n600), .A2(KEYINPUT85), .ZN(n453) );
  INV_X1 U490 ( .A(KEYINPUT82), .ZN(n507) );
  XNOR2_X1 U491 ( .A(n440), .B(n432), .ZN(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n542) );
  INV_X1 U493 ( .A(G125), .ZN(n497) );
  XOR2_X1 U494 ( .A(n353), .B(G140), .Z(n576) );
  NAND2_X1 U495 ( .A1(n375), .A2(n413), .ZN(n412) );
  INV_X1 U496 ( .A(KEYINPUT30), .ZN(n460) );
  NAND2_X1 U497 ( .A1(n355), .A2(n495), .ZN(n629) );
  NOR2_X1 U498 ( .A1(n622), .A2(n496), .ZN(n495) );
  INV_X1 U499 ( .A(n623), .ZN(n496) );
  XNOR2_X1 U500 ( .A(n397), .B(n483), .ZN(n657) );
  XNOR2_X1 U501 ( .A(n523), .B(n484), .ZN(n483) );
  INV_X1 U502 ( .A(n532), .ZN(n484) );
  AND2_X1 U503 ( .A1(n761), .A2(KEYINPUT2), .ZN(n492) );
  NOR2_X1 U504 ( .A1(n707), .A2(n704), .ZN(n646) );
  NOR2_X1 U505 ( .A1(n688), .A2(n389), .ZN(n650) );
  XNOR2_X1 U506 ( .A(n502), .B(n774), .ZN(n501) );
  XNOR2_X1 U507 ( .A(n459), .B(n585), .ZN(n502) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n753) );
  XNOR2_X1 U509 ( .A(n446), .B(n548), .ZN(n445) );
  XNOR2_X1 U510 ( .A(n560), .B(n558), .ZN(n464) );
  NOR2_X1 U511 ( .A1(G952), .A2(n784), .ZN(n760) );
  NOR2_X1 U512 ( .A1(n639), .A2(n640), .ZN(n472) );
  BUF_X1 U513 ( .A(n788), .Z(n458) );
  XNOR2_X1 U514 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n512) );
  NAND2_X1 U515 ( .A1(n409), .A2(n653), .ZN(n408) );
  XNOR2_X1 U516 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U517 ( .A(KEYINPUT106), .ZN(n410) );
  AND2_X1 U518 ( .A1(n634), .A2(n498), .ZN(n672) );
  NOR2_X1 U519 ( .A1(n636), .A2(n389), .ZN(n498) );
  INV_X1 U520 ( .A(n429), .ZN(n683) );
  AND2_X1 U521 ( .A1(n419), .A2(KEYINPUT33), .ZN(n375) );
  AND2_X1 U522 ( .A1(n643), .A2(n423), .ZN(n376) );
  XOR2_X1 U523 ( .A(KEYINPUT72), .B(G469), .Z(n377) );
  XOR2_X1 U524 ( .A(n578), .B(n577), .Z(n378) );
  INV_X1 U525 ( .A(n624), .ZN(n416) );
  AND2_X1 U526 ( .A1(n453), .A2(n456), .ZN(n380) );
  NOR2_X1 U527 ( .A1(n669), .A2(n791), .ZN(n381) );
  INV_X1 U528 ( .A(KEYINPUT33), .ZN(n418) );
  AND2_X1 U529 ( .A1(n595), .A2(n603), .ZN(n382) );
  XOR2_X1 U530 ( .A(n657), .B(KEYINPUT62), .Z(n383) );
  INV_X1 U531 ( .A(KEYINPUT83), .ZN(n506) );
  OR2_X1 U532 ( .A1(n656), .A2(n719), .ZN(n384) );
  INV_X1 U533 ( .A(n457), .ZN(n386) );
  INV_X1 U534 ( .A(n373), .ZN(n531) );
  BUF_X1 U535 ( .A(n467), .Z(n422) );
  AND2_X1 U536 ( .A1(n505), .A2(n504), .ZN(n387) );
  XNOR2_X1 U537 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U538 ( .A(n632), .B(n485), .ZN(n388) );
  XNOR2_X1 U539 ( .A(n486), .B(n377), .ZN(n389) );
  NAND2_X1 U540 ( .A1(n400), .A2(n401), .ZN(n402) );
  NAND2_X1 U541 ( .A1(n406), .A2(KEYINPUT83), .ZN(n404) );
  BUF_X1 U542 ( .A(n710), .Z(n390) );
  NAND2_X1 U543 ( .A1(n414), .A2(n412), .ZN(n710) );
  BUF_X1 U544 ( .A(n652), .Z(n467) );
  BUF_X1 U545 ( .A(n388), .Z(n465) );
  AND2_X1 U546 ( .A1(n456), .A2(n466), .ZN(n438) );
  NAND2_X1 U547 ( .A1(n788), .A2(KEYINPUT44), .ZN(n456) );
  INV_X1 U548 ( .A(n489), .ZN(n392) );
  NAND2_X1 U549 ( .A1(n581), .A2(G217), .ZN(n444) );
  NOR2_X1 U550 ( .A1(n609), .A2(n608), .ZN(n513) );
  BUF_X1 U551 ( .A(n435), .Z(n393) );
  BUF_X1 U552 ( .A(n735), .Z(n395) );
  INV_X1 U553 ( .A(n396), .ZN(n790) );
  NAND2_X1 U554 ( .A1(n438), .A2(n396), .ZN(n437) );
  XNOR2_X2 U555 ( .A(n593), .B(KEYINPUT103), .ZN(n396) );
  NAND2_X1 U556 ( .A1(n396), .A2(n380), .ZN(n439) );
  XNOR2_X2 U557 ( .A(n773), .B(n517), .ZN(n397) );
  NAND2_X1 U558 ( .A1(n399), .A2(KEYINPUT83), .ZN(n398) );
  INV_X1 U559 ( .A(n406), .ZN(n405) );
  NAND2_X1 U560 ( .A1(n426), .A2(n655), .ZN(n407) );
  NOR2_X1 U561 ( .A1(n624), .A2(n388), .ZN(n413) );
  NAND2_X1 U562 ( .A1(n415), .A2(n418), .ZN(n414) );
  NAND2_X1 U563 ( .A1(n417), .A2(n416), .ZN(n415) );
  INV_X1 U564 ( .A(n447), .ZN(n417) );
  NOR2_X2 U565 ( .A1(n710), .A2(n601), .ZN(n602) );
  NAND2_X1 U566 ( .A1(n379), .A2(n419), .ZN(n447) );
  NAND2_X1 U567 ( .A1(n448), .A2(KEYINPUT44), .ZN(n452) );
  XNOR2_X1 U568 ( .A(n461), .B(n460), .ZN(n618) );
  NAND2_X1 U569 ( .A1(n435), .A2(n434), .ZN(n486) );
  NAND2_X1 U570 ( .A1(n421), .A2(n611), .ZN(n454) );
  NAND2_X1 U571 ( .A1(n452), .A2(n449), .ZN(n421) );
  XNOR2_X1 U572 ( .A(n559), .B(n464), .ZN(n564) );
  XNOR2_X1 U573 ( .A(n638), .B(n424), .ZN(n423) );
  AND2_X1 U574 ( .A1(n425), .A2(n382), .ZN(n682) );
  XNOR2_X1 U575 ( .A(n620), .B(KEYINPUT39), .ZN(n425) );
  NAND2_X1 U576 ( .A1(n428), .A2(n427), .ZN(n426) );
  XNOR2_X1 U577 ( .A(n789), .B(KEYINPUT77), .ZN(n427) );
  INV_X1 U578 ( .A(n376), .ZN(n431) );
  INV_X1 U579 ( .A(n394), .ZN(n601) );
  NAND2_X1 U580 ( .A1(n394), .A2(n650), .ZN(n598) );
  NAND2_X1 U581 ( .A1(n394), .A2(n696), .ZN(n597) );
  XNOR2_X1 U582 ( .A(n393), .B(n742), .ZN(n744) );
  NAND2_X1 U583 ( .A1(n436), .A2(n439), .ZN(n455) );
  NAND2_X1 U584 ( .A1(n437), .A2(KEYINPUT85), .ZN(n436) );
  XNOR2_X2 U585 ( .A(n441), .B(KEYINPUT19), .ZN(n635) );
  NAND2_X2 U586 ( .A1(n652), .A2(n700), .ZN(n441) );
  XNOR2_X1 U587 ( .A(n442), .B(n793), .ZN(G39) );
  XNOR2_X1 U588 ( .A(n647), .B(KEYINPUT42), .ZN(n442) );
  XNOR2_X1 U589 ( .A(n549), .B(n550), .ZN(n446) );
  NOR2_X1 U590 ( .A1(n753), .A2(G902), .ZN(n551) );
  NOR2_X1 U591 ( .A1(n447), .A2(n630), .ZN(n696) );
  NAND2_X1 U592 ( .A1(n451), .A2(n450), .ZN(n449) );
  INV_X1 U593 ( .A(n669), .ZN(n450) );
  NOR2_X1 U594 ( .A1(n791), .A2(KEYINPUT44), .ZN(n451) );
  NAND2_X1 U595 ( .A1(n454), .A2(n455), .ZN(n612) );
  XNOR2_X1 U596 ( .A(n537), .B(n536), .ZN(n735) );
  NAND2_X1 U597 ( .A1(n694), .A2(n700), .ZN(n461) );
  XNOR2_X2 U598 ( .A(n482), .B(G472), .ZN(n694) );
  INV_X1 U599 ( .A(n529), .ZN(n490) );
  XNOR2_X1 U600 ( .A(n736), .B(n737), .ZN(n738) );
  NAND2_X1 U601 ( .A1(n701), .A2(n700), .ZN(n707) );
  NAND2_X1 U602 ( .A1(n479), .A2(n384), .ZN(n493) );
  XNOR2_X1 U603 ( .A(n609), .B(KEYINPUT84), .ZN(n592) );
  XNOR2_X1 U604 ( .A(n612), .B(KEYINPUT45), .ZN(n718) );
  NAND2_X1 U605 ( .A1(n368), .A2(n649), .ZN(n620) );
  XNOR2_X1 U606 ( .A(n646), .B(KEYINPUT41), .ZN(n699) );
  XNOR2_X1 U607 ( .A(n480), .B(n494), .ZN(n479) );
  XNOR2_X1 U608 ( .A(n488), .B(n766), .ZN(n537) );
  XNOR2_X2 U609 ( .A(n463), .B(n547), .ZN(n773) );
  NAND2_X1 U610 ( .A1(n385), .A2(G210), .ZN(n736) );
  INV_X1 U611 ( .A(n600), .ZN(n466) );
  XNOR2_X1 U612 ( .A(n469), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U613 ( .A1(n750), .A2(n760), .ZN(n469) );
  XNOR2_X1 U614 ( .A(n470), .B(KEYINPUT122), .ZN(G66) );
  NOR2_X2 U615 ( .A1(n759), .A2(n760), .ZN(n470) );
  AND2_X1 U616 ( .A1(n681), .A2(n642), .ZN(n643) );
  NAND2_X1 U617 ( .A1(n471), .A2(n641), .ZN(n681) );
  XNOR2_X1 U618 ( .A(n472), .B(KEYINPUT36), .ZN(n471) );
  NAND2_X1 U619 ( .A1(n474), .A2(n416), .ZN(n625) );
  NAND2_X1 U620 ( .A1(n476), .A2(n624), .ZN(n609) );
  NAND2_X1 U621 ( .A1(n476), .A2(n465), .ZN(n610) );
  NAND2_X1 U622 ( .A1(n481), .A2(n782), .ZN(n480) );
  XNOR2_X1 U623 ( .A(n508), .B(n507), .ZN(n481) );
  NAND2_X1 U624 ( .A1(n385), .A2(G217), .ZN(n758) );
  INV_X1 U625 ( .A(KEYINPUT81), .ZN(n494) );
  XNOR2_X2 U626 ( .A(G131), .B(KEYINPUT70), .ZN(n516) );
  NOR2_X2 U627 ( .A1(n738), .A2(n760), .ZN(n739) );
  NAND2_X1 U628 ( .A1(n634), .A2(n633), .ZN(n499) );
  INV_X1 U629 ( .A(n655), .ZN(n500) );
  NAND2_X1 U630 ( .A1(n718), .A2(n613), .ZN(n508) );
  AND2_X2 U631 ( .A1(n509), .A2(n355), .ZN(n669) );
  XNOR2_X1 U632 ( .A(n511), .B(n510), .ZN(n509) );
  INV_X1 U633 ( .A(KEYINPUT65), .ZN(n510) );
  NOR2_X2 U634 ( .A1(n610), .A2(n354), .ZN(n511) );
  XNOR2_X2 U635 ( .A(n539), .B(n514), .ZN(n652) );
  BUF_X1 U636 ( .A(n385), .Z(n751) );
  BUF_X1 U637 ( .A(n718), .Z(n761) );
  INV_X1 U638 ( .A(KEYINPUT48), .ZN(n654) );
  XNOR2_X1 U639 ( .A(n654), .B(KEYINPUT71), .ZN(n655) );
  XNOR2_X1 U640 ( .A(n589), .B(KEYINPUT25), .ZN(n590) );
  INV_X1 U641 ( .A(n760), .ZN(n659) );
  XNOR2_X1 U642 ( .A(n749), .B(n748), .ZN(n750) );
  INV_X1 U643 ( .A(n656), .ZN(n613) );
  INV_X1 U644 ( .A(n518), .ZN(n520) );
  XNOR2_X1 U645 ( .A(KEYINPUT3), .B(G119), .ZN(n519) );
  XOR2_X1 U646 ( .A(n534), .B(KEYINPUT5), .Z(n522) );
  NAND2_X1 U647 ( .A1(n557), .A2(G210), .ZN(n521) );
  XNOR2_X1 U648 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X1 U649 ( .A1(G898), .A2(n784), .ZN(n770) );
  NAND2_X1 U650 ( .A1(G234), .A2(G237), .ZN(n524) );
  XNOR2_X1 U651 ( .A(n524), .B(KEYINPUT14), .ZN(n526) );
  NAND2_X1 U652 ( .A1(G902), .A2(n526), .ZN(n614) );
  INV_X1 U653 ( .A(n614), .ZN(n525) );
  NAND2_X1 U654 ( .A1(n770), .A2(n525), .ZN(n528) );
  NAND2_X1 U655 ( .A1(G952), .A2(n526), .ZN(n717) );
  NOR2_X1 U656 ( .A1(n717), .A2(G953), .ZN(n527) );
  XNOR2_X1 U657 ( .A(n527), .B(KEYINPUT91), .ZN(n617) );
  NAND2_X1 U658 ( .A1(n528), .A2(n617), .ZN(n541) );
  AND2_X1 U659 ( .A1(G224), .A2(n784), .ZN(n529) );
  XNOR2_X2 U660 ( .A(KEYINPUT76), .B(KEYINPUT89), .ZN(n530) );
  XOR2_X2 U661 ( .A(G122), .B(G107), .Z(n546) );
  XNOR2_X1 U662 ( .A(G104), .B(KEYINPUT88), .ZN(n533) );
  XNOR2_X1 U663 ( .A(n535), .B(n578), .ZN(n536) );
  NAND2_X1 U664 ( .A1(n735), .A2(n656), .ZN(n539) );
  AND2_X1 U665 ( .A1(G210), .A2(n540), .ZN(n538) );
  XNOR2_X1 U666 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n550) );
  XNOR2_X1 U667 ( .A(n542), .B(KEYINPUT79), .ZN(n543) );
  XOR2_X1 U668 ( .A(KEYINPUT68), .B(n543), .Z(n545) );
  NAND2_X1 U669 ( .A1(G234), .A2(n784), .ZN(n544) );
  XNOR2_X1 U670 ( .A(n545), .B(n544), .ZN(n581) );
  XOR2_X1 U671 ( .A(KEYINPUT100), .B(n546), .Z(n549) );
  XNOR2_X1 U672 ( .A(G116), .B(n547), .ZN(n548) );
  XOR2_X1 U673 ( .A(G478), .B(n551), .Z(n595) );
  INV_X1 U674 ( .A(n595), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n553), .B(n552), .ZN(n560) );
  XNOR2_X1 U676 ( .A(n555), .B(n554), .ZN(n556) );
  NAND2_X1 U677 ( .A1(G214), .A2(n557), .ZN(n558) );
  XNOR2_X1 U678 ( .A(n561), .B(G140), .ZN(n562) );
  INV_X1 U679 ( .A(n774), .ZN(n563) );
  XNOR2_X1 U680 ( .A(n564), .B(n563), .ZN(n747) );
  XNOR2_X1 U681 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n565) );
  XNOR2_X1 U682 ( .A(n566), .B(n565), .ZN(n567) );
  NAND2_X1 U683 ( .A1(n604), .A2(n603), .ZN(n704) );
  XOR2_X1 U684 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n571) );
  NAND2_X1 U685 ( .A1(n656), .A2(G234), .ZN(n568) );
  XNOR2_X1 U686 ( .A(n568), .B(KEYINPUT20), .ZN(n569) );
  XNOR2_X1 U687 ( .A(KEYINPUT94), .B(n569), .ZN(n588) );
  NAND2_X1 U688 ( .A1(G221), .A2(n588), .ZN(n570) );
  XNOR2_X1 U689 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U690 ( .A(KEYINPUT21), .B(n572), .Z(n686) );
  INV_X1 U691 ( .A(n686), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n704), .A2(n622), .ZN(n573) );
  NAND2_X1 U693 ( .A1(G227), .A2(n784), .ZN(n575) );
  XNOR2_X1 U694 ( .A(n576), .B(n575), .ZN(n577) );
  INV_X1 U695 ( .A(KEYINPUT1), .ZN(n579) );
  INV_X1 U696 ( .A(KEYINPUT66), .ZN(n580) );
  INV_X1 U697 ( .A(n465), .ZN(n641) );
  NAND2_X1 U698 ( .A1(G221), .A2(n581), .ZN(n587) );
  XOR2_X1 U699 ( .A(KEYINPUT78), .B(KEYINPUT93), .Z(n583) );
  XNOR2_X1 U700 ( .A(G137), .B(G110), .ZN(n582) );
  XNOR2_X1 U701 ( .A(n583), .B(n582), .ZN(n585) );
  NAND2_X1 U702 ( .A1(G217), .A2(n588), .ZN(n589) );
  NOR2_X2 U703 ( .A1(n592), .A2(n515), .ZN(n593) );
  INV_X1 U704 ( .A(n603), .ZN(n594) );
  NAND2_X1 U705 ( .A1(n594), .A2(n604), .ZN(n644) );
  INV_X1 U706 ( .A(n644), .ZN(n675) );
  XNOR2_X1 U707 ( .A(n596), .B(KEYINPUT101), .ZN(n637) );
  INV_X1 U708 ( .A(n637), .ZN(n706) );
  INV_X1 U709 ( .A(n468), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n686), .A2(n621), .ZN(n688) );
  XNOR2_X1 U711 ( .A(KEYINPUT31), .B(n597), .ZN(n678) );
  NOR2_X1 U712 ( .A1(n354), .A2(n598), .ZN(n664) );
  NOR2_X1 U713 ( .A1(n678), .A2(n664), .ZN(n599) );
  NOR2_X1 U714 ( .A1(n706), .A2(n599), .ZN(n600) );
  XNOR2_X1 U715 ( .A(n602), .B(KEYINPUT34), .ZN(n605) );
  NOR2_X1 U716 ( .A1(n604), .A2(n603), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n605), .A2(n653), .ZN(n606) );
  NOR2_X1 U718 ( .A1(n465), .A2(n685), .ZN(n607) );
  XOR2_X1 U719 ( .A(KEYINPUT104), .B(n607), .Z(n608) );
  NAND2_X1 U720 ( .A1(n381), .A2(n458), .ZN(n611) );
  NOR2_X1 U721 ( .A1(G900), .A2(n614), .ZN(n615) );
  NAND2_X1 U722 ( .A1(G953), .A2(n615), .ZN(n616) );
  NAND2_X1 U723 ( .A1(n617), .A2(n616), .ZN(n623) );
  AND2_X1 U724 ( .A1(n623), .A2(n618), .ZN(n649) );
  XNOR2_X1 U725 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n619) );
  XOR2_X1 U726 ( .A(KEYINPUT105), .B(n639), .Z(n626) );
  XNOR2_X1 U727 ( .A(n627), .B(KEYINPUT43), .ZN(n628) );
  XNOR2_X1 U728 ( .A(n631), .B(KEYINPUT28), .ZN(n634) );
  INV_X1 U729 ( .A(n389), .ZN(n633) );
  INV_X1 U730 ( .A(n635), .ZN(n636) );
  INV_X1 U731 ( .A(n422), .ZN(n640) );
  AND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n719) );
  NAND2_X1 U734 ( .A1(G472), .A2(n385), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(n383), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U737 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U738 ( .A1(n664), .A2(n675), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n662), .B(KEYINPUT108), .ZN(n663) );
  XNOR2_X1 U740 ( .A(G104), .B(n663), .ZN(G6) );
  XOR2_X1 U741 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n666) );
  NAND2_X1 U742 ( .A1(n664), .A2(n382), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U744 ( .A(n353), .B(KEYINPUT26), .Z(n667) );
  XNOR2_X1 U745 ( .A(n668), .B(n667), .ZN(G9) );
  XOR2_X1 U746 ( .A(n669), .B(G110), .Z(G12) );
  XOR2_X1 U747 ( .A(G128), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U748 ( .A1(n672), .A2(n382), .ZN(n670) );
  XNOR2_X1 U749 ( .A(n671), .B(n670), .ZN(G30) );
  NAND2_X1 U750 ( .A1(n672), .A2(n675), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT110), .ZN(n674) );
  XNOR2_X1 U752 ( .A(G146), .B(n674), .ZN(G48) );
  XOR2_X1 U753 ( .A(G113), .B(KEYINPUT111), .Z(n677) );
  NAND2_X1 U754 ( .A1(n678), .A2(n675), .ZN(n676) );
  XNOR2_X1 U755 ( .A(n677), .B(n676), .ZN(G15) );
  NAND2_X1 U756 ( .A1(n678), .A2(n382), .ZN(n679) );
  XNOR2_X1 U757 ( .A(n679), .B(G116), .ZN(G18) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n680) );
  XNOR2_X1 U759 ( .A(n681), .B(n680), .ZN(G27) );
  XOR2_X1 U760 ( .A(G134), .B(n682), .Z(G36) );
  XOR2_X1 U761 ( .A(G140), .B(n683), .Z(G42) );
  XOR2_X1 U762 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n731) );
  NOR2_X1 U763 ( .A1(n699), .A2(n390), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G953), .A2(n684), .ZN(n729) );
  NOR2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U766 ( .A(KEYINPUT49), .B(n687), .ZN(n692) );
  NAND2_X1 U767 ( .A1(n688), .A2(n465), .ZN(n689) );
  XNOR2_X1 U768 ( .A(n689), .B(KEYINPUT112), .ZN(n690) );
  XNOR2_X1 U769 ( .A(KEYINPUT50), .B(n690), .ZN(n691) );
  NAND2_X1 U770 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n354), .A2(n693), .ZN(n695) );
  NOR2_X1 U772 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n697), .Z(n698) );
  NOR2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U776 ( .A(KEYINPUT113), .B(n702), .Z(n703) );
  NOR2_X1 U777 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U778 ( .A(n705), .B(KEYINPUT114), .ZN(n709) );
  NOR2_X1 U779 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U780 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U781 ( .A1(n711), .A2(n390), .ZN(n712) );
  NOR2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U783 ( .A(n714), .B(KEYINPUT52), .Z(n715) );
  XNOR2_X1 U784 ( .A(KEYINPUT115), .B(n715), .ZN(n716) );
  NOR2_X1 U785 ( .A1(n717), .A2(n716), .ZN(n727) );
  INV_X1 U786 ( .A(n761), .ZN(n720) );
  NAND2_X1 U787 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U788 ( .A(n721), .B(KEYINPUT80), .ZN(n723) );
  OR2_X1 U789 ( .A1(n387), .A2(KEYINPUT2), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U794 ( .A(n731), .B(n730), .ZN(G75) );
  XOR2_X1 U795 ( .A(KEYINPUT54), .B(KEYINPUT117), .Z(n733) );
  XNOR2_X1 U796 ( .A(KEYINPUT86), .B(KEYINPUT55), .ZN(n732) );
  XNOR2_X1 U797 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U798 ( .A(n395), .B(n734), .ZN(n737) );
  XNOR2_X1 U799 ( .A(n739), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U800 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n741) );
  XNOR2_X1 U801 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n740) );
  XNOR2_X1 U802 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U803 ( .A1(n751), .A2(G469), .ZN(n743) );
  XNOR2_X1 U804 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U805 ( .A1(n760), .A2(n745), .ZN(G54) );
  NAND2_X1 U806 ( .A1(n385), .A2(G475), .ZN(n749) );
  INV_X1 U807 ( .A(KEYINPUT59), .ZN(n746) );
  NAND2_X1 U808 ( .A1(G478), .A2(n751), .ZN(n752) );
  XNOR2_X1 U809 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U810 ( .A1(n760), .A2(n754), .ZN(G63) );
  XOR2_X1 U811 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n755) );
  XNOR2_X1 U812 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U813 ( .A1(n784), .A2(n761), .ZN(n765) );
  NAND2_X1 U814 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U815 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U816 ( .A1(n763), .A2(G898), .ZN(n764) );
  NAND2_X1 U817 ( .A1(n765), .A2(n764), .ZN(n772) );
  XNOR2_X1 U818 ( .A(G101), .B(n766), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(n767), .ZN(n769) );
  NOR2_X1 U820 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(G69) );
  BUF_X1 U822 ( .A(n773), .Z(n777) );
  XNOR2_X1 U823 ( .A(KEYINPUT4), .B(n774), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n775), .B(KEYINPUT123), .ZN(n776) );
  XOR2_X1 U825 ( .A(n777), .B(n776), .Z(n783) );
  XOR2_X1 U826 ( .A(G227), .B(n783), .Z(n778) );
  NAND2_X1 U827 ( .A1(n778), .A2(G900), .ZN(n779) );
  XOR2_X1 U828 ( .A(KEYINPUT124), .B(n779), .Z(n780) );
  NOR2_X1 U829 ( .A1(n784), .A2(n780), .ZN(n781) );
  XNOR2_X1 U830 ( .A(n781), .B(KEYINPUT125), .ZN(n787) );
  XNOR2_X1 U831 ( .A(n783), .B(n387), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U833 ( .A1(n787), .A2(n786), .ZN(G72) );
  XOR2_X1 U834 ( .A(n458), .B(G122), .Z(G24) );
  XOR2_X1 U835 ( .A(n789), .B(G143), .Z(G45) );
  XOR2_X1 U836 ( .A(n790), .B(G101), .Z(G3) );
  XOR2_X1 U837 ( .A(n791), .B(G119), .Z(n792) );
  XNOR2_X1 U838 ( .A(KEYINPUT126), .B(n792), .ZN(G21) );
  XNOR2_X1 U839 ( .A(G137), .B(KEYINPUT127), .ZN(n793) );
  XOR2_X1 U840 ( .A(n794), .B(G131), .Z(G33) );
endmodule

