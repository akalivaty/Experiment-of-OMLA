//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(G122), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT14), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT97), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G122), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(new_n188), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G107), .ZN(new_n197));
  INV_X1    g011(.A(new_n193), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n189), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(KEYINPUT95), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G128), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n202), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n202), .A3(new_n207), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT98), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n197), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n210), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n200), .B1(new_n214), .B2(new_n208), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n199), .B1(new_n191), .B2(new_n195), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT98), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT13), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n207), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n205), .A2(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(G134), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT96), .ZN(new_n224));
  OAI21_X1  g038(.A(G107), .B1(new_n188), .B2(new_n193), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n210), .A2(new_n224), .B1(new_n200), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n223), .B(new_n226), .C1(new_n224), .C2(new_n210), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT9), .B(G234), .ZN(new_n229));
  INV_X1    g043(.A(G217), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n229), .A2(new_n230), .A3(G953), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n218), .A2(new_n227), .A3(new_n231), .ZN(new_n234));
  AOI21_X1  g048(.A(G902), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G478), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT15), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n238), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(G475), .A2(G902), .ZN(new_n243));
  INV_X1    g057(.A(G140), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G125), .ZN(new_n245));
  INV_X1    g059(.A(G125), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G140), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT16), .ZN(new_n248));
  OR3_X1    g062(.A1(new_n246), .A2(KEYINPUT16), .A3(G140), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT75), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n248), .A2(new_n249), .A3(new_n252), .A4(G146), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n249), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G214), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(G143), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT17), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n261), .B(new_n262), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n258), .B(new_n264), .C1(new_n265), .C2(KEYINPUT17), .ZN(new_n266));
  XNOR2_X1  g080(.A(G113), .B(G122), .ZN(new_n267));
  INV_X1    g081(.A(G104), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(KEYINPUT18), .A2(G131), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n261), .B(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n245), .A2(new_n247), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(new_n255), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n255), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(KEYINPUT94), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n273), .A2(KEYINPUT94), .A3(new_n274), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n266), .A2(new_n269), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n272), .B(KEYINPUT19), .Z(new_n280));
  OAI211_X1 g094(.A(new_n265), .B(new_n250), .C1(G146), .C2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n269), .B1(new_n281), .B2(new_n277), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n243), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT20), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT20), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(new_n243), .C1(new_n279), .C2(new_n282), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n269), .B1(new_n266), .B2(new_n277), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n287), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n284), .A2(new_n286), .B1(G475), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(G234), .A2(G237), .ZN(new_n292));
  INV_X1    g106(.A(G953), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(G952), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(G902), .A3(G953), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT21), .B(G898), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n242), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  OR3_X1    g114(.A1(new_n192), .A2(KEYINPUT5), .A3(G119), .ZN(new_n301));
  XOR2_X1   g115(.A(G116), .B(G119), .Z(new_n302));
  INV_X1    g116(.A(KEYINPUT5), .ZN(new_n303));
  OAI211_X1 g117(.A(G113), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT2), .B(G113), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT82), .B(G101), .Z(new_n308));
  OAI21_X1  g122(.A(KEYINPUT3), .B1(new_n268), .B2(G107), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n268), .A2(G107), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n199), .A3(G104), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n199), .A2(G104), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G101), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n317), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT91), .B(KEYINPUT8), .Z(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G122), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n255), .A2(G143), .ZN(new_n326));
  INV_X1    g140(.A(G143), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(G143), .B2(new_n255), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n206), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G143), .B(G146), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n330), .A3(G128), .ZN(new_n334));
  AOI21_X1  g148(.A(G125), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(KEYINPUT0), .A2(G128), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT64), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT0), .B(G128), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n339), .A3(KEYINPUT64), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n335), .B1(G125), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G224), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G953), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT7), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n342), .A2(new_n346), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n322), .A2(new_n325), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT68), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n302), .A2(new_n305), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n306), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n302), .A2(KEYINPUT68), .A3(new_n305), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n309), .A2(new_n312), .A3(new_n310), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G101), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n358), .B2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n357), .A2(KEYINPUT83), .A3(new_n360), .A4(G101), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n313), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n355), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n324), .A3(new_n320), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n349), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n320), .ZN(new_n367));
  INV_X1    g181(.A(new_n324), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT90), .A2(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n342), .B(new_n344), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT90), .A2(KEYINPUT6), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G210), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n366), .A2(new_n375), .A3(new_n377), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT93), .A3(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(KEYINPUT93), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G214), .B1(G237), .B2(G902), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n385), .B(KEYINPUT89), .Z(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(G221), .B1(new_n229), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n389));
  INV_X1    g203(.A(G137), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G134), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT11), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT65), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT65), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT11), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(KEYINPUT65), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n202), .A2(G137), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n390), .A2(G134), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G131), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n394), .A2(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n397), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n202), .A2(G137), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n391), .A2(new_n406), .ZN(new_n407));
  AOI22_X1  g221(.A1(new_n391), .A2(new_n405), .B1(new_n407), .B2(new_n397), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n403), .B1(new_n408), .B2(new_n262), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n396), .A2(new_n400), .A3(new_n403), .A4(new_n262), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n402), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n329), .B1(new_n331), .B2(new_n203), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n334), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n313), .A3(new_n316), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n332), .A2(new_n334), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n317), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT12), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n389), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n419), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n412), .A2(new_n417), .A3(KEYINPUT85), .A4(KEYINPUT12), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G110), .B(G140), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n293), .A2(G227), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT10), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(new_n332), .B2(new_n334), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n415), .A2(new_n430), .B1(new_n317), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n362), .A2(new_n341), .A3(new_n363), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n396), .A2(new_n400), .A3(new_n262), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT66), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n435), .A2(new_n410), .B1(G131), .B2(new_n401), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT84), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT87), .A4(new_n422), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n425), .A2(new_n429), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n432), .A2(new_n433), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n412), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT88), .A3(new_n428), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n439), .A2(new_n440), .B1(new_n412), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n429), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n443), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G469), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n287), .ZN(new_n453));
  NAND2_X1  g267(.A1(G469), .A2(G902), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n441), .A2(new_n455), .A3(new_n423), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n441), .B2(new_n423), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n428), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n441), .A2(new_n429), .A3(new_n445), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(G469), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  AND4_X1   g275(.A1(new_n300), .A2(new_n387), .A3(new_n388), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n230), .B1(G234), .B2(new_n287), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n203), .A2(G119), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n206), .B2(G119), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT24), .B(G110), .Z(new_n466));
  OAI21_X1  g280(.A(KEYINPUT77), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT23), .B1(new_n203), .B2(G119), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(G110), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n465), .A2(KEYINPUT77), .A3(new_n466), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n250), .B(new_n274), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n471), .A2(G110), .B1(new_n465), .B2(new_n466), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n257), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n257), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n293), .A2(G221), .A3(G234), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT78), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G137), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n474), .B(new_n483), .C1(new_n477), .C2(new_n478), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT25), .B1(new_n487), .B2(new_n287), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n489), .B(G902), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n463), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT79), .B(new_n463), .C1(new_n488), .C2(new_n490), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n463), .A2(G902), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT80), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(KEYINPUT81), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT74), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n332), .A2(new_n334), .B1(G131), .B2(new_n407), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n503), .B1(new_n409), .B2(new_n411), .ZN(new_n504));
  INV_X1    g318(.A(new_n341), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n354), .C1(new_n436), .C2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g322(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n509));
  NAND2_X1  g323(.A1(new_n259), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(G101), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(KEYINPUT29), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n435), .A2(new_n410), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n505), .B1(new_n516), .B2(new_n402), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n407), .A2(G131), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n416), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n410), .B2(new_n435), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n355), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n506), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n412), .A2(new_n341), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(KEYINPUT69), .A3(new_n354), .A4(new_n504), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n523), .A2(KEYINPUT72), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT72), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n515), .B1(new_n528), .B2(KEYINPUT28), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT73), .B1(new_n529), .B2(G902), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(new_n525), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n523), .A2(new_n525), .A3(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n507), .B1(new_n536), .B2(new_n521), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n531), .B(new_n287), .C1(new_n537), .C2(new_n515), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n507), .B1(new_n523), .B2(new_n525), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n508), .A2(new_n521), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(new_n513), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n523), .A2(new_n525), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n524), .B2(new_n504), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n517), .A2(KEYINPUT30), .A3(new_n520), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n355), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n514), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n539), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n530), .A2(new_n538), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(new_n548), .A3(new_n514), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT31), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n513), .B1(new_n540), .B2(new_n541), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n544), .A2(new_n548), .A3(new_n556), .A4(new_n514), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G472), .A2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT32), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT32), .B1(new_n558), .B2(new_n559), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT71), .ZN(new_n567));
  AOI221_X4 g381(.A(new_n502), .B1(new_n552), .B2(G472), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n552), .A2(G472), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT74), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n462), .B(new_n501), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n572), .B(new_n308), .Z(G3));
  NAND2_X1  g387(.A1(new_n461), .A2(new_n388), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n558), .A2(new_n287), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n560), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n575), .A2(new_n500), .A3(new_n579), .A4(new_n499), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n236), .A2(new_n287), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n235), .B2(new_n236), .ZN(new_n582));
  INV_X1    g396(.A(new_n234), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n231), .B1(new_n218), .B2(new_n227), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT33), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n233), .A2(new_n586), .A3(new_n234), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(G478), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n291), .ZN(new_n590));
  INV_X1    g404(.A(new_n299), .ZN(new_n591));
  INV_X1    g405(.A(new_n386), .ZN(new_n592));
  INV_X1    g406(.A(new_n380), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n377), .B1(new_n366), .B2(new_n375), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  OR3_X1    g409(.A1(new_n590), .A2(new_n595), .A3(KEYINPUT99), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT99), .B1(new_n590), .B2(new_n595), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n580), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT34), .B(G104), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  INV_X1    g414(.A(new_n595), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n289), .A2(G475), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n286), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n284), .ZN(new_n605));
  INV_X1    g419(.A(new_n286), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n607), .B2(new_n603), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n601), .A2(new_n602), .A3(new_n242), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n580), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT35), .B(G107), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G9));
  NOR2_X1   g426(.A1(new_n483), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n479), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n496), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n493), .A2(new_n615), .A3(new_n494), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n300), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(new_n387), .A3(new_n575), .A4(new_n579), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT37), .B(G110), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G12));
  NAND2_X1  g434(.A1(new_n608), .A2(new_n242), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n294), .B(KEYINPUT101), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(new_n297), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n602), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n574), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n379), .A2(new_n380), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n616), .A2(new_n592), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n628), .B(new_n630), .C1(new_n568), .C2(new_n571), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  XOR2_X1   g446(.A(new_n384), .B(KEYINPUT38), .Z(new_n633));
  AOI21_X1  g447(.A(new_n290), .B1(new_n240), .B2(new_n241), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n592), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n616), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n625), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n575), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n640), .A2(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n549), .A2(new_n514), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n287), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n528), .A2(new_n514), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n569), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n637), .A2(new_n641), .A3(new_n642), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n327), .ZN(G45));
  NOR2_X1   g464(.A1(new_n590), .A2(new_n625), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n574), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n630), .B(new_n653), .C1(new_n568), .C2(new_n571), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n566), .A3(KEYINPUT71), .ZN(new_n658));
  INV_X1    g472(.A(new_n567), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n570), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n502), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n569), .A2(KEYINPUT74), .A3(new_n570), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n663), .A2(KEYINPUT103), .A3(new_n630), .A4(new_n653), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  AOI21_X1  g480(.A(new_n452), .B1(new_n451), .B2(new_n287), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n388), .A3(new_n453), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n596), .B2(new_n597), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n501), .C1(new_n568), .C2(new_n571), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT41), .B(G113), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G15));
  NOR2_X1   g487(.A1(new_n609), .A2(new_n669), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n674), .B(new_n501), .C1(new_n568), .C2(new_n571), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G116), .ZN(G18));
  NAND2_X1  g490(.A1(new_n629), .A2(new_n592), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n617), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(new_n661), .B2(new_n662), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(G119), .Z(G21));
  INV_X1    g495(.A(new_n453), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n667), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n601), .A3(new_n388), .A4(new_n634), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n537), .B1(new_n507), .B2(new_n506), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n554), .B(new_n557), .C1(new_n685), .C2(new_n514), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n559), .B(KEYINPUT104), .Z(new_n687));
  AOI22_X1  g501(.A1(new_n686), .A2(new_n687), .B1(G472), .B2(new_n576), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n498), .B(KEYINPUT105), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n684), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n187), .ZN(G24));
  AND2_X1   g509(.A1(new_n688), .A2(new_n616), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n651), .A3(new_n678), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  AOI211_X1 g512(.A(new_n566), .B(new_n657), .C1(new_n552), .C2(G472), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n498), .B(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  OR3_X1    g516(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n699), .B2(new_n701), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n384), .A2(new_n592), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n651), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT107), .B1(new_n461), .B2(new_n388), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n461), .A2(KEYINPUT107), .A3(new_n388), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n708), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n711), .A2(new_n706), .A3(new_n710), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n501), .B(new_n715), .C1(new_n568), .C2(new_n571), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n709), .B1(new_n716), .B2(new_n652), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g533(.A(KEYINPUT108), .B(new_n709), .C1(new_n716), .C2(new_n652), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n262), .ZN(G33));
  NOR2_X1   g536(.A1(new_n621), .A2(new_n627), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n663), .A2(new_n501), .A3(new_n723), .A4(new_n715), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(new_n388), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n458), .A2(new_n459), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n452), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n728), .B2(new_n727), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT46), .B1(new_n730), .B2(new_n454), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n682), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n454), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n726), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n582), .A2(new_n588), .A3(new_n290), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT43), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT43), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n578), .A3(new_n616), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n706), .B1(new_n740), .B2(new_n741), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n734), .A2(new_n742), .A3(new_n639), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G137), .ZN(G39));
  NOR3_X1   g559(.A1(new_n663), .A2(new_n501), .A3(new_n708), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  AOI211_X1 g562(.A(new_n748), .B(new_n726), .C1(new_n732), .C2(new_n733), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G140), .ZN(G42));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n623), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT113), .Z(new_n753));
  NOR2_X1   g567(.A1(new_n706), .A2(new_n669), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n705), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT48), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n648), .A2(new_n501), .A3(new_n295), .A4(new_n754), .ZN(new_n758));
  OAI211_X1 g572(.A(G952), .B(new_n293), .C1(new_n758), .C2(new_n590), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n691), .A2(new_n693), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n759), .B1(new_n761), .B2(new_n678), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n633), .A2(new_n592), .A3(new_n669), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n753), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n758), .A2(new_n291), .A3(new_n589), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n696), .B2(new_n755), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n747), .A2(new_n749), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n683), .A2(new_n726), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT115), .Z(new_n775));
  NOR3_X1   g589(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n761), .A2(new_n707), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n763), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n774), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n707), .B(new_n761), .C1(new_n771), .C2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n767), .A2(new_n782), .A3(KEYINPUT51), .A4(new_n769), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n631), .A2(new_n697), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n574), .A2(new_n616), .A3(new_n625), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT112), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n635), .B1(new_n380), .B2(new_n379), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n647), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n665), .A2(new_n788), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n787), .B1(new_n656), .B2(new_n664), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .A3(new_n792), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n572), .A2(new_n671), .A3(new_n675), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n589), .A2(new_n290), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n242), .A2(new_n291), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n387), .A3(new_n591), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n618), .B1(new_n580), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n694), .A2(new_n680), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n696), .A2(new_n651), .ZN(new_n806));
  INV_X1    g620(.A(new_n608), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n242), .A3(new_n627), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n575), .A2(new_n707), .A3(new_n616), .A4(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n806), .A2(new_n715), .B1(new_n663), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n799), .A2(new_n805), .A3(new_n724), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n721), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n798), .A2(new_n812), .A3(KEYINPUT53), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT53), .B1(new_n798), .B2(new_n812), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n796), .B2(new_n792), .ZN(new_n817));
  AND4_X1   g631(.A1(KEYINPUT52), .A2(new_n665), .A3(new_n788), .A4(new_n792), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n720), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n663), .A2(new_n501), .A3(new_n651), .A4(new_n715), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT108), .B1(new_n821), .B2(new_n709), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n713), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n799), .A2(new_n805), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n810), .A2(new_n724), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n816), .B1(new_n819), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n798), .A2(new_n812), .A3(KEYINPUT53), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n780), .A2(new_n833), .A3(new_n784), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n786), .A2(new_n815), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(G952), .B2(G953), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n735), .A2(new_n386), .A3(new_n726), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT49), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n689), .B(new_n837), .C1(new_n838), .C2(new_n683), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT111), .Z(new_n840));
  AOI21_X1  g654(.A(new_n633), .B1(new_n838), .B2(new_n683), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n648), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(G75));
  NOR2_X1   g657(.A1(new_n293), .A2(G952), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n829), .A2(new_n831), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(G902), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT56), .B1(new_n848), .B2(G210), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n371), .A2(new_n374), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n372), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT55), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n845), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n849), .B2(new_n853), .ZN(G51));
  NAND3_X1  g669(.A1(new_n815), .A2(KEYINPUT118), .A3(new_n832), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n857), .A3(KEYINPUT54), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n454), .B(KEYINPUT57), .Z(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(new_n858), .A3(KEYINPUT119), .A4(new_n859), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n451), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n730), .B(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n848), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n844), .B1(new_n864), .B2(new_n866), .ZN(G54));
  NOR2_X1   g681(.A1(new_n279), .A2(new_n282), .ZN(new_n868));
  NAND2_X1  g682(.A1(KEYINPUT58), .A2(G475), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n847), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n847), .B2(new_n869), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n845), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT121), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n870), .A2(new_n874), .A3(new_n845), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(G60));
  XNOR2_X1  g690(.A(new_n581), .B(KEYINPUT59), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n585), .B2(new_n587), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n856), .A2(new_n858), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n815), .B2(new_n832), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n585), .A2(new_n587), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n845), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT122), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n879), .A4(new_n845), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(G63));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n889));
  NAND2_X1  g703(.A1(G217), .A2(G902), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT60), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n846), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT123), .ZN(new_n893));
  INV_X1    g707(.A(new_n487), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n846), .A2(new_n895), .A3(new_n891), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n845), .ZN(new_n898));
  INV_X1    g712(.A(new_n614), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n893), .B2(new_n896), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n889), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n893), .A2(new_n896), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n614), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT61), .A3(new_n845), .A4(new_n897), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(G66));
  NOR3_X1   g719(.A1(new_n298), .A2(new_n343), .A3(new_n293), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n825), .B2(new_n293), .ZN(new_n907));
  INV_X1    g721(.A(G898), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n850), .B1(new_n908), .B2(G953), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n907), .B(new_n909), .Z(G69));
  OR2_X1    g724(.A1(new_n546), .A2(new_n547), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n280), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n665), .A2(new_n788), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(new_n649), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT62), .ZN(new_n916));
  OR3_X1    g730(.A1(new_n914), .A2(KEYINPUT62), .A3(new_n649), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n640), .A2(new_n801), .A3(new_n706), .A4(new_n800), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n663), .A3(new_n501), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT124), .B1(new_n744), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n744), .A2(KEYINPUT124), .A3(new_n919), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n921), .A2(new_n922), .B1(new_n771), .B2(new_n746), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n913), .B1(new_n924), .B2(new_n293), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n912), .B1(G900), .B2(G953), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n705), .A2(new_n639), .A3(new_n734), .A4(new_n791), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n750), .A2(new_n928), .A3(new_n724), .A4(new_n744), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n929), .A2(new_n721), .A3(new_n914), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n930), .B2(new_n293), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT125), .B1(new_n925), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n293), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n926), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n935));
  INV_X1    g749(.A(new_n922), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n750), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n915), .B2(KEYINPUT62), .ZN(new_n938));
  AOI21_X1  g752(.A(G953), .B1(new_n938), .B2(new_n917), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n934), .B(new_n935), .C1(new_n939), .C2(new_n913), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n932), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n932), .B2(new_n940), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n293), .B1(G227), .B2(G900), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n932), .A2(new_n940), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n949), .B2(new_n942), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n947), .A2(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n550), .A2(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n846), .A2(new_n643), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n938), .A2(new_n825), .A3(new_n917), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n643), .B1(new_n957), .B2(new_n953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n954), .B1(new_n930), .B2(new_n825), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n550), .B(KEYINPUT127), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n845), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(G57));
endmodule


