//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n203), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT66), .B(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n203), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n214), .B1(new_n217), .B2(new_n219), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT69), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n250), .A2(new_n252), .A3(new_n254), .A4(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n222), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n250), .A2(new_n252), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n258), .A2(G222), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G1698), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n263), .B(KEYINPUT70), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n215), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n267), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G274), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(G226), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(G190), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n215), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n208), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(G50), .B2(new_n284), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n205), .A2(G20), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n209), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n293), .B1(G150), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n215), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n271), .A2(new_n282), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n283), .B1(new_n301), .B2(new_n302), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT75), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n301), .B2(new_n302), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n296), .A2(new_n297), .ZN(new_n311));
  INV_X1    g0111(.A(new_n289), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(new_n300), .A3(KEYINPUT73), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n303), .A2(G200), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n317), .A2(new_n283), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n308), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n310), .A2(new_n315), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n283), .B(new_n319), .C1(new_n304), .C2(new_n305), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT75), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n307), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n298), .B1(new_n303), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(G179), .B2(new_n303), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n294), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n330), .A2(new_n201), .B1(new_n209), .B2(G68), .ZN(new_n331));
  INV_X1    g0131(.A(G77), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n292), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n297), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT11), .Z(new_n335));
  OAI22_X1  g0135(.A1(new_n284), .A2(G68), .B1(KEYINPUT77), .B2(KEYINPUT12), .ZN(new_n336));
  NAND2_X1  g0136(.A1(KEYINPUT77), .A2(KEYINPUT12), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n286), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G68), .A3(new_n287), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n254), .A2(new_n256), .A3(G226), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n234), .A2(new_n253), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n260), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT76), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT76), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT69), .B(G1698), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n346), .B1(new_n353), .B2(G226), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n352), .B(new_n349), .C1(new_n354), .C2(new_n260), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n351), .A2(new_n355), .A3(new_n270), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n279), .B1(G238), .B2(new_n281), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n357), .B1(new_n356), .B2(new_n358), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n344), .B(G169), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n356), .A2(new_n358), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G179), .A3(new_n359), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n359), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n344), .B1(new_n367), .B2(G169), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n343), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(G200), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n342), .C1(new_n371), .C2(new_n367), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(KEYINPUT78), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n262), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n203), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G159), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n381), .A2(G20), .A3(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G58), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT80), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT80), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(G58), .A3(G68), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n386), .A3(new_n218), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n387), .B2(G20), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n376), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n376), .B(new_n382), .C1(new_n387), .C2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n249), .A2(KEYINPUT79), .A3(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n252), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT79), .B1(new_n249), .B2(G33), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n377), .B(new_n209), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G68), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(new_n252), .A3(new_n392), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n377), .B1(new_n399), .B2(new_n209), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n391), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n390), .A2(new_n401), .A3(new_n297), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n291), .B1(new_n208), .B2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(new_n284), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n403), .A2(new_n339), .B1(new_n404), .B2(new_n291), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n254), .A2(new_n256), .A3(G223), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G226), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n398), .A2(new_n252), .A3(new_n392), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n269), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n275), .A2(G232), .A3(new_n276), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n278), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n326), .B2(new_n419), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n408), .A2(new_n409), .A3(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n423), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n408), .A2(new_n409), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n278), .A2(new_n417), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n412), .A2(new_n413), .B1(G33), .B2(G87), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(G190), .C1(new_n269), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n416), .B2(new_n418), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n402), .A2(new_n405), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT17), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n431), .A2(new_n430), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(KEYINPUT83), .A3(new_n402), .A4(new_n405), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT83), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n439), .B2(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n222), .A2(new_n404), .ZN(new_n441));
  XOR2_X1   g0241(.A(new_n441), .B(KEYINPUT72), .Z(new_n442));
  NAND3_X1  g0242(.A1(new_n339), .A2(G77), .A3(new_n287), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n291), .B(KEYINPUT71), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n330), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n209), .A2(new_n222), .B1(new_n447), .B2(new_n292), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n444), .B1(new_n450), .B2(new_n297), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n258), .A2(G232), .B1(G107), .B2(new_n260), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n264), .B2(new_n221), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n270), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n279), .B1(G244), .B2(new_n281), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n451), .B1(new_n326), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G179), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(G190), .A3(new_n455), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n451), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n427), .A2(new_n440), .A3(new_n460), .A4(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n329), .A2(new_n375), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n374), .A2(KEYINPUT78), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n208), .A2(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G274), .A3(new_n275), .ZN(new_n474));
  INV_X1    g0274(.A(new_n472), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n208), .B(G45), .C1(new_n475), .C2(new_n470), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n275), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n398), .A2(new_n392), .A3(G244), .A4(new_n252), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n254), .A2(new_n256), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n480), .A2(new_n223), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT85), .B1(new_n257), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n353), .A2(new_n262), .A3(new_n490), .A4(new_n484), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n486), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n479), .B1(new_n492), .B2(new_n270), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n458), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n495), .A2(new_n496), .A3(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(G97), .B(G107), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n499), .A2(new_n209), .B1(new_n332), .B2(new_n330), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n378), .B2(new_n379), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n297), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n404), .A2(new_n496), .ZN(new_n504));
  OR3_X1    g0304(.A1(new_n251), .A2(KEYINPUT84), .A3(G1), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT84), .B1(new_n251), .B2(G1), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n286), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n494), .B(new_n510), .C1(G169), .C2(new_n493), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n492), .A2(new_n270), .ZN(new_n512));
  INV_X1    g0312(.A(new_n479), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(G190), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n504), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n498), .A2(new_n495), .ZN(new_n516));
  INV_X1    g0316(.A(new_n497), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n378), .A2(new_n379), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n515), .B1(new_n522), .B2(new_n297), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n514), .B(new_n523), .C1(new_n305), .C2(new_n493), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n209), .A2(G87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n260), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n209), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n501), .A2(KEYINPUT23), .A3(G20), .ZN(new_n530));
  INV_X1    g0330(.A(G116), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n251), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n529), .A2(new_n530), .B1(new_n532), .B2(new_n209), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n398), .A2(new_n392), .A3(new_n209), .A4(new_n252), .ZN(new_n535));
  NAND2_X1  g0335(.A1(KEYINPUT22), .A2(G87), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT24), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT24), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n297), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n476), .A2(new_n275), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G264), .ZN(new_n543));
  INV_X1    g0343(.A(G250), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n482), .A2(new_n544), .B1(new_n478), .B2(new_n253), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n413), .B1(G33), .B2(G294), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n543), .B(new_n474), .C1(new_n546), .C2(new_n269), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT25), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n284), .B2(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n404), .A2(KEYINPUT25), .A3(new_n501), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n508), .A2(G107), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n353), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G294), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n553), .A2(new_n399), .B1(new_n251), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n270), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(G190), .A3(new_n474), .A4(new_n543), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n541), .A2(new_n548), .A3(new_n552), .A4(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n511), .A2(new_n524), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n482), .A2(new_n221), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n532), .B1(new_n560), .B2(new_n413), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT86), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n413), .A2(new_n562), .A3(G244), .A4(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT86), .B1(new_n481), .B2(new_n253), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n270), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n469), .A2(G274), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n469), .A2(new_n544), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n275), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(G190), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  INV_X1    g0371(.A(G87), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(new_n496), .A3(new_n501), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n349), .A2(new_n209), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n571), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n292), .A2(KEYINPUT19), .A3(new_n496), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(new_n535), .B2(new_n203), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n297), .B1(new_n404), .B2(new_n447), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n508), .A2(G87), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n570), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n569), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n565), .B2(new_n270), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n305), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n339), .A2(new_n505), .A3(new_n506), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n578), .B1(new_n447), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n583), .B2(G169), .ZN(new_n587));
  AOI211_X1 g0387(.A(G179), .B(new_n582), .C1(new_n565), .C2(new_n270), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n581), .A2(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n559), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n284), .A2(G116), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n508), .B2(G116), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n488), .B(new_n209), .C1(G33), .C2(new_n496), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n531), .A2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n297), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n326), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT87), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n254), .A2(new_n256), .A3(G257), .ZN(new_n600));
  NAND2_X1  g0400(.A1(G264), .A2(G1698), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n413), .ZN(new_n603));
  INV_X1    g0403(.A(G303), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n262), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n269), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n476), .A2(G270), .A3(new_n275), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n474), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n599), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n399), .B1(new_n601), .B2(new_n600), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n270), .B1(new_n611), .B2(new_n605), .ZN(new_n612));
  INV_X1    g0412(.A(new_n609), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n598), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n607), .A2(new_n609), .A3(new_n458), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n592), .A2(new_n597), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n610), .A2(new_n598), .A3(new_n614), .A4(KEYINPUT21), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n610), .A2(new_n614), .A3(G200), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n371), .B1(new_n610), .B2(new_n614), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n619), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n547), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n458), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n547), .A2(new_n326), .ZN(new_n629));
  INV_X1    g0429(.A(new_n541), .ZN(new_n630));
  INV_X1    g0430(.A(new_n552), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n590), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n468), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT88), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n512), .A2(new_n513), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n326), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n637), .A2(new_n494), .A3(new_n510), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n570), .B(new_n580), .C1(new_n305), .C2(new_n583), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n583), .A2(new_n458), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n640), .B(new_n586), .C1(G169), .C2(new_n583), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g0442(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n632), .A2(new_n617), .A3(new_n620), .A4(new_n621), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n590), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n646), .A3(new_n641), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n468), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n421), .A2(new_n406), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT18), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT18), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n421), .A2(new_n652), .A3(new_n406), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n369), .A2(new_n460), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n440), .A2(new_n372), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n325), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n328), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT90), .ZN(G369));
  NAND3_X1  g0462(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n619), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n626), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n622), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n668), .B1(new_n630), .B2(new_n631), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n558), .A3(new_n632), .ZN(new_n676));
  INV_X1    g0476(.A(new_n668), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n676), .B1(new_n632), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n622), .A2(new_n677), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n632), .A2(new_n668), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n679), .A2(new_n683), .ZN(G399));
  INV_X1    g0484(.A(new_n212), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(G41), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n573), .A2(G116), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G1), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n219), .B2(new_n687), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT28), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n648), .A2(new_n677), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  INV_X1    g0493(.A(new_n589), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(new_n638), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n642), .A2(new_n643), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n641), .B(KEYINPUT92), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT93), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n646), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n677), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n693), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  INV_X1    g0505(.A(G330), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n627), .A2(new_n493), .A3(G179), .ZN(new_n707));
  INV_X1    g0507(.A(new_n583), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n610), .A2(new_n614), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n555), .A2(new_n270), .B1(G264), .B2(new_n542), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n618), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(KEYINPUT30), .A3(new_n583), .A4(new_n493), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n583), .A2(new_n618), .A3(new_n493), .A4(new_n711), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n668), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n633), .A2(new_n677), .B1(new_n720), .B2(KEYINPUT91), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT91), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n706), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n705), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n691), .B1(new_n729), .B2(G1), .ZN(G364));
  XOR2_X1   g0530(.A(new_n673), .B(KEYINPUT94), .Z(new_n731));
  AND2_X1   g0531(.A1(new_n209), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n208), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n686), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n731), .B(new_n736), .C1(G330), .C2(new_n672), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n212), .A2(new_n262), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n739), .B1(G116), .B2(new_n212), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n685), .A2(new_n413), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n219), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n244), .A2(new_n743), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n215), .B1(G20), .B2(new_n326), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n735), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(G190), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G179), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G159), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g0562(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n209), .B1(new_n757), .B2(G190), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n765), .A2(new_n203), .B1(new_n766), .B2(new_n496), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n763), .A2(new_n371), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G50), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n305), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n756), .A2(new_n758), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n209), .A2(new_n371), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n458), .A2(G200), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n260), .B1(new_n777), .B2(G58), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n770), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n755), .A2(new_n775), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n780), .A2(G87), .B1(new_n782), .B2(new_n259), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n769), .A2(new_n773), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G317), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT33), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT33), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n764), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(G326), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n554), .C2(new_n766), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n760), .A2(G329), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n772), .A2(G283), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G322), .A2(new_n777), .B1(new_n782), .B2(G311), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n262), .B1(new_n780), .B2(G303), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n762), .A2(new_n784), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n754), .B1(new_n796), .B2(new_n751), .ZN(new_n797));
  INV_X1    g0597(.A(new_n750), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n672), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n737), .A2(new_n800), .ZN(G396));
  AND2_X1   g0601(.A1(new_n648), .A2(new_n677), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n451), .A2(new_n677), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n463), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n460), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n457), .A2(new_n459), .A3(new_n677), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n802), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n463), .A2(new_n803), .B1(new_n457), .B2(new_n459), .ZN(new_n810));
  INV_X1    g0610(.A(new_n806), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT99), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT99), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n805), .A2(new_n813), .A3(new_n806), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n809), .B1(new_n802), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n735), .B1(new_n816), .B2(new_n727), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n727), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n771), .A2(new_n572), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G311), .B2(new_n760), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n260), .B1(new_n779), .B2(new_n501), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n776), .A2(new_n554), .B1(new_n781), .B2(new_n531), .ZN(new_n823));
  INV_X1    g0623(.A(new_n766), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(G97), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT97), .B(G283), .Z(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(new_n764), .B1(new_n768), .B2(G303), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n820), .A2(new_n822), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n777), .B1(new_n782), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(new_n768), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n830), .B1(new_n831), .B2(new_n832), .C1(new_n833), .C2(new_n765), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n413), .B1(new_n201), .B2(new_n779), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G58), .B2(new_n824), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n760), .A2(G132), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n772), .A2(G68), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n834), .A2(new_n835), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n829), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n751), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n751), .A2(new_n748), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n736), .B1(new_n332), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(new_n808), .C2(new_n749), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n818), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  AND2_X1   g0649(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n850), .A2(new_n851), .A3(new_n531), .A4(new_n217), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  OR3_X1    g0653(.A1(new_n387), .A2(new_n201), .A3(new_n222), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n201), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n208), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n343), .A2(new_n668), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT101), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n373), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n858), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n369), .A3(new_n372), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n807), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n590), .A2(new_n626), .A3(new_n632), .A4(new_n677), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n720), .A3(new_n722), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT104), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n396), .A2(new_n400), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT16), .B1(new_n868), .B2(new_n388), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n401), .A2(new_n297), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n405), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n666), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n421), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n438), .A3(new_n436), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n408), .B(new_n409), .C1(new_n421), .C2(new_n872), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n438), .A4(new_n436), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n427), .A2(new_n440), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n871), .A2(new_n872), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT102), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n884), .B(new_n881), .C1(new_n427), .C2(new_n440), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n879), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n875), .B2(new_n878), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n883), .B2(new_n885), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n867), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n866), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT40), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n655), .A2(new_n440), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n408), .A2(new_n409), .A3(new_n872), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n650), .A2(new_n432), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n895), .A2(new_n896), .B1(new_n878), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n890), .B1(KEYINPUT38), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n864), .A2(KEYINPUT40), .A3(new_n866), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n894), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n866), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n467), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n903), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n906), .A2(new_n907), .A3(new_n706), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n888), .A2(new_n890), .ZN(new_n909));
  INV_X1    g0709(.A(new_n889), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n880), .A2(new_n882), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n884), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n880), .A2(KEYINPUT102), .A3(new_n882), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT103), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n898), .A2(new_n878), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n433), .B1(new_n436), .B2(new_n438), .ZN(new_n919));
  NOR3_X1   g0719(.A1(new_n654), .A2(new_n919), .A3(new_n434), .ZN(new_n920));
  INV_X1    g0720(.A(new_n896), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT39), .B1(new_n922), .B2(new_n887), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT103), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n890), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(KEYINPUT39), .A2(new_n909), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n369), .A2(new_n668), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n806), .B(KEYINPUT100), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n809), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n860), .A2(new_n863), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n912), .A2(new_n913), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n887), .A2(new_n886), .B1(new_n933), .B2(new_n889), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n932), .A2(new_n934), .B1(new_n655), .B2(new_n872), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n928), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n660), .B1(new_n705), .B2(new_n467), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OAI22_X1  g0738(.A1(new_n908), .A2(new_n938), .B1(new_n208), .B2(new_n732), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n908), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n857), .B1(new_n939), .B2(new_n940), .ZN(G367));
  OAI211_X1 g0741(.A(new_n511), .B(new_n524), .C1(new_n523), .C2(new_n677), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n638), .A2(new_n668), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n681), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT106), .Z(new_n947));
  OR2_X1    g0747(.A1(new_n942), .A2(new_n632), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n668), .B1(new_n948), .B2(new_n511), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n945), .B2(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT43), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n580), .A2(new_n677), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT105), .Z(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n694), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n641), .B2(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n954), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n958), .B2(new_n954), .ZN(new_n960));
  INV_X1    g0760(.A(new_n679), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n944), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n959), .B(new_n964), .C1(new_n958), .C2(new_n954), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n686), .B(KEYINPUT41), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n678), .B1(new_n622), .B2(new_n677), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n967), .A2(KEYINPUT109), .A3(new_n681), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(KEYINPUT109), .B2(new_n681), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n731), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n673), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n728), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n683), .A2(new_n944), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n683), .A2(new_n944), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n973), .B1(new_n978), .B2(new_n961), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n961), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n978), .A2(new_n973), .A3(new_n961), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n972), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n966), .B1(new_n983), .B2(new_n729), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n963), .B(new_n965), .C1(new_n984), .C2(new_n734), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n741), .A2(new_n240), .ZN(new_n986));
  INV_X1    g0786(.A(new_n447), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n753), .B1(new_n685), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n736), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n751), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n776), .A2(new_n833), .B1(new_n781), .B2(new_n201), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n260), .B(new_n991), .C1(G58), .C2(new_n780), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n765), .A2(new_n381), .B1(new_n766), .B2(new_n203), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G143), .B2(new_n768), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n760), .A2(G137), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n772), .A2(new_n259), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(KEYINPUT110), .B(G317), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G97), .A2(new_n772), .B1(new_n760), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n780), .A2(G116), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT46), .ZN(new_n1001));
  INV_X1    g0801(.A(G311), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n831), .A2(new_n1002), .B1(new_n766), .B2(new_n501), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G294), .B2(new_n764), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n826), .A2(new_n781), .B1(new_n776), .B2(new_n604), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n413), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n999), .A2(new_n1001), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n997), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT47), .Z(new_n1009));
  OAI221_X1 g0809(.A(new_n989), .B1(new_n990), .B2(new_n1009), .C1(new_n958), .C2(new_n798), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  NOR2_X1   g0811(.A1(new_n972), .A2(new_n687), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n971), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1012), .B1(new_n729), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n678), .A2(new_n798), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n738), .A2(new_n688), .B1(G107), .B2(new_n212), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n445), .A2(G50), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT50), .ZN(new_n1018));
  AOI21_X1  g0818(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n688), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n742), .B1(new_n237), .B2(G45), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1016), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n735), .B1(new_n1022), .B2(new_n753), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n781), .A2(new_n203), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n779), .A2(new_n222), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G50), .C2(new_n777), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n496), .B2(new_n771), .C1(new_n833), .C2(new_n759), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n766), .A2(new_n447), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n381), .A2(new_n831), .B1(new_n765), .B2(new_n291), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1027), .A2(new_n399), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT111), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n777), .A2(new_n998), .B1(new_n782), .B2(G303), .ZN(new_n1032));
  INV_X1    g0832(.A(G322), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1032), .B1(new_n831), .B2(new_n1033), .C1(new_n1002), .C2(new_n765), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n826), .A2(new_n766), .B1(new_n779), .B2(new_n554), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n413), .B1(new_n760), .B2(G326), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n531), .C2(new_n771), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT49), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1031), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1023), .B1(new_n1043), .B2(new_n751), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1013), .A2(new_n734), .B1(new_n1015), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1014), .A2(new_n1045), .ZN(G393));
  XNOR2_X1  g0846(.A(new_n978), .B(new_n679), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n983), .B(new_n686), .C1(new_n972), .C2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n942), .A2(new_n943), .A3(new_n750), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n752), .B1(new_n496), .B2(new_n212), .C1(new_n742), .C2(new_n247), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n735), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n760), .A2(G143), .B1(G68), .B2(new_n780), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT112), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n766), .A2(new_n332), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n764), .B2(G50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n445), .B2(new_n781), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT113), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n831), .A2(new_n833), .B1(new_n776), .B2(new_n381), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT51), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1060), .A2(new_n1061), .A3(new_n819), .A4(new_n399), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1053), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n262), .B1(new_n827), .B2(new_n780), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n773), .B(new_n1064), .C1(new_n1033), .C2(new_n759), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT114), .Z(new_n1066));
  OAI22_X1  g0866(.A1(new_n831), .A2(new_n785), .B1(new_n776), .B2(new_n1002), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT52), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n781), .A2(new_n554), .B1(new_n766), .B2(new_n531), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G303), .B2(new_n764), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1063), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT115), .Z(new_n1073));
  AOI21_X1  g0873(.A(new_n1051), .B1(new_n1073), .B2(new_n751), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1047), .A2(new_n734), .B1(new_n1049), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1048), .A2(KEYINPUT116), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(KEYINPUT116), .B1(new_n1048), .B2(new_n1075), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(G390));
  AOI22_X1  g0880(.A1(new_n699), .A2(KEYINPUT93), .B1(new_n590), .B2(new_n645), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n668), .B1(new_n1081), .B2(new_n702), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n811), .B1(new_n1082), .B2(new_n805), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n931), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n927), .B(new_n900), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n726), .A2(new_n864), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n890), .A2(new_n924), .A3(new_n923), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n924), .B1(new_n890), .B2(new_n923), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n915), .A2(new_n934), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n927), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n930), .B2(new_n931), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1085), .B(new_n1086), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n899), .A2(KEYINPUT38), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n927), .B1(new_n914), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n806), .B1(new_n704), .B2(new_n810), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n931), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n932), .A2(new_n927), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n926), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n904), .A2(new_n706), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n864), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1092), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n733), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n926), .A2(new_n748), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n845), .A2(new_n291), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n776), .A2(new_n531), .B1(new_n781), .B2(new_n496), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n262), .B(new_n1105), .C1(G87), .C2(new_n780), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n840), .C1(new_n554), .C2(new_n759), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1054), .B1(new_n764), .B2(G107), .ZN(new_n1108));
  INV_X1    g0908(.A(G283), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n831), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n824), .A2(G159), .B1(G128), .B2(new_n768), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT53), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n779), .A2(new_n833), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G50), .A2(new_n772), .B1(new_n760), .B2(G125), .ZN(new_n1115));
  INV_X1    g0915(.A(G132), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n262), .B1(new_n776), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n782), .B2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1113), .A2(new_n1112), .B1(G137), .B2(new_n764), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1115), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1107), .A2(new_n1110), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n736), .B(new_n1104), .C1(new_n1123), .C2(new_n751), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1102), .B1(new_n1103), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n720), .A2(KEYINPUT91), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n865), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT91), .B1(new_n720), .B2(new_n722), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n808), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1084), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1100), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n815), .A2(new_n866), .A3(G330), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n726), .A2(new_n864), .B1(new_n1084), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1131), .A2(new_n930), .B1(new_n1133), .B2(new_n1083), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n465), .A2(new_n466), .A3(new_n1099), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n660), .B(new_n1135), .C1(new_n705), .C2(new_n467), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1101), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1092), .B(new_n1137), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n686), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1125), .A2(new_n1141), .ZN(G378));
  INV_X1    g0942(.A(KEYINPUT119), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n706), .B1(new_n900), .B2(new_n902), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n894), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n934), .A2(new_n892), .A3(new_n867), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1144), .B(KEYINPUT119), .C1(new_n1147), .C2(KEYINPUT40), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n298), .A2(new_n666), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n329), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n329), .A2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1146), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1154), .B(new_n1143), .C1(new_n894), .C2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n936), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1156), .A2(new_n936), .A3(new_n1157), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1155), .A2(new_n748), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n771), .A2(new_n202), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n776), .A2(new_n501), .B1(new_n781), .B2(new_n447), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1164), .A2(new_n1165), .A3(G41), .A4(new_n1025), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n765), .A2(new_n496), .B1(new_n831), .B2(new_n531), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n413), .B(new_n1167), .C1(G68), .C2(new_n824), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n1109), .C2(new_n759), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT58), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n413), .B2(G33), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G128), .A2(new_n777), .B1(new_n780), .B2(new_n1119), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n782), .A2(G137), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n768), .A2(G125), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n824), .A2(G150), .B1(G132), .B2(new_n764), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n760), .A2(G124), .ZN(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n772), .C2(G159), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1170), .B1(G50), .B2(new_n1171), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT117), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n751), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT118), .Z(new_n1185));
  AOI211_X1 g0985(.A(new_n736), .B(new_n1185), .C1(new_n201), .C2(new_n845), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1162), .A2(new_n734), .B1(new_n1163), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1136), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1188), .B1(new_n1140), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1160), .A2(new_n1190), .A3(new_n1161), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(KEYINPUT120), .A3(new_n686), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1140), .A2(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1160), .A2(new_n1161), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1188), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT120), .B1(new_n1191), .B2(new_n686), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1187), .B1(new_n1196), .B2(new_n1197), .ZN(G375));
  AOI21_X1  g0998(.A(new_n736), .B1(new_n203), .B2(new_n845), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1164), .A2(new_n399), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT123), .Z(new_n1201));
  OAI22_X1  g1001(.A1(new_n831), .A2(new_n1116), .B1(new_n766), .B2(new_n201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n780), .A2(G159), .B1(new_n782), .B2(G150), .ZN(new_n1203));
  INV_X1    g1003(.A(G128), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1203), .B1(new_n1204), .B2(new_n759), .C1(new_n832), .C2(new_n776), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(new_n764), .C2(new_n1119), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n765), .A2(new_n531), .B1(new_n447), .B2(new_n766), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n780), .A2(G97), .B1(new_n782), .B2(G107), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n1109), .B2(new_n776), .C1(new_n604), .C2(new_n759), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(G294), .C2(new_n768), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n260), .B1(new_n771), .B2(new_n332), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  AOI22_X1  g1012(.A1(new_n1201), .A2(new_n1206), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1199), .B1(new_n1213), .B2(new_n990), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1084), .B2(new_n748), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1134), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n734), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n966), .B(KEYINPUT121), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1138), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1216), .A2(new_n1189), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(G381));
  INV_X1    g1021(.A(G375), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1125), .A2(new_n1224), .A3(new_n1141), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1222), .A2(new_n1227), .A3(new_n1228), .A4(new_n1230), .ZN(G407));
  NAND2_X1  g1031(.A1(new_n667), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1222), .A2(new_n1227), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(G407), .A2(G213), .A3(new_n1234), .ZN(G409));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1162), .A2(new_n1193), .A3(new_n1218), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1187), .A2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G378), .B(new_n1187), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1220), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n686), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1242), .A2(new_n1220), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1217), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n848), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1246), .A2(new_n848), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G2897), .B(new_n1233), .C1(new_n1248), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1249), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1233), .A2(G2897), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1247), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1236), .B1(new_n1241), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1232), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1079), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G390), .A2(new_n1010), .A3(new_n985), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G393), .B(G396), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1263), .B2(KEYINPUT126), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1265), .B(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1260), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1256), .A2(new_n1262), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1259), .A2(KEYINPUT62), .A3(new_n1261), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1241), .B2(new_n1260), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1272), .A2(new_n1255), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1271), .B1(new_n1275), .B2(new_n1269), .ZN(G405));
  NAND2_X1  g1076(.A1(G375), .A2(new_n1227), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n1240), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1277), .B2(new_n1240), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1260), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1268), .B(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1240), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1191), .A2(new_n686), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT120), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1287), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1226), .B1(new_n1288), .B2(new_n1187), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT127), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1277), .A2(new_n1278), .A3(new_n1240), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1261), .A3(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1281), .A2(new_n1283), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1283), .B1(new_n1281), .B2(new_n1292), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G402));
endmodule


