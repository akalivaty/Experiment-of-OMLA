//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n214), .A2(G50), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G20), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G116), .A2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G238), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n202), .C2(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n226), .B(new_n231), .C1(G97), .C2(G257), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n208), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT1), .Z(new_n234));
  AOI211_X1 g0034(.A(new_n220), .B(new_n234), .C1(new_n213), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n247), .B(KEYINPUT67), .Z(new_n248));
  XOR2_X1   g0048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT66), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G50), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n255), .A2(KEYINPUT72), .B1(G20), .B2(new_n202), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n207), .A2(G33), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n256), .B1(KEYINPUT72), .B2(new_n255), .C1(new_n222), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n217), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n206), .B2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n261), .B1(new_n202), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT11), .B1(new_n258), .B2(new_n260), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G68), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT12), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n229), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G232), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(KEYINPUT70), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT70), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n283), .B(new_n280), .C1(new_n275), .C2(new_n276), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n280), .A2(G238), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n285), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G274), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT71), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n282), .A2(new_n284), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT13), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT13), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n293), .B1(new_n289), .B2(new_n290), .C1(new_n282), .C2(new_n284), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n269), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(new_n292), .B2(new_n294), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n292), .A2(new_n294), .A3(G179), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT14), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n295), .A2(new_n304), .A3(G169), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n269), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n309));
  INV_X1    g0109(.A(G150), .ZN(new_n310));
  INV_X1    g0110(.A(new_n254), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT8), .B(G58), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n309), .B1(new_n310), .B2(new_n311), .C1(new_n312), .C2(new_n257), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n260), .ZN(new_n314));
  INV_X1    g0114(.A(new_n266), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n228), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n262), .A2(G50), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT69), .B(G200), .Z(new_n319));
  NOR2_X1   g0119(.A1(new_n281), .A2(new_n287), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G226), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G223), .A2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n271), .A2(G222), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n270), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n281), .C1(G77), .C2(new_n270), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n325), .A3(new_n288), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n318), .A2(KEYINPUT9), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n327), .B1(KEYINPUT9), .B2(new_n318), .C1(new_n296), .C2(new_n326), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT10), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n318), .B1(new_n330), .B2(new_n326), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT68), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G179), .B2(new_n326), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G238), .A2(G1698), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n270), .B(new_n334), .C1(new_n273), .C2(G1698), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n335), .B(new_n281), .C1(G107), .C2(new_n270), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n320), .A2(G244), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n288), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G20), .A2(G77), .ZN(new_n340));
  XOR2_X1   g0140(.A(KEYINPUT15), .B(G87), .Z(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n340), .B1(new_n311), .B2(new_n312), .C1(new_n342), .C2(new_n257), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n260), .B1(new_n222), .B2(new_n315), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n262), .A2(G77), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(new_n330), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n339), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n308), .A2(new_n329), .A3(new_n333), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n312), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n315), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(new_n263), .B2(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(new_n260), .ZN(new_n353));
  XNOR2_X1  g0153(.A(G58), .B(G68), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(G20), .B1(G159), .B2(new_n254), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G33), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n360), .B2(new_n207), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  AOI211_X1 g0162(.A(new_n362), .B(G20), .C1(new_n357), .C2(new_n359), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n362), .B1(new_n270), .B2(G20), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT73), .A3(G68), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n356), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n353), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT74), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n361), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n374), .A2(G68), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(new_n356), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n352), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n320), .A2(G232), .B1(G274), .B2(new_n287), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n357), .A2(new_n359), .A3(G226), .A4(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n270), .A2(new_n385), .A3(G226), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n270), .A2(G223), .A3(new_n271), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n384), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n281), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(new_n392), .A3(new_n281), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n382), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(G169), .B1(new_n390), .B2(new_n380), .ZN(new_n395));
  OR2_X1    g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT18), .B1(new_n379), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT73), .B1(new_n369), .B2(G68), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n365), .B(new_n202), .C1(new_n367), .C2(new_n368), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT16), .B(new_n355), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n378), .A2(new_n400), .A3(new_n260), .ZN(new_n401));
  INV_X1    g0201(.A(new_n352), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n394), .A2(new_n395), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT18), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n380), .A2(new_n296), .ZN(new_n407));
  INV_X1    g0207(.A(new_n393), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n392), .B1(new_n389), .B2(new_n281), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n390), .A2(new_n380), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n298), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n401), .A3(new_n402), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n413), .A2(new_n401), .A3(KEYINPUT17), .A4(new_n402), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n397), .A2(new_n406), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n338), .A2(new_n296), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n419), .B(new_n346), .C1(new_n319), .C2(new_n338), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n349), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n374), .A2(new_n376), .A3(G107), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT6), .A3(G97), .ZN(new_n425));
  INV_X1    g0225(.A(G97), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n424), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G97), .A2(G107), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n425), .B1(new_n429), .B2(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n254), .A2(G77), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n423), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n260), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n266), .A2(new_n426), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n206), .A2(G33), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n266), .A2(new_n436), .A3(new_n217), .A4(new_n259), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n435), .B1(new_n438), .B2(new_n426), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT77), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT79), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n434), .A2(new_n443), .A3(new_n440), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n206), .B(G45), .C1(new_n279), .C2(KEYINPUT5), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(G257), .A3(new_n280), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n357), .A2(new_n359), .A3(G244), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n450), .A2(new_n451), .B1(G33), .B2(G283), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n270), .B2(G250), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(new_n453), .C1(new_n271), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n449), .B1(new_n455), .B2(new_n281), .ZN(new_n456));
  INV_X1    g0256(.A(G274), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G179), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n458), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G169), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n442), .A2(new_n444), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n434), .A2(new_n440), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n296), .B1(new_n298), .B2(KEYINPUT78), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(KEYINPUT78), .A3(G200), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n422), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n424), .A3(G20), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n470), .A2(new_n472), .A3(new_n473), .A4(KEYINPUT84), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n357), .A2(new_n359), .A3(new_n207), .A4(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n270), .A2(new_n481), .A3(new_n207), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT83), .B(KEYINPUT24), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n478), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n478), .B2(new_n483), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n260), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n266), .A2(G107), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT25), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n489), .A2(KEYINPUT25), .B1(new_n437), .B2(new_n424), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n280), .B(G264), .C1(new_n445), .C2(new_n446), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n357), .B(new_n359), .C1(G250), .C2(G1698), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n271), .A2(G257), .ZN(new_n497));
  INV_X1    g0297(.A(G294), .ZN(new_n498));
  OAI22_X1  g0298(.A1(new_n496), .A2(new_n497), .B1(new_n278), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n281), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n500), .A3(new_n458), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n330), .ZN(new_n503));
  INV_X1    g0303(.A(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n381), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n493), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(G238), .A2(G1698), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n223), .B2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n270), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n281), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n514));
  INV_X1    g0314(.A(G45), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n280), .B(G250), .C1(G1), .C2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n381), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n509), .A2(new_n270), .B1(G33), .B2(G116), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n514), .B(new_n516), .C1(new_n518), .C2(new_n280), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n330), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n224), .A2(new_n426), .A3(new_n424), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n276), .A2(new_n207), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT19), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n357), .A2(new_n359), .A3(new_n207), .A4(G68), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n257), .A2(new_n426), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n523), .B(new_n524), .C1(KEYINPUT19), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n260), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n438), .A2(new_n341), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n342), .A2(new_n315), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n517), .A2(new_n520), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n438), .A2(G87), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n513), .A2(new_n296), .A3(new_n514), .A4(new_n516), .ZN(new_n534));
  INV_X1    g0334(.A(new_n319), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n519), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT81), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n534), .A2(new_n536), .ZN(new_n539));
  INV_X1    g0339(.A(new_n533), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT81), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n517), .A2(new_n520), .A3(new_n530), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n502), .A2(G200), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n487), .A2(new_n546), .A3(new_n490), .A4(new_n492), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n502), .A2(new_n296), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n507), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G264), .A2(G1698), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n271), .A2(G257), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n270), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n281), .C1(G303), .C2(new_n270), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n447), .A2(G270), .A3(new_n280), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n458), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n438), .A2(G116), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n315), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n259), .A2(new_n217), .B1(G20), .B2(new_n559), .ZN(new_n561));
  AOI21_X1  g0361(.A(G20), .B1(G33), .B2(G283), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G33), .B2(new_n426), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT20), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT20), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n558), .B(new_n560), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n557), .B(new_n567), .C1(new_n296), .C2(new_n556), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(G169), .A3(new_n566), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n458), .A2(new_n554), .A3(G179), .A4(new_n555), .ZN(new_n572));
  OR2_X1    g0372(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n556), .A2(KEYINPUT21), .A3(new_n566), .A4(G169), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n568), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n462), .B1(new_n381), .B2(new_n461), .ZN(new_n578));
  INV_X1    g0378(.A(new_n444), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n443), .B1(new_n434), .B2(new_n440), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(KEYINPUT80), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n469), .A2(new_n550), .A3(new_n577), .A4(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n421), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g0386(.A(new_n586), .B(KEYINPUT86), .Z(G372));
  INV_X1    g0387(.A(new_n333), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n397), .A2(new_n406), .ZN(new_n589));
  INV_X1    g0389(.A(new_n300), .ZN(new_n590));
  INV_X1    g0390(.A(new_n348), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n306), .B2(new_n307), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT88), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n416), .A2(new_n417), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n589), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n588), .B1(new_n596), .B2(new_n329), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n463), .A2(new_n468), .ZN(new_n598));
  INV_X1    g0398(.A(new_n549), .ZN(new_n599));
  XOR2_X1   g0399(.A(new_n533), .B(KEYINPUT87), .Z(new_n600));
  AOI21_X1  g0400(.A(new_n531), .B1(new_n600), .B2(new_n539), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n506), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n598), .A2(new_n599), .A3(new_n601), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n578), .A2(new_n441), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n601), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n463), .A2(new_n544), .A3(new_n538), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT26), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n604), .A2(new_n543), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n421), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(new_n612), .ZN(G369));
  NOR2_X1   g0413(.A1(new_n209), .A2(G20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n206), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(G213), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(G343), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n577), .B1(new_n567), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n602), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n566), .A3(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G330), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT89), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n493), .A2(new_n620), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n507), .B1(new_n599), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n507), .B2(new_n621), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n602), .A2(new_n620), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n634), .A2(new_n636), .B1(new_n507), .B2(new_n621), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(G399));
  NOR2_X1   g0438(.A1(new_n210), .A2(G41), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n521), .A2(G116), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(G1), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n216), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT28), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n572), .B(KEYINPUT90), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(new_n519), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n459), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT30), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n504), .A2(G179), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n651), .A2(new_n461), .A3(new_n556), .A4(new_n519), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n620), .ZN(new_n655));
  OAI211_X1 g0455(.A(KEYINPUT31), .B(new_n655), .C1(new_n584), .C2(new_n620), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(KEYINPUT31), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n658), .A2(G330), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n609), .A2(new_n607), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT91), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n606), .A2(KEYINPUT26), .A3(new_n601), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n609), .A2(new_n663), .A3(new_n607), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n604), .A2(new_n543), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n620), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT29), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n611), .A2(new_n621), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n659), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n644), .B1(new_n672), .B2(G1), .ZN(G364));
  INV_X1    g0473(.A(new_n631), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n614), .B(KEYINPUT92), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n206), .B1(new_n675), .B2(G45), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n639), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n674), .B(new_n679), .C1(G330), .C2(new_n625), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n217), .B1(G20), .B2(new_n330), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n381), .A2(new_n298), .A3(G190), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G20), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n426), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n207), .A2(new_n381), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G200), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G190), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n270), .B1(new_n689), .B2(new_n202), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n207), .A2(G179), .ZN(new_n691));
  NOR2_X1   g0491(.A1(G190), .A2(G200), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G159), .ZN(new_n695));
  AOI211_X1 g0495(.A(new_n685), .B(new_n690), .C1(KEYINPUT32), .C2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n686), .A2(G190), .A3(new_n298), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n695), .A2(KEYINPUT32), .B1(new_n201), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n687), .A2(new_n296), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(G50), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n686), .A2(new_n692), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G77), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n319), .A2(new_n691), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n296), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(G190), .ZN(new_n706));
  AOI22_X1  g0506(.A1(G87), .A2(new_n705), .B1(new_n706), .B2(G107), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n696), .A2(new_n700), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(KEYINPUT33), .B(G317), .Z(new_n709));
  INV_X1    g0509(.A(G322), .ZN(new_n710));
  OAI22_X1  g0510(.A1(new_n689), .A2(new_n709), .B1(new_n697), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT93), .Z(new_n712));
  AOI22_X1  g0512(.A1(G283), .A2(new_n706), .B1(new_n705), .B2(G303), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n699), .A2(G326), .B1(G294), .B2(new_n683), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n270), .B1(new_n694), .B2(G329), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G311), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n701), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n708), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n252), .A2(G45), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n210), .A2(new_n270), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n720), .B(new_n721), .C1(G45), .C2(new_n216), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n210), .A2(new_n360), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G355), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n722), .B(new_n724), .C1(G116), .C2(new_n211), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G13), .A2(G33), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n681), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n681), .A2(new_n719), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n728), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n678), .B(new_n730), .C1(new_n625), .C2(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n680), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(G396));
  OAI21_X1  g0534(.A(new_n270), .B1(new_n684), .B2(new_n201), .ZN(new_n735));
  INV_X1    g0535(.A(new_n706), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n202), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n735), .B(new_n737), .C1(G50), .C2(new_n705), .ZN(new_n738));
  INV_X1    g0538(.A(new_n697), .ZN(new_n739));
  AOI22_X1  g0539(.A1(G150), .A2(new_n688), .B1(new_n739), .B2(G143), .ZN(new_n740));
  INV_X1    g0540(.A(G137), .ZN(new_n741));
  INV_X1    g0541(.A(new_n699), .ZN(new_n742));
  INV_X1    g0542(.A(G159), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n740), .B1(new_n741), .B2(new_n742), .C1(new_n743), .C2(new_n701), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT34), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n694), .A2(G132), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n738), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n688), .A2(G283), .B1(new_n702), .B2(G116), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(KEYINPUT95), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G303), .A2(new_n699), .B1(new_n739), .B2(G294), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n717), .B2(new_n693), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n753), .A2(new_n270), .A3(new_n685), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n750), .A2(KEYINPUT95), .B1(new_n705), .B2(G107), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(new_n755), .C1(new_n224), .C2(new_n736), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n749), .B1(new_n751), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n681), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n681), .A2(new_n726), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n679), .B1(new_n222), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  AOI21_X1  g0561(.A(new_n621), .B1(new_n344), .B2(new_n345), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n348), .B1(new_n420), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n348), .A2(new_n620), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n758), .B(new_n761), .C1(new_n767), .C2(new_n727), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n766), .B(KEYINPUT96), .Z(new_n769));
  MUX2_X1   g0569(.A(new_n766), .B(new_n769), .S(new_n669), .Z(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(new_n659), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n771), .B2(new_n678), .ZN(G384));
  AND3_X1   g0572(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n773), .A2(new_n269), .A3(new_n620), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT101), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT38), .ZN(new_n776));
  INV_X1    g0576(.A(new_n618), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n400), .A2(new_n260), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n366), .A2(new_n370), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT16), .B1(new_n779), .B2(new_n355), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n402), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT98), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(KEYINPUT98), .B(new_n402), .C1(new_n778), .C2(new_n780), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n418), .A2(new_n777), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n618), .B1(new_n394), .B2(new_n395), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n403), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT37), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n788), .A2(new_n789), .A3(new_n414), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n783), .A2(new_n784), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n414), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(new_n792), .B2(KEYINPUT37), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n776), .B1(new_n786), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n418), .A2(new_n777), .A3(new_n785), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n789), .B1(new_n791), .B2(new_n414), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(KEYINPUT38), .C1(new_n796), .C2(new_n790), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n794), .A2(KEYINPUT99), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT99), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n776), .C1(new_n786), .C2(new_n793), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT39), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n418), .A2(new_n403), .A3(new_n777), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n789), .B1(new_n788), .B2(new_n414), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n790), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT38), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT39), .B1(new_n807), .B2(new_n797), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n775), .B1(new_n802), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT39), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n798), .B2(new_n800), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n812), .A2(KEYINPUT101), .A3(new_n808), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n774), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n669), .C2(new_n766), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n307), .A2(new_n620), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n590), .B(new_n818), .C1(new_n773), .C2(new_n269), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n307), .B(new_n620), .C1(new_n306), .C2(new_n300), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n817), .A2(new_n800), .A3(new_n798), .A4(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n589), .A2(new_n777), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(KEYINPUT100), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT100), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n814), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n668), .A2(new_n421), .A3(new_n671), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n597), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n827), .B(new_n829), .Z(new_n830));
  AOI21_X1  g0630(.A(new_n766), .B1(new_n819), .B2(new_n820), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT40), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n656), .A2(new_n831), .A3(new_n832), .A4(new_n657), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT102), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT102), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n656), .A2(new_n831), .A3(new_n835), .A4(new_n657), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n834), .A2(new_n800), .A3(new_n798), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n807), .A2(new_n797), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n656), .A2(new_n657), .A3(new_n831), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT40), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n658), .A2(new_n421), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G330), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n830), .B(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n206), .B2(new_n675), .ZN(new_n847));
  OAI211_X1 g0647(.A(G20), .B(new_n218), .C1(new_n430), .C2(KEYINPUT35), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n559), .B(new_n848), .C1(KEYINPUT35), .C2(new_n430), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  OAI21_X1  g0650(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n216), .A2(new_n851), .B1(G50), .B2(new_n202), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(G1), .A3(new_n209), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n847), .A2(new_n850), .A3(new_n853), .ZN(G367));
  AOI22_X1  g0654(.A1(new_n702), .A2(G283), .B1(G107), .B2(new_n683), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(KEYINPUT106), .ZN(new_n856));
  INV_X1    g0656(.A(new_n705), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n857), .A2(new_n559), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n858), .B2(KEYINPUT46), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT46), .B2(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(G303), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n742), .A2(new_n717), .B1(new_n861), .B2(new_n697), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n270), .B(new_n862), .C1(G317), .C2(new_n694), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n863), .B1(new_n426), .B2(new_n736), .C1(new_n498), .C2(new_n689), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n860), .B(new_n864), .C1(KEYINPUT106), .C2(new_n855), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n699), .A2(G143), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n683), .A2(G68), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n866), .B(new_n867), .C1(new_n310), .C2(new_n697), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT107), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n270), .B1(new_n701), .B2(new_n228), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G159), .B2(new_n688), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n705), .A2(G58), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n706), .A2(G77), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n870), .B(new_n876), .C1(G137), .C2(new_n694), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n865), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT47), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n681), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n600), .A2(new_n621), .ZN(new_n881));
  MUX2_X1   g0681(.A(new_n601), .B(new_n531), .S(new_n881), .Z(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(new_n731), .ZN(new_n883));
  INV_X1    g0683(.A(new_n721), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n729), .B1(new_n211), .B2(new_n342), .C1(new_n243), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n678), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT105), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n598), .B1(new_n464), .B2(new_n621), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n606), .A2(new_n620), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR3_X1    g0691(.A1(new_n637), .A2(KEYINPUT44), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT44), .B1(new_n637), .B2(new_n891), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n637), .A2(KEYINPUT45), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT45), .B1(new_n637), .B2(new_n891), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n631), .A3(new_n634), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n635), .A2(new_n897), .A3(new_n894), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n634), .B(new_n636), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n629), .A2(new_n630), .B1(KEYINPUT103), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(KEYINPUT103), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n674), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n672), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n672), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n639), .B(KEYINPUT41), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n677), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n891), .A2(new_n634), .A3(new_n636), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT42), .Z(new_n912));
  AOI21_X1  g0712(.A(new_n463), .B1(new_n891), .B2(new_n507), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n620), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n891), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n635), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n916), .A2(new_n918), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n922), .B1(new_n920), .B2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT104), .B1(new_n910), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n910), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n888), .B1(new_n928), .B2(new_n929), .ZN(G387));
  XOR2_X1   g0730(.A(new_n639), .B(KEYINPUT111), .Z(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n905), .B2(new_n672), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n672), .B2(new_n905), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n884), .B1(new_n240), .B2(G45), .ZN(new_n934));
  INV_X1    g0734(.A(new_n641), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n935), .B2(new_n723), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n350), .A2(new_n228), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n935), .B1(new_n937), .B2(KEYINPUT50), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n515), .C1(KEYINPUT50), .C2(new_n937), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G68), .B2(G77), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n936), .A2(new_n940), .B1(G107), .B2(new_n211), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n679), .B1(new_n941), .B2(new_n729), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n943));
  INV_X1    g0743(.A(new_n681), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n683), .A2(G283), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G311), .A2(new_n688), .B1(new_n739), .B2(G317), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n861), .B2(new_n701), .C1(new_n710), .C2(new_n742), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT48), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n945), .B1(new_n498), .B2(new_n857), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT110), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(KEYINPUT49), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n694), .A2(G326), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(KEYINPUT49), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n270), .B1(new_n706), .B2(G116), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n954), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n360), .B1(new_n694), .B2(G150), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(new_n202), .B2(new_n701), .C1(new_n742), .C2(new_n743), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n857), .A2(new_n222), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G97), .C2(new_n706), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n341), .A2(new_n683), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n228), .B2(new_n697), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT109), .Z(new_n964));
  OAI211_X1 g0764(.A(new_n961), .B(new_n964), .C1(new_n312), .C2(new_n689), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n944), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n634), .A2(new_n731), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n942), .A2(KEYINPUT108), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n905), .A2(new_n677), .B1(new_n943), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n933), .A2(new_n970), .ZN(G393));
  INV_X1    g0771(.A(new_n931), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n901), .A2(new_n906), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n907), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n899), .A2(new_n900), .A3(new_n677), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G317), .A2(new_n699), .B1(new_n739), .B2(G311), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT52), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n688), .A2(G303), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n360), .B1(new_n693), .B2(new_n710), .C1(new_n498), .C2(new_n701), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G116), .B2(new_n683), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G107), .A2(new_n706), .B1(new_n705), .B2(G283), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n736), .A2(new_n224), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G150), .A2(new_n699), .B1(new_n739), .B2(G159), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT51), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n684), .A2(new_n222), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n270), .B1(new_n312), .B2(new_n701), .C1(new_n689), .C2(new_n228), .ZN(new_n987));
  OR4_X1    g0787(.A1(new_n983), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n705), .A2(G68), .B1(G143), .B2(new_n694), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT112), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n982), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT113), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n678), .B1(new_n992), .B2(new_n944), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n247), .A2(new_n721), .B1(G97), .B2(new_n210), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n729), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT114), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n731), .B2(new_n891), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n974), .A2(new_n975), .A3(new_n997), .ZN(G390));
  NAND3_X1  g0798(.A1(new_n802), .A2(new_n775), .A3(new_n809), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT101), .B1(new_n812), .B2(new_n808), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n999), .A2(new_n726), .A3(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n360), .B1(new_n693), .B2(new_n498), .C1(new_n689), .C2(new_n424), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G97), .B2(new_n702), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n705), .A2(G87), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n737), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n697), .A2(new_n559), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1006), .B(new_n986), .C1(G283), .C2(new_n699), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT54), .B(G143), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n270), .B1(new_n701), .B2(new_n1010), .C1(new_n689), .C2(new_n741), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G50), .B2(new_n706), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT53), .B1(new_n857), .B2(new_n310), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n857), .A2(KEYINPUT53), .A3(new_n310), .ZN(new_n1014));
  INV_X1    g0814(.A(G132), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n684), .A2(new_n743), .B1(new_n697), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G128), .B2(new_n699), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(G125), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n693), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1008), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1021), .A2(new_n681), .B1(new_n312), .B2(new_n759), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n1001), .A2(new_n678), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n817), .A2(new_n821), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n774), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n999), .A2(new_n1000), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n764), .B1(new_n667), .B2(new_n763), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n821), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1025), .B(new_n838), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n656), .A2(new_n657), .A3(G330), .A4(new_n767), .ZN(new_n1031));
  OR3_X1    g0831(.A1(new_n1031), .A2(KEYINPUT115), .A3(new_n1029), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT115), .B1(new_n1031), .B2(new_n1029), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1027), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1031), .A2(new_n1029), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1023), .B1(new_n1040), .B2(new_n677), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT117), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n769), .A2(new_n656), .A3(G330), .A4(new_n657), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n1029), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1032), .A2(new_n1028), .A3(new_n1033), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1031), .A2(new_n1029), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n817), .B1(new_n1046), .B2(new_n1037), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n658), .A2(G330), .A3(new_n421), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n597), .A2(new_n828), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1027), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1038), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1051), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n931), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1042), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1039), .A2(KEYINPUT116), .A3(new_n1051), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT116), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n1060), .ZN(new_n1061));
  AND4_X1   g0861(.A1(new_n1042), .A2(new_n1057), .A3(new_n1059), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1041), .B1(new_n1058), .B2(new_n1062), .ZN(G378));
  NAND2_X1  g0863(.A1(new_n329), .A2(new_n333), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT55), .Z(new_n1065));
  NOR2_X1   g0865(.A1(new_n318), .A2(new_n618), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT56), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1065), .B(new_n1067), .Z(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(G330), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n837), .B2(new_n841), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n999), .A2(new_n1000), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n825), .B1(new_n1073), .B2(new_n774), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n1074), .B2(new_n824), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1025), .B1(new_n999), .B2(new_n1000), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n824), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n1071), .A4(new_n825), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1069), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n827), .A2(new_n1071), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1074), .A2(new_n824), .A3(new_n1072), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1068), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1050), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT119), .B1(new_n1056), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT119), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n1050), .C1(new_n1039), .C2(new_n1051), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1083), .A2(new_n1085), .A3(KEYINPUT57), .A4(new_n1087), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n972), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n739), .A2(G128), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n742), .B2(new_n1019), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n689), .A2(new_n1015), .B1(new_n310), .B2(new_n684), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(new_n705), .C2(new_n1009), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n741), .B2(new_n701), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n694), .A2(G124), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(KEYINPUT59), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(G33), .A2(G41), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT118), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n706), .B2(G159), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n228), .C1(G41), .C2(new_n270), .ZN(new_n1105));
  AOI211_X1 g0905(.A(G41), .B(new_n270), .C1(new_n694), .C2(G283), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n426), .B2(new_n689), .C1(new_n342), .C2(new_n701), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n736), .A2(new_n201), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n867), .B1(new_n424), .B2(new_n697), .C1(new_n742), .C2(new_n559), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1107), .A2(new_n960), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT58), .Z(new_n1111));
  AND3_X1   g0911(.A1(new_n1104), .A2(new_n1105), .A3(new_n1111), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n678), .B1(new_n944), .B2(new_n1112), .C1(new_n1069), .C2(new_n727), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n228), .B2(new_n759), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1083), .B2(new_n677), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1092), .A2(new_n1115), .ZN(G375));
  NAND3_X1  g0916(.A1(new_n1084), .A2(new_n1047), .A3(new_n1045), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1117), .A2(new_n1051), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n909), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT120), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n1029), .A2(new_n726), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n701), .A2(new_n424), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n688), .A2(G116), .B1(G303), .B2(new_n694), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n875), .A2(new_n360), .A3(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n857), .A2(new_n426), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n739), .A2(G283), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n962), .B(new_n1126), .C1(new_n742), .C2(new_n498), .ZN(new_n1127));
  OR4_X1    g0927(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n270), .B1(new_n701), .B2(new_n310), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1129), .B(new_n1108), .C1(G128), .C2(new_n694), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n684), .A2(new_n228), .B1(new_n697), .B2(new_n741), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G132), .B2(new_n699), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n743), .C2(new_n857), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n689), .A2(new_n1010), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n681), .B1(new_n202), .B2(new_n759), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1121), .A2(new_n678), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1048), .B2(new_n677), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1120), .A2(new_n1138), .ZN(G381));
  NAND2_X1  g0939(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1041), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(G375), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n933), .A2(new_n733), .A3(new_n970), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(G384), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n910), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT104), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n926), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n927), .ZN(new_n1149));
  INV_X1    g0949(.A(G390), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n888), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(G381), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1142), .A2(new_n1144), .A3(new_n1152), .ZN(G407));
  INV_X1    g0953(.A(G213), .ZN(new_n1154));
  OR3_X1    g0954(.A1(new_n1154), .A2(KEYINPUT121), .A3(G343), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT121), .B1(new_n1154), .B2(G343), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1154), .B1(new_n1142), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(G407), .ZN(G409));
  NAND3_X1  g0960(.A1(G378), .A2(new_n1092), .A3(new_n1115), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1141), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n909), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1115), .B1(new_n1088), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1158), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT60), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1118), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1117), .A2(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n972), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1138), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(G384), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT63), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(G393), .A2(G396), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n1143), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1150), .B1(new_n1149), .B2(new_n888), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n888), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1180), .B(G390), .C1(new_n1148), .C2(new_n927), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(G387), .A2(G390), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1151), .A3(new_n1177), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1173), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1166), .A2(KEYINPUT122), .A3(new_n1172), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1188), .A2(new_n1174), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT61), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1172), .B1(KEYINPUT123), .B2(new_n1157), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1158), .A2(G2897), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(new_n1166), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1186), .A2(new_n1190), .A3(new_n1191), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1191), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1198), .A2(KEYINPUT62), .A3(new_n1157), .A4(new_n1172), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT124), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1166), .A2(KEYINPUT124), .A3(KEYINPUT62), .A4(new_n1172), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT62), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1188), .A2(new_n1204), .A3(new_n1189), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1197), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1185), .B(KEYINPUT125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1196), .B1(new_n1206), .B2(new_n1207), .ZN(G405));
  AND3_X1   g1008(.A1(G378), .A2(new_n1092), .A3(new_n1115), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1141), .B1(new_n1092), .B2(new_n1115), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1172), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(G375), .A2(new_n1162), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1172), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1161), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1185), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT126), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT127), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1185), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1217), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1219), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1225), .A2(new_n1221), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1224), .A2(new_n1227), .ZN(G402));
endmodule


