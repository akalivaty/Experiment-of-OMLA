//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g028(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT67), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(KEYINPUT3), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n482), .A2(G137), .A3(new_n483), .A4(new_n472), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n481), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n485), .A2(G101), .A3(new_n483), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G160));
  AND2_X1   g064(.A1(new_n482), .A2(new_n472), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT70), .Z(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n483), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n483), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n493), .B(new_n496), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT71), .Z(G162));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n471), .A2(new_n474), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n482), .A2(new_n472), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n502), .A2(new_n504), .B1(new_n506), .B2(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n482), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n508));
  OR2_X1    g083(.A1(G102), .A2(G2105), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n509), .B(G2104), .C1(G114), .C2(new_n483), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n501), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n472), .A2(new_n473), .A3(KEYINPUT67), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT67), .B1(new_n472), .B2(new_n473), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n508), .A2(new_n510), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT72), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G164));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n527), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n532), .A2(G88), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(G50), .A3(G543), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n527), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n533), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND2_X1  g114(.A1(new_n532), .A2(G89), .ZN(new_n540));
  OR2_X1    g115(.A1(KEYINPUT6), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g117(.A1(KEYINPUT6), .A2(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(KEYINPUT6), .A2(G651), .ZN(new_n545));
  NOR2_X1   g120(.A1(KEYINPUT6), .A2(G651), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT75), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n547), .A3(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G51), .ZN(new_n550));
  AND2_X1   g125(.A1(G63), .A2(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n527), .A2(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n540), .A2(new_n550), .A3(new_n555), .ZN(G168));
  AND2_X1   g131(.A1(new_n532), .A2(G90), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G52), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n558), .A2(new_n536), .B1(new_n548), .B2(new_n559), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n557), .A2(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  AOI22_X1  g137(.A1(new_n532), .A2(G81), .B1(new_n549), .B2(G43), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n536), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND4_X1  g148(.A1(new_n544), .A2(new_n547), .A3(G53), .A4(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n523), .B1(new_n529), .B2(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n577), .A2(G53), .A3(new_n544), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT79), .B(G65), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n527), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n536), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n532), .B2(G91), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G299));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND2_X1  g166(.A1(new_n532), .A2(G87), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n527), .A2(G74), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n549), .A2(G49), .B1(new_n593), .B2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G288));
  AOI22_X1  g170(.A1(new_n527), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n536), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n529), .A2(G48), .A3(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n532), .A2(G86), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n532), .A2(G85), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n549), .A2(G47), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n536), .C2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n532), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n527), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n612), .A2(new_n536), .B1(new_n548), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n610), .A2(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND2_X1  g200(.A1(new_n565), .A2(new_n567), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n617), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(new_n627), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n485), .A2(new_n483), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n502), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n495), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n491), .A2(G123), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(G111), .ZN(new_n644));
  AOI22_X1  g219(.A1(new_n643), .A2(KEYINPUT81), .B1(new_n644), .B2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(KEYINPUT81), .B2(new_n643), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n639), .A2(new_n640), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI21_X1  g247(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT85), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G2096), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(new_n684), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT20), .Z(new_n688));
  AOI211_X1 g263(.A(new_n686), .B(new_n688), .C1(new_n681), .C2(new_n685), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT86), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G20), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT23), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n621), .B2(new_n697), .ZN(new_n700));
  INV_X1    g275(.A(G1956), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G35), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G162), .B2(new_n703), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2090), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT96), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT97), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n697), .A2(G6), .ZN(new_n712));
  INV_X1    g287(.A(G305), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n697), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT89), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT32), .B(G1981), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n697), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n697), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1971), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n697), .A2(G23), .ZN(new_n722));
  INV_X1    g297(.A(G288), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n697), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n717), .A2(new_n718), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT90), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n703), .A2(G25), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT87), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT87), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n491), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n483), .A2(G107), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G131), .B2(new_n495), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT88), .Z(new_n738));
  OAI211_X1 g313(.A(new_n731), .B(new_n732), .C1(new_n738), .C2(new_n703), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  MUX2_X1   g318(.A(G24), .B(G290), .S(G16), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1986), .ZN(new_n745));
  NOR3_X1   g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n729), .B(new_n746), .C1(KEYINPUT34), .C2(new_n727), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n748), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n483), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n752), .B(new_n754), .C1(G139), .C2(new_n495), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(new_n442), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n703), .B1(new_n759), .B2(G34), .ZN(new_n761));
  OAI22_X1  g336(.A1(new_n488), .A2(new_n703), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n703), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n634), .A2(G105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  NAND3_X1  g342(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT26), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n491), .B2(G129), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n495), .A2(G141), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT27), .B(G1996), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n758), .A2(new_n764), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n697), .A2(G5), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G171), .B2(new_n697), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G1961), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n757), .A2(new_n442), .B1(new_n762), .B2(new_n763), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n703), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n495), .A2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n491), .A2(G128), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n483), .A2(G116), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n777), .A2(new_n780), .A3(new_n781), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT92), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n629), .B2(new_n697), .ZN(new_n795));
  INV_X1    g370(.A(G1348), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n703), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n703), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2078), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n792), .B(new_n801), .C1(new_n706), .C2(G2090), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n697), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n568), .B2(new_n697), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT31), .B(G11), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT30), .B(G28), .Z(new_n807));
  NOR2_X1   g382(.A1(new_n647), .A2(new_n703), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n806), .B1(G29), .B2(new_n807), .C1(new_n808), .C2(KEYINPUT94), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(KEYINPUT94), .B2(new_n808), .ZN(new_n810));
  INV_X1    g385(.A(G1966), .ZN(new_n811));
  NOR2_X1   g386(.A1(G168), .A2(new_n697), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n697), .B2(G21), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n811), .A2(new_n813), .B1(new_n779), .B2(G1961), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n810), .B(new_n814), .C1(new_n811), .C2(new_n813), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT95), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n802), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n711), .A2(new_n749), .A3(new_n750), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n617), .A2(G559), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT38), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n527), .A2(G67), .ZN(new_n822));
  INV_X1    g397(.A(G80), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n523), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n536), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n532), .A2(G93), .B1(new_n549), .B2(G55), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n626), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n821), .B(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(G860), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n836), .ZN(G145));
  XNOR2_X1  g412(.A(G162), .B(new_n488), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n647), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n491), .A2(G130), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n483), .A2(G118), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G142), .B2(new_n495), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(new_n636), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n755), .B(new_n772), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n511), .B1(new_n513), .B2(new_n516), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n788), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n738), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n848), .B(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n840), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n840), .B2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g430(.A1(new_n829), .A2(new_n627), .ZN(new_n856));
  XNOR2_X1  g431(.A(G290), .B(G288), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(G303), .B(G305), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT42), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n830), .B(new_n630), .ZN(new_n866));
  OR2_X1    g441(.A1(G299), .A2(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g442(.A1(G299), .A2(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n617), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT100), .A3(G299), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT41), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n872), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n865), .B1(new_n877), .B2(KEYINPUT102), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(KEYINPUT102), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n878), .B(new_n879), .Z(new_n880));
  OAI21_X1  g455(.A(new_n856), .B1(new_n880), .B2(new_n627), .ZN(G295));
  OAI21_X1  g456(.A(new_n856), .B1(new_n880), .B2(new_n627), .ZN(G331));
  XNOR2_X1  g457(.A(new_n568), .B(new_n829), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n884));
  OR3_X1    g459(.A1(G301), .A2(new_n884), .A3(KEYINPUT104), .ZN(new_n885));
  AOI21_X1  g460(.A(G168), .B1(G301), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT104), .B1(G301), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n883), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n830), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n883), .A2(KEYINPUT105), .A3(new_n888), .A4(new_n891), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n874), .A3(new_n875), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n894), .A3(new_n873), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n864), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n899), .ZN(new_n903));
  INV_X1    g478(.A(new_n864), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(KEYINPUT43), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n871), .B1(new_n896), .B2(new_n897), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n892), .A2(new_n894), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n876), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n901), .B(new_n900), .C1(new_n910), .C2(new_n864), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(KEYINPUT43), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n905), .A2(new_n915), .A3(new_n901), .A4(new_n900), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT106), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n902), .A2(new_n918), .A3(new_n915), .A4(new_n905), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n914), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n914), .C1(new_n923), .C2(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(G397));
  NAND3_X1  g504(.A1(new_n478), .A2(G40), .A3(new_n487), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n478), .A2(KEYINPUT109), .A3(G40), .A4(new_n487), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n849), .B2(G1384), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G290), .A2(G1986), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n941));
  XOR2_X1   g516(.A(new_n940), .B(new_n941), .Z(new_n942));
  OR2_X1    g517(.A1(new_n738), .A2(new_n740), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n788), .B(new_n790), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n772), .B(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n738), .A2(new_n740), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n938), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n944), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n938), .B1(new_n950), .B2(new_n772), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n938), .A2(new_n945), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  NAND2_X1  g531(.A1(new_n946), .A2(new_n944), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n947), .A2(new_n957), .B1(G2067), .B2(new_n788), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n949), .B(new_n956), .C1(new_n938), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT123), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n517), .A2(new_n518), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n932), .A2(new_n933), .A3(new_n963), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n507), .A2(new_n501), .A3(new_n511), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT72), .B1(new_n517), .B2(new_n518), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n936), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n520), .B2(new_n962), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n932), .A2(new_n933), .A3(new_n963), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT110), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(G1971), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n520), .B2(new_n962), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n961), .A2(new_n976), .A3(new_n962), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n932), .A2(new_n933), .A3(new_n978), .ZN(new_n979));
  OR3_X1    g554(.A1(new_n977), .A2(new_n979), .A3(G2090), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G303), .A2(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT55), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(G8), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n527), .A2(new_n529), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT74), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT112), .B(G86), .Z(new_n993));
  NAND3_X1  g568(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n994), .B2(new_n598), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n597), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n989), .A3(new_n598), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n988), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(G305), .A2(G1981), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n987), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n999), .ZN(new_n1001));
  INV_X1    g576(.A(new_n997), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1002), .A2(new_n597), .A3(new_n995), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1001), .B(KEYINPUT49), .C1(new_n1003), .C2(new_n988), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n849), .A2(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n932), .A2(new_n1005), .A3(new_n933), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n723), .A2(G1976), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(G8), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  INV_X1    g586(.A(G1976), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(G288), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1007), .A2(new_n1009), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(G1976), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n999), .B1(new_n1008), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1007), .B(KEYINPUT114), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n986), .A2(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n985), .A2(new_n1016), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(new_n849), .B2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n932), .A2(new_n1023), .A3(new_n933), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2090), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n520), .A2(new_n976), .A3(new_n962), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n975), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT115), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n975), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1022), .B1(new_n983), .B2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n977), .A2(new_n979), .A3(G2084), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n932), .A2(new_n937), .A3(new_n933), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n520), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n932), .A2(new_n937), .A3(KEYINPUT116), .A4(new_n933), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1035), .B1(new_n1041), .B2(new_n811), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(G286), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT63), .B1(new_n1034), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n985), .A3(KEYINPUT63), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n975), .B2(new_n980), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n984), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1049), .B2(new_n1015), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1016), .B(KEYINPUT117), .C1(new_n984), .C2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1021), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1961), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n977), .B2(new_n979), .ZN(new_n1058));
  AOI21_X1  g633(.A(G2078), .B1(new_n970), .B2(new_n973), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1056), .B(new_n1058), .C1(new_n1059), .C2(KEYINPUT53), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1060), .A2(G171), .ZN(new_n1061));
  INV_X1    g636(.A(new_n930), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n937), .A2(new_n1062), .A3(new_n963), .A4(new_n1055), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1058), .C1(new_n1059), .C2(KEYINPUT53), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1054), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n964), .A2(new_n968), .A3(new_n1067), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT50), .B(G1384), .C1(new_n512), .C2(new_n519), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n701), .B1(new_n1024), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n588), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n991), .A2(G91), .A3(new_n992), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n580), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT118), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n576), .A2(new_n579), .A3(KEYINPUT78), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT78), .B1(new_n576), .B2(new_n579), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n589), .B(KEYINPUT57), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n584), .A2(KEYINPUT118), .A3(KEYINPUT57), .A4(new_n589), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1068), .A2(new_n1070), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n796), .B1(new_n977), .B2(new_n979), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n934), .A2(new_n790), .A3(new_n1005), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n629), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1081), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(new_n1081), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n617), .B2(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1082), .A2(new_n1083), .A3(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n617), .A2(KEYINPUT119), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1094), .B(new_n1095), .C1(new_n1084), .C2(KEYINPUT60), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1956), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1067), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n971), .A2(new_n972), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1087), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1091), .A2(new_n1096), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n964), .A2(new_n968), .A3(new_n945), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n1006), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n626), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1088), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1064), .A2(G171), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(KEYINPUT54), .C1(G171), .C2(new_n1060), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1066), .A2(new_n1034), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G168), .A2(new_n1043), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT51), .B1(new_n1118), .B2(KEYINPUT120), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1118), .B(new_n1120), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1041), .A2(new_n811), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n1035), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1043), .B(new_n1120), .C1(new_n1042), .C2(G168), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1116), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1043), .B1(new_n1042), .B2(G168), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1119), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(KEYINPUT121), .A3(new_n1123), .A4(new_n1121), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1115), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n960), .B1(new_n1053), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1129), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1033), .A2(new_n983), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1022), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1061), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT62), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1134), .A2(new_n1137), .A3(KEYINPUT124), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1110), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1107), .A2(KEYINPUT59), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n1096), .A3(new_n1102), .A4(new_n1091), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1060), .A2(G171), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(G171), .B2(new_n1064), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1148), .A2(new_n1088), .B1(new_n1150), .B2(new_n1054), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1141), .A3(new_n1034), .A4(new_n1114), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1135), .A2(new_n1136), .A3(new_n1044), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1052), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1152), .A2(new_n1157), .A3(KEYINPUT123), .A4(new_n1021), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1132), .A2(new_n1144), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G290), .B(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n938), .B1(new_n948), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1159), .A2(KEYINPUT125), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n959), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT127), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n959), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g743(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n854), .A2(new_n912), .A3(new_n1170), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


