//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  INV_X1    g009(.A(G15gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G22gat), .ZN(new_n212));
  INV_X1    g011(.A(G22gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G15gat), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(G1gat), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g015(.A(G8gat), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(G8gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n219), .C1(G1gat), .C2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n225), .A2(KEYINPUT14), .B1(new_n226), .B2(new_n224), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT90), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT90), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G29gat), .A3(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT92), .ZN(new_n234));
  INV_X1    g033(.A(G43gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(G50gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(G50gat), .ZN(new_n237));
  INV_X1    g036(.A(G50gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT92), .A3(G43gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT15), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(G43gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n237), .A2(new_n243), .A3(new_n244), .A4(KEYINPUT15), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT15), .B1(new_n235), .B2(G50gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n238), .A2(G43gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT91), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n242), .A3(new_n245), .A4(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n229), .A2(new_n231), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n251));
  NOR3_X1   g050(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(KEYINPUT89), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT89), .ZN(new_n254));
  NOR4_X1   g053(.A1(new_n254), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n246), .A2(new_n247), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT17), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n222), .B1(new_n259), .B2(KEYINPUT93), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT17), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n222), .B2(KEYINPUT93), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n249), .A2(new_n258), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n208), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT94), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n217), .A2(new_n221), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n226), .A2(new_n224), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n251), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n248), .A2(new_n250), .A3(new_n245), .A4(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n240), .A2(new_n241), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n257), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n269), .A2(new_n254), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n252), .A2(KEYINPUT89), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n251), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n277), .B2(new_n250), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n268), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n249), .A2(new_n258), .A3(new_n217), .A4(new_n221), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n207), .B(KEYINPUT13), .Z(new_n282));
  AOI21_X1  g081(.A(new_n267), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  AOI211_X1 g083(.A(KEYINPUT94), .B(new_n284), .C1(new_n279), .C2(new_n280), .ZN(new_n285));
  OAI22_X1  g084(.A1(new_n266), .A2(KEYINPUT18), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT18), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n287), .B(new_n208), .C1(new_n260), .C2(new_n265), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n206), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n265), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n207), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n263), .A2(new_n268), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n249), .A2(new_n258), .B1(new_n217), .B2(new_n221), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n282), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT94), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n267), .A3(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n266), .A2(KEYINPUT18), .ZN(new_n299));
  INV_X1    g098(.A(new_n206), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n292), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n289), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304));
  XOR2_X1   g103(.A(G211gat), .B(G218gat), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n307), .A2(new_n308), .B1(G211gat), .B2(G218gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n304), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G141gat), .B(G148gat), .Z(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(KEYINPUT77), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI221_X1 g124(.A(new_n321), .B1(new_n323), .B2(new_n318), .C1(new_n320), .C2(KEYINPUT77), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(KEYINPUT78), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n326), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n317), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n313), .B2(new_n314), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n310), .A2(new_n311), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n305), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT75), .A3(new_n312), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT3), .B1(new_n325), .B2(new_n326), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n333), .B(new_n336), .C1(new_n337), .C2(KEYINPUT29), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n331), .A2(G228gat), .A3(G233gat), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(KEYINPUT80), .Z(new_n342));
  AOI21_X1  g141(.A(new_n328), .B1(new_n315), .B2(new_n316), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n343), .A2(KEYINPUT81), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(KEYINPUT81), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT82), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(new_n342), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n340), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT31), .B(G50gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n213), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n213), .A2(KEYINPUT83), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n356), .B2(new_n353), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n350), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n333), .A2(new_n336), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n368));
  INV_X1    g167(.A(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n368), .A2(new_n372), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n367), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT65), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n372), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n378), .B(new_n379), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n380), .A3(new_n366), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n375), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n377), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT68), .ZN(new_n386));
  INV_X1    g185(.A(new_n361), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n386), .B(new_n366), .C1(KEYINPUT26), .C2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT27), .B(G183gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n370), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n390), .A2(KEYINPUT28), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n379), .B1(new_n390), .B2(KEYINPUT28), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G226gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT76), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n395), .B1(new_n384), .B2(new_n393), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n388), .A2(new_n391), .A3(new_n392), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n376), .A2(new_n373), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n400), .A2(new_n367), .B1(new_n382), .B2(new_n375), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n304), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n398), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n360), .B(new_n397), .C1(new_n403), .C2(KEYINPUT76), .ZN(new_n404));
  INV_X1    g203(.A(new_n398), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n405), .B1(new_n396), .B2(new_n394), .ZN(new_n406));
  INV_X1    g205(.A(new_n360), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XOR2_X1   g210(.A(new_n410), .B(new_n411), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n404), .A2(new_n408), .A3(new_n412), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(KEYINPUT30), .A3(new_n415), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n409), .A2(KEYINPUT30), .A3(new_n413), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT70), .B(G120gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G113gat), .ZN(new_n426));
  OR2_X1    g225(.A1(G113gat), .A2(G120gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G127gat), .B(G134gat), .ZN(new_n428));
  XOR2_X1   g227(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n429));
  NAND4_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(KEYINPUT69), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G127gat), .ZN(new_n434));
  OR3_X1    g233(.A1(new_n434), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n328), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT4), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n337), .A2(new_n437), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n330), .A2(new_n327), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n440), .B1(new_n441), .B2(new_n316), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n424), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT39), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n423), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n437), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n330), .A2(new_n446), .A3(new_n327), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n438), .ZN(new_n448));
  INV_X1    g247(.A(new_n424), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT39), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n445), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT40), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n439), .A2(new_n442), .A3(new_n424), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n448), .B2(new_n449), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n439), .A2(new_n442), .A3(new_n455), .A4(new_n424), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n423), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n445), .B(KEYINPUT40), .C1(new_n443), .C2(new_n450), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n453), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n359), .B1(new_n418), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n422), .B1(new_n457), .B2(new_n458), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(new_n422), .A3(new_n458), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n465), .B(new_n415), .C1(new_n468), .C2(new_n464), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n413), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n404), .A2(new_n408), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n406), .B2(new_n360), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n407), .B(new_n397), .C1(new_n403), .C2(KEYINPUT76), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n476), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n475), .B(KEYINPUT87), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n480), .A2(new_n479), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n413), .B(new_n471), .C1(new_n409), .C2(KEYINPUT37), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n409), .A2(KEYINPUT37), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n413), .B1(new_n473), .B2(new_n474), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT88), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(KEYINPUT88), .B(new_n413), .C1(new_n473), .C2(new_n474), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n471), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n463), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n350), .A2(new_n358), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n357), .B(new_n340), .C1(new_n347), .C2(new_n349), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n467), .B(new_n466), .C1(new_n464), .C2(KEYINPUT79), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n465), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n416), .A2(new_n417), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n384), .A2(new_n393), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n437), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n384), .A2(new_n446), .A3(new_n393), .ZN(new_n504));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT64), .Z(new_n506));
  NAND3_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT32), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT33), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(KEYINPUT72), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(new_n211), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(new_n235), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n514), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT32), .B(new_n507), .C1(new_n516), .C2(new_n509), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n504), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n505), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT34), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(KEYINPUT34), .A2(new_n520), .B1(new_n523), .B2(KEYINPUT73), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(new_n515), .A3(new_n526), .A4(new_n517), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n530), .A3(KEYINPUT36), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT36), .B1(new_n528), .B2(new_n530), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT84), .B1(new_n501), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n533), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT79), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n460), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n466), .A2(new_n467), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n543), .A2(new_n465), .B1(new_n417), .B2(new_n416), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n537), .B(new_n538), .C1(new_n544), .C2(new_n496), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n493), .A2(new_n535), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n528), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n518), .A2(new_n527), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n499), .A2(new_n549), .A3(new_n496), .A4(new_n500), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT35), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(new_n460), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT35), .B1(new_n552), .B2(new_n465), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(new_n496), .A3(new_n549), .A4(new_n500), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n303), .B1(new_n546), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT98), .A3(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(G85gat), .A3(G92gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT99), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n561), .A2(new_n564), .A3(new_n568), .A4(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n561), .A2(new_n571), .B1(new_n568), .B2(new_n564), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT41), .ZN(new_n576));
  NAND2_X1  g375(.A1(G232gat), .A2(G233gat), .ZN(new_n577));
  OAI22_X1  g376(.A1(new_n264), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n578), .A2(KEYINPUT100), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n259), .A2(new_n573), .A3(new_n574), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n261), .B2(new_n263), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(KEYINPUT100), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(KEYINPUT101), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(KEYINPUT101), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n577), .A2(new_n576), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n583), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n583), .B2(new_n585), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n594), .A2(new_n597), .B1(new_n600), .B2(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(G64gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(G57gat), .ZN(new_n603));
  INV_X1    g402(.A(G57gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(G64gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n597), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(G64gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n602), .A2(G57gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(G71gat), .A2(G78gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n597), .B(new_n610), .C1(new_n613), .C2(new_n594), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT21), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n268), .B1(KEYINPUT21), .B2(new_n615), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT97), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT96), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n620), .B(new_n627), .Z(new_n628));
  NOR2_X1   g427(.A1(new_n593), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n615), .B1(new_n573), .B2(new_n574), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n561), .A2(new_n571), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n568), .A2(new_n564), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n614), .A3(new_n607), .A4(new_n572), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n615), .B(KEYINPUT10), .C1(new_n573), .C2(new_n574), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n630), .A2(new_n635), .ZN(new_n641));
  INV_X1    g440(.A(new_n639), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G120gat), .B(G148gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(G176gat), .B(G204gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n643), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n629), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n556), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n499), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT102), .B(G1gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1324gat));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n500), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n219), .B2(new_n659), .ZN(new_n662));
  MUX2_X1   g461(.A(new_n661), .B(new_n662), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n655), .B2(new_n537), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n549), .A2(new_n211), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n655), .B2(new_n665), .ZN(G1326gat));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n655), .B2(new_n496), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n556), .A2(KEYINPUT103), .A3(new_n359), .A4(new_n654), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  INV_X1    g471(.A(new_n593), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n628), .A2(new_n652), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n556), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n499), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n223), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n546), .A2(new_n555), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n673), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n501), .A2(new_n534), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n493), .A2(new_n685), .B1(new_n551), .B2(new_n554), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n682), .B1(new_n686), .B2(new_n673), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n289), .A2(KEYINPUT104), .A3(new_n301), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n289), .B2(new_n301), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n674), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n499), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n679), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n695), .A3(new_n696), .ZN(G1328gat));
  NAND4_X1  g496(.A1(new_n556), .A2(new_n224), .A3(new_n418), .A4(new_n675), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT46), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n699), .A2(KEYINPUT106), .A3(new_n700), .A4(new_n701), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n694), .B2(new_n500), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(G1329gat));
  NAND4_X1  g508(.A1(new_n684), .A2(new_n687), .A3(new_n534), .A4(new_n693), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n235), .B1(new_n710), .B2(KEYINPUT108), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT108), .B2(new_n710), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n676), .A2(new_n235), .A3(new_n549), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(G43gat), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n713), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(G1330gat));
  NOR2_X1   g518(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n496), .A2(G50gat), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n676), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n684), .A2(new_n687), .A3(new_n359), .A4(new_n693), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G50gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n493), .A2(new_n685), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n555), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n691), .A2(new_n628), .A3(new_n593), .A4(new_n652), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n499), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(new_n604), .ZN(G1332gat));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n731), .B(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n735), .A2(new_n418), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  NAND3_X1  g539(.A1(new_n735), .A2(G71gat), .A3(new_n534), .ZN(new_n741));
  INV_X1    g540(.A(new_n549), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n598), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n741), .A2(KEYINPUT50), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT50), .B1(new_n741), .B2(new_n743), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(G1334gat));
  NAND2_X1  g545(.A1(new_n735), .A2(new_n359), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(G78gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1335gat));
  INV_X1    g548(.A(new_n628), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n691), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n652), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n688), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(new_n677), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n673), .B1(new_n728), .B2(new_n555), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT51), .B1(new_n756), .B2(new_n751), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n686), .A2(new_n759), .A3(new_n673), .A4(new_n752), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n761), .A3(KEYINPUT112), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n677), .A2(new_n569), .A3(new_n651), .ZN(new_n766));
  OAI22_X1  g565(.A1(new_n755), .A2(new_n569), .B1(new_n765), .B2(new_n766), .ZN(G1336gat));
  NOR3_X1   g566(.A1(new_n500), .A2(G92gat), .A3(new_n652), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n762), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n684), .A2(new_n687), .A3(new_n418), .A4(new_n753), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n768), .B1(new_n757), .B2(new_n760), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n774), .B1(new_n776), .B2(KEYINPUT52), .ZN(new_n777));
  AOI211_X1 g576(.A(KEYINPUT113), .B(new_n770), .C1(new_n772), .C2(new_n775), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(G1337gat));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n534), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n742), .A2(G99gat), .A3(new_n652), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n765), .B2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n496), .A2(G106gat), .A3(new_n652), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n762), .A2(new_n764), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n684), .A2(new_n687), .A3(new_n359), .A4(new_n753), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n758), .A2(new_n761), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n790), .A2(new_n784), .B1(G106gat), .B2(new_n786), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n785), .A2(new_n789), .B1(new_n791), .B2(new_n788), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n291), .A2(new_n287), .B1(new_n296), .B2(new_n297), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n300), .B1(new_n794), .B2(new_n299), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n286), .A2(new_n206), .A3(new_n288), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n642), .B1(new_n636), .B2(new_n637), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n647), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(new_n802), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(new_n650), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n289), .A2(new_n301), .A3(KEYINPUT104), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n800), .A3(new_n801), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n638), .A2(new_n801), .A3(new_n639), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n648), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n809), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n802), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(KEYINPUT115), .A3(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n797), .A2(new_n807), .A3(new_n808), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n260), .A2(new_n265), .A3(new_n208), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n282), .B2(new_n281), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n205), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(new_n301), .A3(new_n651), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n593), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT115), .B1(new_n817), .B2(new_n809), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n815), .B(KEYINPUT55), .C1(new_n799), .C2(new_n802), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n805), .A2(new_n650), .A3(new_n806), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n826), .A2(new_n301), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n593), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT117), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n827), .B1(new_n691), .B2(new_n834), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n839), .B(new_n836), .C1(new_n840), .C2(new_n593), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n841), .A3(new_n628), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n692), .A2(new_n629), .A3(new_n652), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n499), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n549), .A2(new_n496), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n418), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848), .B2(new_n691), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n843), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n496), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT118), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n853), .A3(new_n496), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n677), .A2(new_n500), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n742), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n302), .A2(G113gat), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n849), .B1(new_n859), .B2(new_n860), .ZN(G1340gat));
  OAI21_X1  g660(.A(G120gat), .B1(new_n858), .B2(new_n652), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n652), .A2(new_n425), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n847), .B2(new_n863), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n858), .B2(new_n628), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n434), .A3(new_n750), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1342gat));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n677), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n500), .A2(new_n593), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n868), .A2(G134gat), .A3(new_n845), .A4(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n858), .B2(new_n673), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n537), .A2(new_n359), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n844), .B2(KEYINPUT119), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n303), .A2(G141gat), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT120), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n500), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n856), .A2(new_n534), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n850), .B2(new_n359), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n359), .A2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n807), .A2(new_n302), .A3(new_n814), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n593), .B1(new_n828), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n628), .B1(new_n837), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n889), .B2(new_n843), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n303), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n881), .A2(new_n882), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n877), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n418), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n691), .B(new_n883), .C1(new_n884), .C2(new_n890), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(new_n880), .B1(G141gat), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n897), .B2(new_n882), .ZN(G1344gat));
  AOI21_X1  g697(.A(new_n886), .B1(new_n842), .B2(new_n843), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n654), .A2(new_n303), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n901), .B2(new_n359), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n651), .B(new_n883), .C1(new_n899), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G148gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n651), .B(new_n883), .C1(new_n884), .C2(new_n890), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  AOI22_X1  g706(.A1(KEYINPUT59), .A2(new_n904), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n652), .A2(G148gat), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n418), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT121), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n878), .A2(new_n500), .A3(new_n909), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n905), .A2(new_n907), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n906), .B1(new_n903), .B2(G148gat), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n912), .A2(new_n917), .ZN(G1345gat));
  INV_X1    g717(.A(G155gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n895), .A2(new_n919), .A3(new_n750), .ZN(new_n920));
  OAI21_X1  g719(.A(G155gat), .B1(new_n891), .B2(new_n628), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  OAI21_X1  g721(.A(G162gat), .B1(new_n891), .B2(new_n673), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n869), .A2(G162gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n894), .B2(new_n924), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n677), .B1(new_n842), .B2(new_n843), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n845), .A2(new_n500), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n691), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n418), .A2(new_n499), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n930), .A2(new_n742), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n932), .B1(new_n852), .B2(new_n854), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n302), .A2(G169gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  AOI21_X1  g734(.A(G176gat), .B1(new_n928), .B2(new_n651), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n651), .A2(G176gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n933), .B2(new_n937), .ZN(G1349gat));
  NAND2_X1  g737(.A1(new_n855), .A2(new_n931), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n939), .B2(new_n628), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n750), .A2(new_n389), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT122), .B1(new_n928), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n369), .B1(new_n933), .B2(new_n750), .ZN(new_n946));
  INV_X1    g745(.A(new_n944), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT60), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n939), .B2(new_n673), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g751(.A(KEYINPUT61), .B(G190gat), .C1(new_n939), .C2(new_n673), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n928), .A2(new_n370), .A3(new_n593), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(G1351gat));
  AND4_X1   g756(.A1(new_n359), .A2(new_n926), .A3(new_n418), .A4(new_n537), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n691), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n899), .A2(new_n902), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n534), .A2(new_n930), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT124), .ZN(new_n963));
  INV_X1    g762(.A(G197gat), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n963), .A2(new_n964), .A3(new_n303), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n959), .B1(new_n961), .B2(new_n965), .ZN(G1352gat));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n967), .A3(new_n651), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n961), .A2(new_n651), .ZN(new_n970));
  OAI21_X1  g769(.A(G204gat), .B1(new_n970), .B2(new_n963), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(G1353gat));
  INV_X1    g772(.A(G211gat), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n958), .A2(new_n974), .A3(new_n750), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n750), .B(new_n962), .C1(new_n899), .C2(new_n902), .ZN(new_n976));
  AND2_X1   g775(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n977));
  OAI21_X1  g776(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n975), .B(KEYINPUT126), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1354gat));
  AOI21_X1  g785(.A(G218gat), .B1(new_n958), .B2(new_n593), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n593), .A2(G218gat), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n960), .A2(new_n963), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n987), .A2(new_n990), .ZN(G1355gat));
endmodule


