

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736;

  INV_X1 U371 ( .A(G953), .ZN(n728) );
  NOR2_X1 U372 ( .A1(n561), .A2(n560), .ZN(n633) );
  NAND2_X2 U373 ( .A1(n605), .A2(n604), .ZN(n691) );
  XNOR2_X2 U374 ( .A(n570), .B(n394), .ZN(n560) );
  XNOR2_X1 U375 ( .A(n351), .B(KEYINPUT66), .ZN(n436) );
  INV_X1 U376 ( .A(G101), .ZN(n351) );
  NOR2_X1 U377 ( .A1(n540), .A2(n539), .ZN(n559) );
  XNOR2_X1 U378 ( .A(n540), .B(KEYINPUT1), .ZN(n502) );
  OR2_X1 U379 ( .A1(n607), .A2(n388), .ZN(n391) );
  XNOR2_X1 U380 ( .A(G122), .B(G104), .ZN(n409) );
  NAND2_X1 U381 ( .A1(n621), .A2(n630), .ZN(n484) );
  XNOR2_X1 U382 ( .A(n461), .B(n460), .ZN(n540) );
  NAND2_X1 U383 ( .A1(n358), .A2(n356), .ZN(n355) );
  AND2_X1 U384 ( .A1(n360), .A2(n348), .ZN(n359) );
  NOR2_X1 U385 ( .A1(n357), .A2(n400), .ZN(n356) );
  AND2_X1 U386 ( .A1(n492), .A2(n734), .ZN(n495) );
  XNOR2_X1 U387 ( .A(n556), .B(KEYINPUT46), .ZN(n557) );
  AND2_X1 U388 ( .A1(n498), .A2(n499), .ZN(n500) );
  NOR2_X1 U389 ( .A1(n547), .A2(n536), .ZN(n564) );
  XNOR2_X1 U390 ( .A(KEYINPUT16), .B(G110), .ZN(n381) );
  AND2_X1 U391 ( .A1(n724), .A2(n603), .ZN(n352) );
  XNOR2_X1 U392 ( .A(n366), .B(n365), .ZN(n364) );
  INV_X1 U393 ( .A(KEYINPUT34), .ZN(n365) );
  NAND2_X1 U394 ( .A1(n677), .A2(n507), .ZN(n366) );
  OR2_X1 U395 ( .A1(n502), .A2(n652), .ZN(n480) );
  INV_X1 U396 ( .A(n648), .ZN(n647) );
  NAND2_X1 U397 ( .A1(n507), .A2(n433), .ZN(n435) );
  BUF_X1 U398 ( .A(n691), .Z(n702) );
  XNOR2_X1 U399 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U400 ( .A(n722), .B(n454), .ZN(n459) );
  INV_X1 U401 ( .A(G110), .ZN(n456) );
  NOR2_X1 U402 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U403 ( .A(G131), .B(G140), .ZN(n401) );
  XOR2_X1 U404 ( .A(n450), .B(KEYINPUT68), .Z(n462) );
  XNOR2_X1 U405 ( .A(G137), .B(G140), .ZN(n450) );
  XNOR2_X1 U406 ( .A(n444), .B(n368), .ZN(n451) );
  XNOR2_X1 U407 ( .A(n369), .B(G134), .ZN(n368) );
  INV_X1 U408 ( .A(G131), .ZN(n369) );
  INV_X1 U409 ( .A(KEYINPUT82), .ZN(n383) );
  AND2_X1 U410 ( .A1(n568), .A2(n635), .ZN(n592) );
  INV_X1 U411 ( .A(n371), .ZN(n357) );
  XNOR2_X1 U412 ( .A(G134), .B(G122), .ZN(n417) );
  XNOR2_X1 U413 ( .A(n451), .B(n367), .ZN(n722) );
  INV_X1 U414 ( .A(n462), .ZN(n367) );
  XNOR2_X1 U415 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U416 ( .A(n488), .B(n372), .ZN(n677) );
  NOR2_X1 U417 ( .A1(n502), .A2(n487), .ZN(n488) );
  XNOR2_X1 U418 ( .A(n370), .B(n476), .ZN(n477) );
  INV_X1 U419 ( .A(n656), .ZN(n543) );
  INV_X1 U420 ( .A(KEYINPUT2), .ZN(n353) );
  XNOR2_X1 U421 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n554) );
  XNOR2_X1 U422 ( .A(n491), .B(n490), .ZN(n734) );
  NAND2_X1 U423 ( .A1(n364), .A2(n489), .ZN(n491) );
  NOR2_X1 U424 ( .A1(n480), .A2(n363), .ZN(n362) );
  INV_X1 U425 ( .A(n565), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n505), .B(KEYINPUT31), .ZN(n638) );
  OR2_X1 U427 ( .A1(n504), .A2(n503), .ZN(n505) );
  NOR2_X1 U428 ( .A1(n695), .A2(n706), .ZN(n698) );
  XNOR2_X1 U429 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U430 ( .A1(n611), .A2(n706), .ZN(n612) );
  OR2_X1 U431 ( .A1(n371), .A2(KEYINPUT0), .ZN(n348) );
  XNOR2_X1 U432 ( .A(n391), .B(n390), .ZN(n529) );
  XNOR2_X1 U433 ( .A(n484), .B(KEYINPUT81), .ZN(n498) );
  XOR2_X1 U434 ( .A(n574), .B(n573), .Z(n349) );
  AND2_X1 U435 ( .A1(n601), .A2(KEYINPUT2), .ZN(n350) );
  NOR2_X2 U436 ( .A1(n587), .A2(n586), .ZN(n588) );
  AND2_X2 U437 ( .A1(n600), .A2(n599), .ZN(n724) );
  XNOR2_X1 U438 ( .A(n486), .B(KEYINPUT67), .ZN(n648) );
  NAND2_X1 U439 ( .A1(n352), .A2(n710), .ZN(n604) );
  NAND2_X1 U440 ( .A1(n724), .A2(n710), .ZN(n354) );
  NAND2_X1 U441 ( .A1(n354), .A2(n350), .ZN(n605) );
  XNOR2_X1 U442 ( .A(n354), .B(n353), .ZN(n683) );
  NAND2_X2 U443 ( .A1(n359), .A2(n355), .ZN(n507) );
  INV_X1 U444 ( .A(n560), .ZN(n358) );
  NAND2_X1 U445 ( .A1(n560), .A2(n400), .ZN(n360) );
  XNOR2_X2 U446 ( .A(n361), .B(KEYINPUT32), .ZN(n621) );
  NAND2_X1 U447 ( .A1(n482), .A2(n565), .ZN(n517) );
  NAND2_X1 U448 ( .A1(n482), .A2(n362), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n615), .B(n374), .ZN(n617) );
  AND2_X1 U450 ( .A1(G217), .A2(n473), .ZN(n370) );
  OR2_X1 U451 ( .A1(n399), .A2(n534), .ZN(n371) );
  XNOR2_X1 U452 ( .A(KEYINPUT101), .B(KEYINPUT33), .ZN(n372) );
  AND2_X1 U453 ( .A1(n437), .A2(G210), .ZN(n373) );
  XOR2_X1 U454 ( .A(n614), .B(n613), .Z(n374) );
  NOR2_X1 U455 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U456 ( .A(KEYINPUT109), .ZN(n569) );
  XNOR2_X1 U457 ( .A(n443), .B(n442), .ZN(n445) );
  XNOR2_X1 U458 ( .A(n592), .B(n569), .ZN(n572) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(KEYINPUT110), .ZN(n573) );
  XNOR2_X1 U460 ( .A(n459), .B(n458), .ZN(n687) );
  INV_X1 U461 ( .A(n706), .ZN(n616) );
  XNOR2_X1 U462 ( .A(n687), .B(n686), .ZN(n688) );
  BUF_X1 U463 ( .A(n529), .Z(n596) );
  XNOR2_X1 U464 ( .A(n555), .B(n554), .ZN(n733) );
  XNOR2_X2 U465 ( .A(G146), .B(G125), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n436), .B(n407), .ZN(n375) );
  XNOR2_X2 U467 ( .A(G143), .B(G128), .ZN(n419) );
  XNOR2_X1 U468 ( .A(n419), .B(KEYINPUT4), .ZN(n444) );
  XNOR2_X1 U469 ( .A(n375), .B(n444), .ZN(n380) );
  XOR2_X1 U470 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n378) );
  NAND2_X1 U471 ( .A1(G224), .A2(n728), .ZN(n376) );
  XNOR2_X1 U472 ( .A(n376), .B(KEYINPUT17), .ZN(n377) );
  XNOR2_X1 U473 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U474 ( .A(n380), .B(n379), .ZN(n387) );
  XNOR2_X1 U475 ( .A(n409), .B(n381), .ZN(n382) );
  XNOR2_X1 U476 ( .A(G116), .B(G107), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n382), .B(n420), .ZN(n386) );
  XNOR2_X1 U478 ( .A(n383), .B(KEYINPUT3), .ZN(n385) );
  XNOR2_X1 U479 ( .A(G119), .B(G113), .ZN(n384) );
  XNOR2_X1 U480 ( .A(n385), .B(n384), .ZN(n441) );
  XNOR2_X1 U481 ( .A(n386), .B(n441), .ZN(n715) );
  XNOR2_X1 U482 ( .A(n387), .B(n715), .ZN(n607) );
  XNOR2_X1 U483 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  INV_X1 U484 ( .A(n602), .ZN(n388) );
  INV_X1 U485 ( .A(G902), .ZN(n446) );
  INV_X1 U486 ( .A(G237), .ZN(n389) );
  NAND2_X1 U487 ( .A1(n446), .A2(n389), .ZN(n392) );
  AND2_X1 U488 ( .A1(n392), .A2(G210), .ZN(n390) );
  NAND2_X1 U489 ( .A1(n392), .A2(G214), .ZN(n393) );
  XNOR2_X1 U490 ( .A(n393), .B(KEYINPUT83), .ZN(n664) );
  INV_X1 U491 ( .A(n664), .ZN(n591) );
  NAND2_X1 U492 ( .A1(n529), .A2(n591), .ZN(n570) );
  INV_X1 U493 ( .A(KEYINPUT19), .ZN(n394) );
  NAND2_X1 U494 ( .A1(G234), .A2(G237), .ZN(n395) );
  XNOR2_X1 U495 ( .A(n395), .B(KEYINPUT14), .ZN(n398) );
  NAND2_X1 U496 ( .A1(G902), .A2(n398), .ZN(n396) );
  XOR2_X1 U497 ( .A(KEYINPUT84), .B(n396), .Z(n397) );
  NAND2_X1 U498 ( .A1(G953), .A2(n397), .ZN(n532) );
  NOR2_X1 U499 ( .A1(n532), .A2(G898), .ZN(n399) );
  NAND2_X1 U500 ( .A1(G952), .A2(n398), .ZN(n675) );
  NOR2_X1 U501 ( .A1(n675), .A2(G953), .ZN(n534) );
  INV_X1 U502 ( .A(KEYINPUT0), .ZN(n400) );
  XNOR2_X1 U503 ( .A(KEYINPUT13), .B(KEYINPUT93), .ZN(n414) );
  XOR2_X1 U504 ( .A(KEYINPUT12), .B(KEYINPUT92), .Z(n402) );
  XNOR2_X1 U505 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U506 ( .A(KEYINPUT11), .B(KEYINPUT91), .Z(n404) );
  NOR2_X1 U507 ( .A1(G953), .A2(G237), .ZN(n437) );
  NAND2_X1 U508 ( .A1(G214), .A2(n437), .ZN(n403) );
  XNOR2_X1 U509 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U510 ( .A(n406), .B(n405), .ZN(n412) );
  XNOR2_X1 U511 ( .A(n407), .B(KEYINPUT10), .ZN(n721) );
  XNOR2_X1 U512 ( .A(G143), .B(G113), .ZN(n408) );
  XNOR2_X1 U513 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U514 ( .A(n721), .B(n410), .ZN(n411) );
  XNOR2_X1 U515 ( .A(n412), .B(n411), .ZN(n692) );
  NOR2_X1 U516 ( .A1(G902), .A2(n692), .ZN(n413) );
  XNOR2_X1 U517 ( .A(n414), .B(n413), .ZN(n416) );
  INV_X1 U518 ( .A(G475), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n416), .B(n415), .ZN(n511) );
  XNOR2_X1 U520 ( .A(KEYINPUT97), .B(G478), .ZN(n429) );
  XOR2_X1 U521 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n418) );
  XNOR2_X1 U522 ( .A(n418), .B(n417), .ZN(n424) );
  XNOR2_X1 U523 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U524 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n421) );
  XNOR2_X1 U525 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U526 ( .A(n424), .B(n423), .Z(n427) );
  NAND2_X1 U527 ( .A1(G234), .A2(n728), .ZN(n425) );
  XOR2_X1 U528 ( .A(KEYINPUT8), .B(n425), .Z(n463) );
  NAND2_X1 U529 ( .A1(G217), .A2(n463), .ZN(n426) );
  XNOR2_X1 U530 ( .A(n427), .B(n426), .ZN(n699) );
  NOR2_X1 U531 ( .A1(G902), .A2(n699), .ZN(n428) );
  XNOR2_X1 U532 ( .A(n429), .B(n428), .ZN(n512) );
  OR2_X1 U533 ( .A1(n511), .A2(n512), .ZN(n528) );
  XOR2_X1 U534 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n431) );
  NAND2_X1 U535 ( .A1(G234), .A2(n602), .ZN(n430) );
  XNOR2_X1 U536 ( .A(n431), .B(n430), .ZN(n473) );
  AND2_X1 U537 ( .A1(n473), .A2(G221), .ZN(n432) );
  XNOR2_X1 U538 ( .A(n432), .B(KEYINPUT21), .ZN(n651) );
  INV_X1 U539 ( .A(n651), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n528), .A2(n485), .ZN(n433) );
  INV_X1 U541 ( .A(KEYINPUT22), .ZN(n434) );
  XNOR2_X2 U542 ( .A(n435), .B(n434), .ZN(n482) );
  XOR2_X1 U543 ( .A(n436), .B(G146), .Z(n455) );
  XNOR2_X1 U544 ( .A(n455), .B(n373), .ZN(n443) );
  XOR2_X1 U545 ( .A(G116), .B(KEYINPUT90), .Z(n439) );
  XNOR2_X1 U546 ( .A(G137), .B(KEYINPUT5), .ZN(n438) );
  XNOR2_X1 U547 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U548 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U549 ( .A(n445), .B(n451), .ZN(n614) );
  NAND2_X1 U550 ( .A1(n614), .A2(n446), .ZN(n448) );
  INV_X1 U551 ( .A(G472), .ZN(n447) );
  XNOR2_X2 U552 ( .A(n448), .B(n447), .ZN(n656) );
  INV_X1 U553 ( .A(KEYINPUT6), .ZN(n449) );
  XNOR2_X1 U554 ( .A(n656), .B(n449), .ZN(n565) );
  NAND2_X1 U555 ( .A1(G227), .A2(n728), .ZN(n453) );
  INV_X1 U556 ( .A(G107), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n455), .B(G104), .ZN(n457) );
  NOR2_X1 U558 ( .A1(G902), .A2(n687), .ZN(n461) );
  XNOR2_X1 U559 ( .A(KEYINPUT70), .B(G469), .ZN(n460) );
  XNOR2_X1 U560 ( .A(n721), .B(n462), .ZN(n465) );
  NAND2_X1 U561 ( .A1(G221), .A2(n463), .ZN(n464) );
  XNOR2_X1 U562 ( .A(n465), .B(n464), .ZN(n472) );
  XOR2_X1 U563 ( .A(KEYINPUT23), .B(KEYINPUT74), .Z(n467) );
  XNOR2_X1 U564 ( .A(KEYINPUT85), .B(KEYINPUT24), .ZN(n466) );
  XNOR2_X1 U565 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U566 ( .A(n468), .B(G110), .Z(n470) );
  XNOR2_X1 U567 ( .A(G128), .B(G119), .ZN(n469) );
  XNOR2_X1 U568 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n472), .B(n471), .ZN(n704) );
  NOR2_X1 U570 ( .A1(n704), .A2(G902), .ZN(n478) );
  XOR2_X1 U571 ( .A(KEYINPUT86), .B(KEYINPUT25), .Z(n475) );
  XNOR2_X1 U572 ( .A(KEYINPUT73), .B(KEYINPUT88), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X2 U574 ( .A(n478), .B(n477), .ZN(n535) );
  INV_X1 U575 ( .A(KEYINPUT100), .ZN(n479) );
  XNOR2_X1 U576 ( .A(n535), .B(n479), .ZN(n652) );
  AND2_X1 U577 ( .A1(n656), .A2(n535), .ZN(n481) );
  AND2_X1 U578 ( .A1(n502), .A2(n481), .ZN(n483) );
  NAND2_X1 U579 ( .A1(n483), .A2(n482), .ZN(n630) );
  XNOR2_X1 U580 ( .A(n498), .B(KEYINPUT80), .ZN(n492) );
  NOR2_X1 U581 ( .A1(n485), .A2(n535), .ZN(n486) );
  OR2_X1 U582 ( .A1(n648), .A2(n565), .ZN(n487) );
  NAND2_X1 U583 ( .A1(n511), .A2(n512), .ZN(n577) );
  INV_X1 U584 ( .A(n577), .ZN(n489) );
  INV_X1 U585 ( .A(KEYINPUT35), .ZN(n490) );
  INV_X1 U586 ( .A(KEYINPUT44), .ZN(n493) );
  NAND2_X1 U587 ( .A1(n495), .A2(n493), .ZN(n494) );
  INV_X1 U588 ( .A(KEYINPUT71), .ZN(n499) );
  NAND2_X1 U589 ( .A1(n494), .A2(n499), .ZN(n497) );
  NAND2_X1 U590 ( .A1(n495), .A2(KEYINPUT71), .ZN(n496) );
  NAND2_X1 U591 ( .A1(n497), .A2(n496), .ZN(n525) );
  NAND2_X1 U592 ( .A1(n734), .A2(n500), .ZN(n501) );
  NAND2_X1 U593 ( .A1(n501), .A2(KEYINPUT44), .ZN(n523) );
  NOR2_X1 U594 ( .A1(n502), .A2(n656), .ZN(n646) );
  INV_X1 U595 ( .A(n646), .ZN(n504) );
  NAND2_X1 U596 ( .A1(n647), .A2(n507), .ZN(n503) );
  INV_X1 U597 ( .A(n540), .ZN(n506) );
  NAND2_X1 U598 ( .A1(n506), .A2(n647), .ZN(n548) );
  INV_X1 U599 ( .A(n507), .ZN(n508) );
  NOR2_X1 U600 ( .A1(n548), .A2(n508), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n509), .B(KEYINPUT89), .ZN(n510) );
  NOR2_X1 U602 ( .A1(n543), .A2(n510), .ZN(n627) );
  NOR2_X1 U603 ( .A1(n638), .A2(n627), .ZN(n515) );
  XOR2_X1 U604 ( .A(KEYINPUT94), .B(n511), .Z(n513) );
  NOR2_X1 U605 ( .A1(n513), .A2(n512), .ZN(n635) );
  INV_X1 U606 ( .A(n635), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U608 ( .A(n514), .B(KEYINPUT98), .Z(n639) );
  INV_X1 U609 ( .A(n639), .ZN(n589) );
  NAND2_X1 U610 ( .A1(n553), .A2(n589), .ZN(n662) );
  INV_X1 U611 ( .A(n662), .ZN(n580) );
  OR2_X1 U612 ( .A1(n515), .A2(n580), .ZN(n516) );
  XNOR2_X1 U613 ( .A(n516), .B(KEYINPUT99), .ZN(n521) );
  AND2_X1 U614 ( .A1(n502), .A2(n652), .ZN(n519) );
  XNOR2_X1 U615 ( .A(n517), .B(KEYINPUT79), .ZN(n518) );
  NAND2_X1 U616 ( .A1(n519), .A2(n518), .ZN(n622) );
  INV_X1 U617 ( .A(n622), .ZN(n520) );
  NOR2_X1 U618 ( .A1(n521), .A2(n520), .ZN(n522) );
  AND2_X1 U619 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U620 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U621 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n526) );
  XNOR2_X1 U622 ( .A(n527), .B(n526), .ZN(n710) );
  XOR2_X1 U623 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n542) );
  XOR2_X1 U624 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n531) );
  INV_X1 U625 ( .A(n528), .ZN(n667) );
  XNOR2_X1 U626 ( .A(n596), .B(KEYINPUT38), .ZN(n665) );
  NOR2_X1 U627 ( .A1(n665), .A2(n664), .ZN(n663) );
  NAND2_X1 U628 ( .A1(n667), .A2(n663), .ZN(n530) );
  XNOR2_X1 U629 ( .A(n531), .B(n530), .ZN(n676) );
  XOR2_X1 U630 ( .A(KEYINPUT105), .B(KEYINPUT28), .Z(n538) );
  NOR2_X1 U631 ( .A1(G900), .A2(n532), .ZN(n533) );
  NOR2_X1 U632 ( .A1(n534), .A2(n533), .ZN(n547) );
  NAND2_X1 U633 ( .A1(n535), .A2(n651), .ZN(n536) );
  NAND2_X1 U634 ( .A1(n564), .A2(n543), .ZN(n537) );
  XNOR2_X1 U635 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U636 ( .A1(n676), .A2(n559), .ZN(n541) );
  XNOR2_X1 U637 ( .A(n542), .B(n541), .ZN(n735) );
  XNOR2_X1 U638 ( .A(KEYINPUT30), .B(KEYINPUT104), .ZN(n545) );
  NAND2_X1 U639 ( .A1(n543), .A2(n591), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n545), .B(n544), .ZN(n546) );
  NOR2_X1 U641 ( .A1(n547), .A2(n546), .ZN(n550) );
  INV_X1 U642 ( .A(n548), .ZN(n549) );
  NAND2_X1 U643 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U644 ( .A(n551), .B(KEYINPUT72), .ZN(n578) );
  NOR2_X1 U645 ( .A1(n578), .A2(n665), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n552), .B(KEYINPUT39), .ZN(n590) );
  NOR2_X1 U647 ( .A1(n590), .A2(n553), .ZN(n555) );
  NOR2_X1 U648 ( .A1(n735), .A2(n733), .ZN(n558) );
  INV_X1 U649 ( .A(KEYINPUT78), .ZN(n556) );
  XNOR2_X1 U650 ( .A(n558), .B(n557), .ZN(n587) );
  INV_X1 U651 ( .A(n559), .ZN(n561) );
  XOR2_X1 U652 ( .A(KEYINPUT47), .B(n633), .Z(n563) );
  NAND2_X1 U653 ( .A1(n633), .A2(n580), .ZN(n562) );
  NAND2_X1 U654 ( .A1(n563), .A2(n562), .ZN(n576) );
  INV_X1 U655 ( .A(n502), .ZN(n575) );
  INV_X1 U656 ( .A(n564), .ZN(n566) );
  XNOR2_X1 U657 ( .A(KEYINPUT102), .B(n567), .ZN(n568) );
  INV_X1 U658 ( .A(n570), .ZN(n571) );
  NAND2_X1 U659 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n575), .A2(n349), .ZN(n641) );
  NAND2_X1 U661 ( .A1(n576), .A2(n641), .ZN(n584) );
  NOR2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U663 ( .A1(n596), .A2(n579), .ZN(n619) );
  NAND2_X1 U664 ( .A1(n580), .A2(KEYINPUT47), .ZN(n581) );
  NAND2_X1 U665 ( .A1(n619), .A2(n581), .ZN(n582) );
  XNOR2_X1 U666 ( .A(n582), .B(KEYINPUT76), .ZN(n583) );
  XNOR2_X1 U667 ( .A(n585), .B(KEYINPUT69), .ZN(n586) );
  XNOR2_X1 U668 ( .A(n588), .B(KEYINPUT48), .ZN(n600) );
  OR2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n644) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U671 ( .A(n593), .B(KEYINPUT103), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(n502), .ZN(n595) );
  XNOR2_X1 U673 ( .A(n595), .B(KEYINPUT43), .ZN(n598) );
  INV_X1 U674 ( .A(n596), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n620) );
  AND2_X1 U676 ( .A1(n644), .A2(n620), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n602), .B(KEYINPUT77), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(KEYINPUT2), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n691), .A2(G210), .ZN(n609) );
  XOR2_X1 U680 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n606) );
  XNOR2_X1 U681 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n611) );
  INV_X1 U683 ( .A(G952), .ZN(n610) );
  AND2_X1 U684 ( .A1(n610), .A2(G953), .ZN(n706) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U686 ( .A1(n691), .A2(G472), .ZN(n615) );
  XNOR2_X1 U687 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U689 ( .A(n618), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U690 ( .A(n619), .B(G143), .ZN(G45) );
  XNOR2_X1 U691 ( .A(n620), .B(G140), .ZN(G42) );
  XNOR2_X1 U692 ( .A(n621), .B(G119), .ZN(G21) );
  XNOR2_X1 U693 ( .A(G101), .B(n622), .ZN(G3) );
  NAND2_X1 U694 ( .A1(n627), .A2(n635), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n623), .B(G104), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n625) );
  XNOR2_X1 U697 ( .A(G107), .B(KEYINPUT26), .ZN(n624) );
  XNOR2_X1 U698 ( .A(n625), .B(n624), .ZN(n626) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(n626), .Z(n629) );
  NAND2_X1 U700 ( .A1(n627), .A2(n639), .ZN(n628) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(G9) );
  XNOR2_X1 U702 ( .A(G110), .B(n630), .ZN(G12) );
  XOR2_X1 U703 ( .A(G128), .B(KEYINPUT29), .Z(n632) );
  NAND2_X1 U704 ( .A1(n633), .A2(n639), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(G30) );
  NAND2_X1 U706 ( .A1(n633), .A2(n635), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n638), .A2(n635), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT114), .ZN(n637) );
  XNOR2_X1 U710 ( .A(G113), .B(n637), .ZN(G15) );
  NAND2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(G116), .ZN(G18) );
  XNOR2_X1 U713 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(G125), .B(n643), .ZN(G27) );
  INV_X1 U716 ( .A(n644), .ZN(n645) );
  XOR2_X1 U717 ( .A(G134), .B(n645), .Z(G36) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n659) );
  XOR2_X1 U719 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n650) );
  NAND2_X1 U720 ( .A1(n502), .A2(n648), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n655) );
  NOR2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U723 ( .A(KEYINPUT49), .B(n653), .Z(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U727 ( .A(KEYINPUT51), .B(n660), .Z(n661) );
  NAND2_X1 U728 ( .A1(n676), .A2(n661), .ZN(n672) );
  NAND2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U733 ( .A1(n677), .A2(n670), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U735 ( .A(KEYINPUT52), .B(n673), .Z(n674) );
  NOR2_X1 U736 ( .A1(n675), .A2(n674), .ZN(n679) );
  AND2_X1 U737 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U738 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n680), .B(KEYINPUT117), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n681), .A2(G953), .ZN(n682) );
  NAND2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U742 ( .A(KEYINPUT118), .B(n684), .ZN(n685) );
  XOR2_X1 U743 ( .A(KEYINPUT53), .B(n685), .Z(G75) );
  NAND2_X1 U744 ( .A1(n702), .A2(G469), .ZN(n689) );
  XOR2_X1 U745 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n686) );
  NOR2_X1 U746 ( .A1(n706), .A2(n690), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n691), .A2(G475), .ZN(n694) );
  XOR2_X1 U748 ( .A(n692), .B(KEYINPUT59), .Z(n693) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U750 ( .A(KEYINPUT60), .B(KEYINPUT65), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n696), .B(KEYINPUT119), .ZN(n697) );
  XNOR2_X1 U752 ( .A(n698), .B(n697), .ZN(G60) );
  NAND2_X1 U753 ( .A1(n702), .A2(G478), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n706), .A2(n701), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n702), .A2(G217), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  NAND2_X1 U759 ( .A1(G953), .A2(G224), .ZN(n707) );
  XNOR2_X1 U760 ( .A(KEYINPUT61), .B(n707), .ZN(n708) );
  NAND2_X1 U761 ( .A1(n708), .A2(G898), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT120), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n710), .A2(n728), .ZN(n711) );
  XOR2_X1 U764 ( .A(KEYINPUT121), .B(n711), .Z(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n720) );
  XNOR2_X1 U766 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n714) );
  XNOR2_X1 U767 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n716), .B(G101), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n728), .A2(G898), .ZN(n717) );
  NOR2_X1 U770 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n720), .B(n719), .ZN(G69) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n723), .B(KEYINPUT124), .ZN(n726) );
  XNOR2_X1 U774 ( .A(n726), .B(n724), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(n728), .ZN(n731) );
  XOR2_X1 U776 ( .A(G227), .B(n726), .Z(n727) );
  NOR2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U778 ( .A1(G900), .A2(n729), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT125), .B(n732), .ZN(G72) );
  XOR2_X1 U781 ( .A(n733), .B(G131), .Z(G33) );
  XNOR2_X1 U782 ( .A(G122), .B(n734), .ZN(G24) );
  XOR2_X1 U783 ( .A(G137), .B(n735), .Z(n736) );
  XNOR2_X1 U784 ( .A(KEYINPUT126), .B(n736), .ZN(G39) );
endmodule

