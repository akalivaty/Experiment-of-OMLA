//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(KEYINPUT79), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT79), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(G125), .A3(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT80), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(new_n190), .A3(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(new_n196), .ZN(new_n201));
  OR3_X1    g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n200), .B1(new_n199), .B2(new_n201), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT72), .B(G237), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(G214), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(KEYINPUT95), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(KEYINPUT95), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n208), .B1(new_n212), .B2(new_n210), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n217), .A3(new_n213), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n211), .B2(new_n213), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT98), .B1(new_n220), .B2(KEYINPUT17), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(KEYINPUT98), .A3(KEYINPUT17), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n205), .B(new_n219), .C1(new_n221), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n211), .B(new_n213), .C1(new_n225), .C2(new_n217), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n192), .A2(G146), .A3(new_n194), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT65), .B(G146), .ZN(new_n228));
  XNOR2_X1  g042(.A(G125), .B(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n226), .B(new_n231), .C1(new_n215), .C2(new_n225), .ZN(new_n232));
  XNOR2_X1  g046(.A(G113), .B(G122), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT97), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n224), .B2(new_n232), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n188), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G475), .ZN(new_n241));
  XNOR2_X1  g055(.A(G116), .B(G122), .ZN(new_n242));
  INV_X1    g056(.A(G107), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT100), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(G128), .B(G143), .Z(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(G134), .ZN(new_n248));
  INV_X1    g062(.A(G116), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT14), .A3(G122), .ZN(new_n250));
  INV_X1    g064(.A(new_n242), .ZN(new_n251));
  OAI211_X1 g065(.A(G107), .B(new_n250), .C1(new_n251), .C2(KEYINPUT14), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT99), .B(KEYINPUT13), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(G128), .A3(new_n209), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(G134), .C1(new_n247), .C2(new_n254), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n242), .B(new_n243), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(new_n257), .C1(G134), .C2(new_n247), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT9), .B(G234), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(G217), .A3(new_n207), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n253), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n253), .B2(new_n258), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT101), .B1(new_n265), .B2(G902), .ZN(new_n266));
  INV_X1    g080(.A(G478), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT15), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT101), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(new_n188), .C1(new_n263), .C2(new_n264), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  OR3_X1    g085(.A1(new_n265), .A2(G902), .A3(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(G234), .A2(G237), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n274), .A2(G952), .A3(new_n207), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT21), .B(G898), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT102), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n274), .A2(G902), .A3(G953), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n192), .A2(KEYINPUT19), .A3(new_n194), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT19), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n283), .B2(new_n229), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n228), .ZN(new_n285));
  INV_X1    g099(.A(new_n218), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n202), .B(new_n285), .C1(new_n286), .C2(new_n220), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n235), .B1(new_n287), .B2(new_n232), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT96), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI211_X1 g104(.A(KEYINPUT96), .B(new_n235), .C1(new_n287), .C2(new_n232), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n237), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT20), .ZN(new_n293));
  NOR2_X1   g107(.A1(G475), .A2(G902), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n292), .B2(new_n294), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n241), .B(new_n281), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n234), .A2(G107), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n234), .A2(G107), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT82), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n243), .A2(G104), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G101), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n306), .A2(KEYINPUT82), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n311), .B2(new_n308), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n301), .A2(new_n302), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n305), .A4(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(KEYINPUT4), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n249), .A2(G119), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n322), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n320), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(G101), .C1(new_n304), .C2(new_n309), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n316), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(KEYINPUT5), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n318), .A2(KEYINPUT5), .ZN(new_n331));
  INV_X1    g145(.A(G113), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT83), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n243), .B2(G104), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n308), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n305), .A2(new_n335), .ZN(new_n338));
  OAI21_X1  g152(.A(G101), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n334), .A2(new_n325), .A3(new_n315), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n329), .A2(new_n340), .A3(KEYINPUT88), .ZN(new_n345));
  XNOR2_X1  g159(.A(G110), .B(G122), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n344), .A3(new_n345), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT90), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n346), .B1(new_n341), .B2(new_n342), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n344), .A4(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G128), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(KEYINPUT1), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT66), .B1(new_n200), .B2(G143), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n228), .B2(G143), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n200), .A2(KEYINPUT65), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G146), .ZN(new_n361));
  AND4_X1   g175(.A1(new_n358), .A2(new_n359), .A3(new_n361), .A4(G143), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n355), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n359), .A2(new_n361), .A3(G143), .ZN(new_n366));
  INV_X1    g180(.A(new_n356), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n359), .A2(new_n361), .A3(new_n358), .A4(G143), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT70), .A3(new_n355), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n200), .A2(G143), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n228), .B2(G143), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(KEYINPUT1), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G128), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n365), .A2(new_n371), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n191), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n207), .A2(G224), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT91), .ZN(new_n379));
  AND2_X1   g193(.A1(KEYINPUT0), .A2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n377), .A2(new_n379), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n379), .B1(new_n377), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n329), .A2(new_n340), .A3(new_n346), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n391), .A2(KEYINPUT6), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT89), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n390), .A2(KEYINPUT89), .A3(new_n392), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n353), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n340), .A2(KEYINPUT92), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n340), .A2(KEYINPUT92), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n334), .A2(new_n325), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n315), .A2(new_n339), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n346), .B(KEYINPUT8), .Z(new_n402));
  OAI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n379), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n377), .B2(new_n386), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n377), .A2(new_n386), .A3(new_n405), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n395), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n395), .A2(new_n409), .A3(new_n411), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT93), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n416), .A3(new_n412), .ZN(new_n417));
  AND4_X1   g231(.A1(new_n187), .A2(new_n299), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n207), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n399), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT84), .B1(new_n376), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n375), .A2(new_n373), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT70), .B1(new_n370), .B2(new_n355), .ZN(new_n429));
  INV_X1    g243(.A(new_n355), .ZN(new_n430));
  AOI211_X1 g244(.A(new_n364), .B(new_n430), .C1(new_n368), .C2(new_n369), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n425), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT67), .ZN(new_n436));
  INV_X1    g250(.A(G134), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(G137), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT11), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n436), .B(new_n440), .C1(new_n437), .C2(G137), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n437), .A2(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n439), .A2(new_n217), .A3(new_n441), .A4(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n316), .A2(new_n328), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n385), .ZN(new_n449));
  INV_X1    g263(.A(new_n370), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n372), .A2(KEYINPUT1), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n429), .B2(new_n431), .ZN(new_n454));
  INV_X1    g268(.A(new_n399), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n456), .B2(new_n424), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n435), .A2(new_n447), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n447), .B1(new_n435), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n423), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n435), .A2(new_n457), .A3(new_n447), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n428), .B(new_n399), .C1(new_n429), .C2(new_n431), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n365), .A2(new_n371), .B1(new_n450), .B2(new_n452), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n399), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n446), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT12), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n467), .A3(new_n446), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n461), .A2(new_n466), .A3(new_n422), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n188), .A3(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(G469), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n461), .A2(new_n466), .A3(new_n423), .A4(new_n468), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n376), .A2(new_n426), .A3(KEYINPUT84), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n433), .B1(new_n432), .B2(new_n425), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n365), .A2(new_n371), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n399), .B1(new_n476), .B2(new_n453), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n477), .A2(KEYINPUT10), .B1(new_n448), .B2(new_n385), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n446), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n423), .B1(new_n479), .B2(new_n461), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n472), .B1(new_n480), .B2(KEYINPUT86), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n472), .A2(KEYINPUT86), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT85), .B(G469), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n471), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G221), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(new_n260), .B2(new_n188), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n419), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n422), .B1(new_n458), .B2(new_n459), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n482), .B1(new_n494), .B2(new_n472), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n495), .A2(G902), .A3(new_n485), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT87), .B(new_n491), .C1(new_n496), .C2(new_n471), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n418), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT103), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G234), .ZN(new_n501));
  OAI21_X1  g315(.A(G217), .B1(new_n501), .B2(G902), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT77), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n317), .A2(G128), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n354), .A2(KEYINPUT23), .A3(G119), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n317), .A2(G128), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n504), .B(new_n505), .C1(new_n506), .C2(KEYINPUT23), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G110), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(KEYINPUT78), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n504), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n204), .B(new_n508), .C1(new_n509), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n507), .A2(G110), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n512), .A2(new_n509), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n202), .B(new_n230), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT22), .B(G137), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n488), .A2(new_n501), .A3(G953), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n518), .B(new_n519), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n516), .A3(new_n520), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n188), .A3(new_n523), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n503), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n502), .A2(new_n188), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT81), .Z(new_n531));
  AND2_X1   g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n437), .B2(G137), .ZN(new_n537));
  INV_X1    g351(.A(G137), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT68), .A3(G134), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n442), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n540), .B2(G131), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n445), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n540), .A2(new_n535), .A3(G131), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT71), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n432), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n326), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n446), .A2(new_n381), .A3(new_n384), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT75), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n551), .A2(KEYINPUT75), .A3(new_n552), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n548), .A2(new_n550), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n326), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n551), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n557), .B1(KEYINPUT28), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n206), .A2(G210), .A3(new_n207), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT27), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT26), .B(G101), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(KEYINPUT29), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n561), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n544), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n445), .B2(new_n541), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n550), .B1(new_n376), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n548), .A2(KEYINPUT30), .A3(new_n550), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n326), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n551), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n565), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n569), .B1(new_n476), .B2(new_n428), .ZN(new_n578));
  INV_X1    g392(.A(new_n550), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n577), .B(new_n326), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n551), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n570), .B2(new_n326), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT28), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  INV_X1    g400(.A(new_n556), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT75), .B1(new_n551), .B2(new_n552), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n576), .B1(new_n590), .B2(new_n565), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n567), .B1(new_n591), .B2(KEYINPUT29), .ZN(new_n592));
  NOR2_X1   g406(.A1(G472), .A2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n565), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT31), .B1(new_n575), .B2(new_n595), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT31), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n574), .A2(new_n598), .A3(new_n565), .A4(new_n551), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n594), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n592), .A2(G472), .B1(new_n602), .B2(KEYINPUT32), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n590), .B2(new_n595), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT76), .B1(new_n604), .B2(new_n594), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT76), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n557), .B1(new_n584), .B2(new_n583), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n565), .B1(new_n607), .B2(new_n586), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n606), .B(new_n593), .C1(new_n608), .C2(new_n600), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT32), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n534), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n418), .A2(new_n490), .A3(KEYINPUT103), .A4(new_n497), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n500), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  OAI21_X1  g429(.A(G472), .B1(new_n604), .B2(G902), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n605), .A2(new_n616), .A3(new_n609), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n490), .A2(new_n497), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n534), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n265), .A2(KEYINPUT33), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT106), .Z(new_n622));
  NAND2_X1  g436(.A1(new_n265), .A2(KEYINPUT33), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(KEYINPUT107), .Z(new_n624));
  NAND4_X1  g438(.A1(new_n622), .A2(new_n624), .A3(G478), .A4(new_n188), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n241), .B1(new_n295), .B2(new_n297), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n395), .A2(new_n409), .A3(new_n411), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n411), .B1(new_n395), .B2(new_n409), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT104), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n395), .A2(new_n409), .A3(KEYINPUT104), .A4(new_n411), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n187), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n631), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n280), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n413), .A2(new_n639), .A3(new_n414), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(KEYINPUT105), .A3(new_n187), .A4(new_n635), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n637), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n620), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AND3_X1   g459(.A1(new_n292), .A2(new_n296), .A3(new_n294), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n241), .B(new_n273), .C1(new_n646), .C2(new_n297), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n637), .A2(new_n641), .A3(new_n638), .A4(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(KEYINPUT108), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(KEYINPUT108), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n620), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT109), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n517), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n531), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n529), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n617), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n500), .A2(new_n613), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AOI21_X1  g479(.A(new_n660), .B1(new_n603), .B2(new_n611), .ZN(new_n666));
  AND4_X1   g480(.A1(new_n461), .A2(new_n423), .A3(new_n466), .A4(new_n468), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n493), .B2(new_n492), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n188), .B(new_n486), .C1(new_n668), .C2(new_n482), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n470), .A2(G469), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n489), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(KEYINPUT87), .ZN(new_n672));
  AOI211_X1 g486(.A(new_n419), .B(new_n489), .C1(new_n669), .C2(new_n670), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n637), .A2(new_n641), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n275), .B1(new_n279), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n241), .B(new_n678), .C1(new_n646), .C2(new_n297), .ZN(new_n679));
  INV_X1    g493(.A(new_n273), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n666), .A2(new_n674), .A3(new_n675), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n415), .A2(new_n417), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT38), .ZN(new_n685));
  INV_X1    g499(.A(new_n187), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n628), .A2(new_n273), .ZN(new_n687));
  NOR4_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n661), .A4(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n560), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n595), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n575), .A2(new_n565), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n602), .A2(KEYINPUT32), .B1(G472), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n611), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n677), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n674), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n688), .B(new_n694), .C1(KEYINPUT40), .C2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(KEYINPUT40), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n209), .ZN(G45));
  NOR2_X1   g513(.A1(new_n629), .A2(new_n677), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n666), .A2(new_n674), .A3(new_n675), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  OAI21_X1  g516(.A(G469), .B1(new_n495), .B2(G902), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n491), .A3(new_n669), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n612), .A2(new_n642), .A3(new_n630), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  OAI211_X1 g521(.A(new_n612), .B(new_n704), .C1(new_n650), .C2(new_n651), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  AND3_X1   g523(.A1(new_n704), .A2(new_n637), .A3(new_n641), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n666), .A2(new_n710), .A3(new_n299), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND2_X1  g526(.A1(new_n637), .A2(new_n641), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n687), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n561), .A2(new_n565), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n593), .B1(new_n715), .B2(new_n600), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n616), .A2(new_n533), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n703), .A2(new_n491), .A3(new_n669), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n280), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n704), .A2(new_n637), .A3(new_n641), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n700), .A2(new_n616), .A3(new_n661), .A4(new_n716), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n191), .ZN(G27));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n686), .B1(new_n415), .B2(new_n417), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n700), .A2(new_n728), .A3(new_n671), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n612), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n610), .B1(new_n604), .B2(new_n594), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n534), .B1(new_n603), .B2(new_n731), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n732), .A2(new_n729), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n726), .B(new_n730), .C1(new_n733), .C2(new_n727), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n612), .A2(new_n727), .A3(new_n729), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n727), .B1(new_n732), .B2(new_n729), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT110), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n217), .ZN(G33));
  AND3_X1   g553(.A1(new_n728), .A2(new_n671), .A3(new_n681), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n603), .A2(new_n611), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n740), .A2(new_n741), .A3(new_n533), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n437), .ZN(G36));
  INV_X1    g557(.A(new_n627), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(KEYINPUT43), .A3(new_n628), .ZN(new_n745));
  INV_X1    g559(.A(new_n628), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT111), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n628), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n627), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n745), .B1(new_n750), .B2(KEYINPUT43), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n618), .A3(new_n661), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n728), .ZN(new_n755));
  INV_X1    g569(.A(G469), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n460), .A2(new_n469), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n757), .B2(KEYINPUT45), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(KEYINPUT45), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g573(.A1(G469), .A2(G902), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT46), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n496), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(KEYINPUT46), .A3(new_n760), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n489), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n695), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n754), .A2(new_n755), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n753), .B2(new_n752), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT112), .B(G137), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G39));
  XOR2_X1   g583(.A(new_n764), .B(KEYINPUT47), .Z(new_n770));
  AND2_X1   g584(.A1(new_n603), .A2(new_n611), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n534), .A3(new_n700), .A4(new_n728), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  AND3_X1   g588(.A1(new_n704), .A2(new_n275), .A3(new_n728), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n611), .A3(new_n533), .A4(new_n693), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT117), .Z(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n630), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n775), .A2(new_n751), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT48), .A4(new_n732), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n616), .A2(new_n716), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n751), .A2(new_n533), .A3(new_n275), .A4(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(G952), .B(new_n207), .C1(new_n783), .C2(new_n722), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n732), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n778), .A2(new_n781), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  INV_X1    g605(.A(new_n685), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n783), .A2(new_n792), .A3(new_n187), .A4(new_n718), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n782), .A2(new_n661), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(new_n779), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n777), .A2(new_n746), .A3(new_n744), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n703), .A2(new_n669), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT113), .Z(new_n801));
  OAI21_X1  g615(.A(new_n770), .B1(new_n491), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n783), .A2(new_n755), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT51), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n790), .B(new_n791), .C1(new_n799), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n797), .A2(KEYINPUT118), .A3(new_n798), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(new_n804), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n705), .A2(new_n711), .A3(new_n720), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n782), .A2(new_n671), .A3(new_n700), .A4(new_n728), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n679), .A2(new_n273), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n490), .A2(new_n497), .A3(new_n728), .A4(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n771), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n742), .B1(new_n817), .B2(new_n661), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n818), .A3(new_n708), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n738), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n722), .A2(new_n723), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n529), .A2(new_n659), .A3(new_n677), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n671), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n611), .B2(new_n693), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n714), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n682), .A2(new_n701), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(new_n681), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n619), .A2(new_n713), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n724), .B1(new_n829), .B2(new_n666), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n701), .A4(new_n825), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n629), .B1(new_n628), .B2(new_n680), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n638), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n835), .A2(new_n686), .A3(new_n684), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n533), .A3(new_n674), .A4(new_n617), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n614), .A2(new_n837), .A3(new_n663), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n614), .A2(new_n837), .A3(new_n663), .A4(KEYINPUT114), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n833), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n830), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT53), .B1(new_n846), .B2(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n735), .A2(new_n736), .A3(new_n844), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n831), .B2(new_n830), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n819), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n833), .A3(new_n842), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n833), .A4(new_n842), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n860), .A3(new_n844), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n812), .A2(new_n849), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n801), .B(KEYINPUT49), .ZN(new_n865));
  OR4_X1    g679(.A1(new_n534), .A2(new_n750), .A3(new_n489), .A4(new_n686), .ZN(new_n866));
  OR4_X1    g680(.A1(new_n694), .A2(new_n865), .A3(new_n792), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(G75));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(G210), .A3(G902), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n353), .B1(new_n393), .B2(new_n394), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n389), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n207), .A2(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G51));
  XOR2_X1   g692(.A(new_n760), .B(KEYINPUT57), .Z(new_n879));
  AND3_X1   g693(.A1(new_n843), .A2(new_n860), .A3(new_n844), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n860), .B1(new_n843), .B2(new_n844), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n859), .B1(new_n882), .B2(new_n857), .ZN(new_n883));
  INV_X1    g697(.A(new_n862), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n495), .B(KEYINPUT121), .Z(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n869), .A2(G902), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(new_n759), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n877), .B1(new_n887), .B2(new_n889), .ZN(G54));
  NAND4_X1  g704(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n892));
  INV_X1    g706(.A(new_n292), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n877), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n891), .B2(new_n893), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n862), .B2(new_n849), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n622), .A2(new_n624), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n900), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n883), .B2(new_n884), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT123), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n905), .C1(new_n883), .C2(new_n884), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT124), .Z(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT60), .Z(new_n913));
  NAND2_X1  g727(.A1(new_n869), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n524), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n882), .B2(new_n857), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n877), .B1(new_n918), .B2(new_n657), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT125), .B1(new_n918), .B2(new_n657), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n916), .B(new_n919), .C1(new_n920), .C2(KEYINPUT61), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n869), .A2(new_n657), .A3(new_n913), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(new_n895), .C1(new_n918), .C2(new_n524), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT61), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n278), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n813), .A2(new_n708), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n842), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(KEYINPUT126), .A3(new_n207), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT126), .B1(new_n931), .B2(new_n207), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n872), .B1(G898), .B2(new_n207), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  NAND4_X1  g750(.A1(new_n764), .A2(new_n714), .A3(new_n695), .A4(new_n732), .ZN(new_n937));
  INV_X1    g751(.A(new_n742), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n767), .A2(new_n773), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n830), .A2(new_n701), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n738), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n941), .A2(new_n945), .A3(new_n942), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n207), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n572), .A2(new_n573), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n284), .Z(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(G900), .B2(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n698), .A2(KEYINPUT62), .A3(new_n940), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n834), .A2(new_n728), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n612), .A2(new_n674), .A3(new_n695), .A4(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n767), .A2(new_n773), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT62), .B1(new_n698), .B2(new_n940), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n950), .B1(new_n958), .B2(G953), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n952), .A2(new_n963), .A3(new_n959), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G72));
  INV_X1    g779(.A(new_n576), .ZN(new_n966));
  INV_X1    g780(.A(new_n931), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n944), .A2(new_n967), .A3(new_n946), .ZN(new_n968));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  AOI21_X1  g784(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n970), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n958), .B2(new_n967), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n895), .B1(new_n973), .B2(new_n691), .ZN(new_n974));
  AND4_X1   g788(.A1(new_n966), .A2(new_n848), .A3(new_n691), .A4(new_n970), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(G57));
endmodule


