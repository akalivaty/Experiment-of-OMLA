//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT1), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n205));
  INV_X1    g0005(.A(G50), .ZN(new_n206));
  INV_X1    g0006(.A(G226), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI221_X1 g0009(.A(new_n205), .B1(new_n206), .B2(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT66), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g0012(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n212), .B(new_n213), .C1(G107), .C2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n203), .B1(KEYINPUT67), .B2(new_n204), .C1(new_n219), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n203), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n221), .B(new_n227), .C1(new_n218), .C2(new_n228), .ZN(new_n229));
  OR2_X1    g0029(.A1(KEYINPUT64), .A2(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(KEYINPUT64), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(G68), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n215), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  OAI22_X1  g0038(.A1(new_n229), .A2(KEYINPUT0), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT0), .B2(new_n229), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT65), .Z(new_n241));
  NOR2_X1   g0041(.A1(new_n225), .A2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G264), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n209), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT73), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT73), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G1698), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n262), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT76), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G87), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n262), .A2(G226), .A3(G1698), .A4(new_n264), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n264), .A4(new_n266), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n233), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT69), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n277), .A2(KEYINPUT69), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n274), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G232), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n275), .A2(new_n284), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT77), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n275), .A2(KEYINPUT77), .A3(new_n284), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g0099(.A(KEYINPUT8), .B(G58), .Z(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT75), .Z(new_n303));
  NAND3_X1  g0103(.A1(new_n276), .A2(G13), .A3(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n233), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n304), .B2(new_n300), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT3), .B1(new_n259), .B2(new_n261), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(KEYINPUT7), .B(new_n232), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT3), .B(G33), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n316), .B1(new_n317), .B2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(KEYINPUT74), .B1(new_n319), .B2(G68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  AOI211_X1 g0121(.A(new_n321), .B(new_n236), .C1(new_n315), .C2(new_n318), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(G58), .B(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(G20), .B1(G159), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT16), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n264), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT73), .B(G33), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n328), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT7), .B1(new_n330), .B2(G20), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n262), .A2(new_n264), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n316), .A3(new_n232), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(G68), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n326), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n307), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n311), .B1(new_n327), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n293), .A2(G179), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n299), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n299), .A2(new_n338), .A3(KEYINPUT18), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n319), .A2(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n321), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n319), .A2(KEYINPUT74), .A3(G68), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n347), .A2(new_n326), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n336), .ZN(new_n350));
  INV_X1    g0150(.A(new_n307), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n334), .A2(new_n326), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(KEYINPUT16), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n310), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(G200), .B1(new_n295), .B2(new_n296), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n293), .A2(G190), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT17), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n297), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n356), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n338), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT17), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n345), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n282), .A2(new_n283), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G97), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n264), .A2(new_n313), .ZN(new_n369));
  INV_X1    g0169(.A(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n207), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n216), .A2(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n368), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n367), .A2(new_n278), .B1(new_n374), .B2(new_n274), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n291), .A2(G238), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n366), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n274), .ZN(new_n378));
  AND4_X1   g0178(.A1(new_n366), .A2(new_n376), .A3(new_n378), .A4(new_n284), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n377), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(G169), .C1(new_n377), .C2(new_n379), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n325), .A2(G50), .B1(G20), .B2(new_n236), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n232), .A2(G33), .ZN(new_n389));
  INV_X1    g0189(.A(G77), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n307), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT11), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n276), .A2(new_n236), .A3(G13), .A4(G20), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT12), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n351), .A2(new_n301), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G68), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT71), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n381), .A2(new_n383), .A3(new_n401), .A4(new_n385), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n387), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n400), .B1(G190), .B2(new_n382), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n360), .B2(new_n382), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n291), .A2(G244), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n284), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G238), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n317), .B(new_n409), .C1(new_n216), .C2(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n274), .C1(G107), .C2(new_n317), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT70), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n406), .A2(new_n412), .A3(new_n284), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n408), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n414), .A2(G179), .ZN(new_n415));
  AND2_X1   g0215(.A1(KEYINPUT64), .A2(G20), .ZN(new_n416));
  NOR2_X1   g0216(.A1(KEYINPUT64), .A2(G20), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n300), .A2(new_n325), .B1(new_n418), .B2(G77), .ZN(new_n419));
  XOR2_X1   g0219(.A(KEYINPUT15), .B(G87), .Z(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n389), .B2(new_n421), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n307), .B1(G77), .B2(new_n397), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n305), .A2(new_n390), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n414), .A2(new_n298), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n415), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n414), .A2(G200), .ZN(new_n428));
  INV_X1    g0228(.A(new_n425), .ZN(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n428), .B(new_n429), .C1(new_n430), .C2(new_n414), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n403), .A2(new_n405), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n370), .A2(G222), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n317), .B(new_n433), .C1(new_n265), .C2(new_n370), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n274), .C1(G77), .C2(new_n317), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n291), .A2(G226), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n284), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(G179), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n325), .A2(G150), .ZN(new_n439));
  OAI21_X1  g0239(.A(G20), .B1(new_n237), .B2(G50), .ZN(new_n440));
  XNOR2_X1  g0240(.A(KEYINPUT8), .B(G58), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n439), .B(new_n440), .C1(new_n389), .C2(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n307), .B1(G50), .B2(new_n397), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G50), .B2(new_n304), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n437), .A2(new_n298), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n438), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n437), .A2(G200), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT9), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n447), .B1(new_n430), .B2(new_n437), .C1(new_n444), .C2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n444), .A2(new_n448), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n451), .A2(KEYINPUT10), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(KEYINPUT10), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n446), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n365), .A2(new_n432), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n286), .A2(G1), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G274), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n457), .B(new_n458), .ZN(new_n459));
  OR3_X1    g0259(.A1(new_n274), .A2(new_n221), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n208), .B1(new_n259), .B2(new_n261), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n370), .A2(G238), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n330), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT82), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n330), .A2(new_n465), .A3(G244), .A4(G1698), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n262), .A2(G244), .A3(G1698), .A4(new_n264), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT82), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n461), .B1(new_n469), .B2(new_n274), .ZN(new_n470));
  INV_X1    g0270(.A(G179), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g0273(.A(G33), .B(G97), .C1(new_n416), .C2(new_n417), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n416), .A2(new_n417), .B1(new_n473), .B2(new_n368), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n220), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n473), .A2(new_n474), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n262), .A2(new_n232), .A3(G68), .A4(new_n264), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n307), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n421), .A2(new_n305), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n276), .A2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n308), .A2(new_n420), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n480), .A2(new_n307), .B1(new_n305), .B2(new_n421), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n484), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n472), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n470), .A2(G169), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n470), .A2(G190), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n351), .A2(new_n304), .A3(new_n483), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n220), .ZN(new_n494));
  XNOR2_X1  g0294(.A(new_n494), .B(KEYINPUT84), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n488), .B(new_n495), .C1(new_n470), .C2(new_n360), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n258), .A2(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n416), .C2(new_n417), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n306), .A2(new_n233), .B1(G20), .B2(new_n208), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT20), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n305), .A2(new_n208), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n493), .B2(new_n208), .ZN(new_n507));
  OAI21_X1  g0307(.A(G169), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n274), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n218), .A2(new_n370), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n228), .A2(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n262), .A2(new_n264), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n369), .A2(G303), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT5), .B(G41), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n456), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n509), .A3(G270), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n282), .A2(new_n456), .A3(new_n515), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n498), .B1(new_n508), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n514), .A2(new_n519), .ZN(new_n522));
  OAI221_X1 g0322(.A(new_n506), .B1(new_n208), .B2(new_n493), .C1(new_n503), .C2(new_n504), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n522), .A2(KEYINPUT21), .A3(G169), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n520), .A3(G179), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n520), .A2(G190), .ZN(new_n528));
  INV_X1    g0328(.A(new_n523), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(new_n360), .C2(new_n520), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n521), .A3(new_n524), .A4(new_n525), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT85), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n497), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT23), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n230), .A2(new_n535), .A3(new_n536), .A4(new_n231), .ZN(new_n537));
  NAND2_X1  g0337(.A1(KEYINPUT23), .A2(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G20), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n462), .B2(KEYINPUT23), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n220), .B1(new_n230), .B2(new_n231), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n543), .A2(new_n262), .A3(KEYINPUT22), .A4(new_n264), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  OAI21_X1  g0345(.A(G87), .B1(new_n416), .B2(new_n417), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n369), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n540), .A2(new_n542), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT24), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT22), .B1(new_n543), .B2(new_n317), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(new_n539), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n552), .A2(KEYINPUT24), .A3(new_n542), .A4(new_n544), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n550), .A2(new_n553), .A3(new_n307), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n304), .A2(G107), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n555), .A2(KEYINPUT25), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT86), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n555), .B2(KEYINPUT25), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n558), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n493), .A2(new_n536), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n221), .A2(new_n370), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n218), .A2(G1698), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n262), .A2(new_n264), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n329), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n274), .B1(new_n456), .B2(new_n515), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(new_n274), .B1(G264), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n571), .A2(new_n518), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n471), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n518), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n298), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n563), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n264), .A2(new_n313), .A3(G250), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n370), .B1(new_n577), .B2(KEYINPUT4), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G1698), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(new_n264), .A3(new_n313), .A4(G244), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n500), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(G244), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n579), .B1(new_n332), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n509), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n570), .A2(G257), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n518), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n360), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n579), .B1(new_n317), .B2(G250), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n500), .B(new_n581), .C1(new_n590), .C2(new_n370), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT4), .B1(new_n330), .B2(G244), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n274), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n587), .A2(new_n518), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n430), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n305), .A2(new_n217), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n493), .B2(new_n217), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n319), .A2(G107), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT78), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(KEYINPUT6), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n603));
  OAI211_X1 g0403(.A(G97), .B(new_n536), .C1(new_n601), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n536), .A2(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(KEYINPUT78), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(KEYINPUT6), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n217), .A2(G107), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n418), .B1(G77), .B2(new_n325), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n599), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n598), .B1(new_n612), .B2(new_n307), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n596), .A2(KEYINPUT79), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT79), .B1(new_n596), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n571), .A2(G190), .A3(new_n518), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n554), .A2(new_n562), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n574), .A2(G200), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT80), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n298), .B1(new_n586), .B2(new_n588), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n593), .A2(new_n471), .A3(new_n594), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n624), .B2(new_n613), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n325), .A2(G77), .ZN(new_n626));
  INV_X1    g0426(.A(new_n610), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n232), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n536), .B1(new_n315), .B2(new_n318), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n307), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n598), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n632), .A2(KEYINPUT80), .A3(new_n623), .A4(new_n622), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n576), .A2(new_n616), .A3(new_n620), .A4(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n455), .A2(new_n534), .A3(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n446), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n364), .A2(new_n359), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n427), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n415), .A2(KEYINPUT90), .A3(new_n425), .A4(new_n426), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n405), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n403), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n345), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n452), .A2(new_n453), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n637), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n496), .A2(new_n492), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n469), .A2(new_n274), .ZN(new_n652));
  INV_X1    g0452(.A(new_n461), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n654), .B2(new_n298), .ZN(new_n655));
  NOR3_X1   g0455(.A1(new_n470), .A2(KEYINPUT87), .A3(G169), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n490), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n650), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n526), .A2(new_n576), .B1(new_n619), .B2(new_n618), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n634), .A3(new_n660), .A4(new_n616), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT89), .B1(new_n624), .B2(new_n613), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT89), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n632), .A2(new_n664), .A3(new_n623), .A4(new_n622), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n659), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT26), .B1(new_n497), .B2(new_n634), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n657), .A2(new_n658), .A3(KEYINPUT88), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n654), .A2(new_n651), .A3(new_n298), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT87), .B1(new_n470), .B2(G169), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n673), .B2(new_n490), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n661), .A2(new_n667), .A3(new_n668), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n455), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n649), .B1(new_n677), .B2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n418), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n276), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT91), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(G213), .A3(G343), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n576), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n563), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n620), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n689), .B2(new_n576), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n685), .A2(new_n529), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n531), .B2(new_n533), .ZN(new_n692));
  INV_X1    g0492(.A(new_n526), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT92), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n696), .A2(KEYINPUT92), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n690), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n686), .A2(new_n526), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n690), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n687), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(G399));
  NOR2_X1   g0504(.A1(new_n227), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n476), .A2(new_n220), .A3(new_n208), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n238), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n676), .A2(new_n685), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT95), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OR3_X1    g0513(.A1(new_n497), .A2(new_n634), .A3(KEYINPUT26), .ZN(new_n714));
  INV_X1    g0514(.A(new_n666), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n673), .A2(new_n490), .B1(new_n492), .B2(new_n496), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT26), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n661), .A3(new_n717), .A4(new_n675), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n718), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n713), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n718), .A2(KEYINPUT95), .A3(KEYINPUT29), .A4(new_n685), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n615), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n596), .A2(KEYINPUT79), .A3(new_n613), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n620), .A2(new_n634), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n534), .A3(new_n576), .A4(new_n685), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT94), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n586), .A2(new_n588), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n572), .A2(new_n728), .A3(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n654), .A3(new_n522), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n729), .A2(KEYINPUT93), .A3(new_n654), .A4(new_n522), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n522), .A2(new_n471), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(new_n728), .A3(new_n470), .A4(new_n571), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT30), .Z(new_n737));
  OAI21_X1  g0537(.A(new_n686), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT94), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n635), .A2(new_n741), .A3(new_n534), .A4(new_n685), .ZN(new_n742));
  INV_X1    g0542(.A(new_n730), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT31), .B(new_n686), .C1(new_n737), .C2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n727), .A2(new_n740), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n722), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n710), .B1(new_n747), .B2(G1), .ZN(G364));
  NOR2_X1   g0548(.A1(new_n698), .A2(new_n699), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n681), .A2(G45), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n707), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n694), .B2(new_n695), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n694), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n317), .A2(G355), .A3(new_n226), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n253), .A2(new_n286), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n330), .A2(new_n227), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n238), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n759), .B1(G116), .B2(new_n226), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n233), .B1(G20), .B2(new_n298), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n430), .A2(new_n360), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n767), .A2(G20), .A3(new_n471), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n220), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n232), .A2(G190), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n471), .A3(new_n360), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT32), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n232), .A2(new_n471), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n430), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G200), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n769), .B(new_n774), .C1(G77), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n767), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G50), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n770), .A2(new_n471), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G107), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n430), .A2(G200), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n775), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n775), .A2(new_n430), .A3(G200), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n215), .B1(new_n236), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n471), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n418), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n217), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n789), .A2(new_n369), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n778), .A2(new_n781), .A3(new_n784), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n779), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n772), .A2(G329), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT33), .B(G317), .Z(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n567), .B2(new_n792), .C1(new_n788), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G311), .B2(new_n777), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(G283), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n786), .A2(G322), .ZN(new_n803));
  INV_X1    g0603(.A(new_n768), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n317), .B1(new_n804), .B2(G303), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n795), .B1(new_n797), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n764), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n758), .A2(new_n766), .A3(new_n752), .A4(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n754), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(G396));
  NAND4_X1  g0611(.A1(new_n640), .A2(new_n425), .A3(new_n641), .A4(new_n686), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n427), .A2(new_n431), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n429), .B2(new_n685), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n676), .A2(new_n815), .A3(new_n685), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(KEYINPUT97), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n746), .B(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n815), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n711), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n818), .B(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n752), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n782), .A2(new_n220), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n787), .A2(new_n567), .B1(new_n825), .B2(new_n771), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n824), .B(new_n826), .C1(G116), .C2(new_n777), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n317), .B(new_n793), .C1(G107), .C2(new_n804), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  INV_X1    g0630(.A(G303), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(new_n830), .B2(new_n788), .C1(new_n831), .C2(new_n779), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n330), .B1(new_n768), .B2(new_n206), .C1(new_n792), .C2(new_n215), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n777), .A2(G159), .B1(G143), .B2(new_n786), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n779), .C1(new_n836), .C2(new_n788), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n772), .A2(G132), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n783), .A2(G68), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n832), .B1(new_n833), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n764), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n764), .A2(new_n755), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n752), .B1(G77), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT96), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n843), .B(new_n847), .C1(new_n756), .C2(new_n815), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n823), .A2(new_n848), .ZN(G384));
  NAND4_X1  g0649(.A1(new_n387), .A2(new_n400), .A3(new_n402), .A4(new_n686), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n686), .A2(new_n400), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n403), .A2(new_n405), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT100), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n850), .A2(new_n853), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n819), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT31), .B(new_n686), .C1(new_n734), .C2(new_n737), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n727), .A2(new_n740), .A3(new_n742), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n684), .A2(G213), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n338), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n341), .A2(new_n357), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  AOI21_X1  g0665(.A(G169), .B1(new_n295), .B2(new_n296), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n335), .A2(new_n336), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n310), .B1(new_n353), .B2(new_n867), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n866), .A2(new_n868), .A3(new_n339), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT101), .B1(new_n363), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n299), .A2(new_n340), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n357), .B(new_n871), .C1(new_n872), .C2(new_n868), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n861), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n865), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n638), .B2(new_n345), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n860), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n365), .A2(new_n874), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n357), .B1(new_n872), .B2(new_n868), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n882), .B2(KEYINPUT101), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n883), .B2(new_n873), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n880), .B(KEYINPUT38), .C1(new_n884), .C2(new_n865), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n859), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n863), .B1(new_n638), .B2(new_n345), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n864), .B(new_n881), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n860), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n859), .A2(KEYINPUT40), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n858), .A2(new_n455), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n895), .B(new_n896), .Z(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n403), .A2(new_n686), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n343), .A2(new_n344), .A3(new_n861), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n686), .A2(new_n427), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT99), .B1(new_n816), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n816), .A2(KEYINPUT99), .A3(new_n906), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n854), .A2(new_n855), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n910), .A2(new_n886), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n903), .A2(new_n904), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n721), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n713), .B2(new_n719), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n649), .B1(new_n915), .B2(new_n678), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n913), .B(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n898), .B(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n919));
  XNOR2_X1  g0719(.A(new_n918), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n276), .B2(new_n681), .ZN(new_n921));
  OAI21_X1  g0721(.A(G77), .B1(new_n215), .B2(new_n236), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n238), .A2(new_n922), .B1(G50), .B2(new_n236), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n680), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n208), .B1(new_n610), .B2(KEYINPUT35), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n925), .B(new_n234), .C1(KEYINPUT35), .C2(new_n610), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT98), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n924), .A3(new_n928), .ZN(G367));
  INV_X1    g0729(.A(new_n788), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n930), .A2(G159), .B1(new_n786), .B2(G150), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n780), .A2(G143), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n791), .A2(G68), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n777), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n317), .B1(new_n935), .B2(new_n206), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n782), .A2(new_n390), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n771), .A2(new_n835), .B1(new_n215), .B2(new_n768), .ZN(new_n938));
  NOR4_X1   g0738(.A1(new_n934), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n783), .A2(G97), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n536), .B2(new_n792), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT107), .B1(new_n804), .B2(G116), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT46), .ZN(new_n943));
  INV_X1    g0743(.A(G317), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n943), .B1(new_n825), .B2(new_n779), .C1(new_n944), .C2(new_n771), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n946), .B(new_n332), .C1(new_n830), .C2(new_n935), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n941), .B(new_n947), .C1(G294), .C2(new_n930), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n786), .A2(G303), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n939), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT47), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n764), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n685), .B1(new_n488), .B2(new_n495), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n669), .A3(new_n674), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n954), .B(new_n757), .C1(new_n716), .C2(new_n953), .ZN(new_n955));
  INV_X1    g0755(.A(new_n761), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n765), .B1(new_n226), .B2(new_n421), .C1(new_n249), .C2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n952), .A2(new_n752), .A3(new_n955), .A4(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n751), .A2(new_n276), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n616), .B(new_n634), .C1(new_n613), .C2(new_n685), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n685), .A2(new_n613), .A3(new_n624), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n702), .B2(new_n687), .ZN(new_n965));
  XOR2_X1   g0765(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n967), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT45), .B1(new_n703), .B2(new_n963), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT105), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n700), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n702), .A2(KEYINPUT106), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n749), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n749), .A2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n690), .B2(new_n701), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n690), .A2(new_n701), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n980), .A3(new_n977), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n747), .B1(new_n974), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n705), .B(KEYINPUT41), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n960), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n954), .B1(new_n716), .B2(new_n953), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n700), .A2(new_n964), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n702), .A2(new_n963), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT42), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n634), .B1(new_n964), .B2(new_n576), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n685), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n995), .A3(new_n994), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n987), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n998), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n987), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n1000), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n958), .B1(new_n985), .B2(new_n1004), .ZN(G387));
  NOR2_X1   g0805(.A1(new_n982), .A2(new_n959), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n441), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n708), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(G68), .A2(G77), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT50), .B1(new_n441), .B2(G50), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1008), .A2(new_n286), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n761), .B(new_n1011), .C1(new_n246), .C2(new_n286), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n317), .A2(new_n708), .A3(new_n226), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G107), .C2(new_n226), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT108), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n765), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G294), .A2(new_n804), .B1(new_n791), .B2(G283), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n777), .A2(G303), .B1(G317), .B2(new_n786), .ZN(new_n1018));
  INV_X1    g0818(.A(G322), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n825), .B2(new_n788), .C1(new_n1019), .C2(new_n779), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT48), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT109), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT49), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n332), .B1(new_n771), .B2(new_n796), .C1(new_n208), .C2(new_n782), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G159), .A2(new_n780), .B1(new_n786), .B2(G50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n791), .A2(new_n420), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(new_n236), .C2(new_n935), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G150), .B2(new_n772), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n804), .A2(G77), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n930), .A2(new_n300), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1034), .A2(new_n940), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n332), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n822), .B1(new_n1039), .B2(new_n764), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n690), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n757), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1006), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n747), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n706), .B1(new_n982), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n982), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(new_n1047), .ZN(G393));
  NOR2_X1   g0848(.A1(new_n982), .A2(new_n1045), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n700), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n973), .B(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n972), .A2(KEYINPUT112), .A3(new_n700), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n700), .A2(KEYINPUT112), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n972), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1052), .B(new_n705), .C1(new_n1049), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1053), .A2(KEYINPUT113), .A3(new_n1057), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(new_n960), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n822), .B1(new_n964), .B2(new_n757), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n765), .B1(new_n217), .B2(new_n226), .C1(new_n956), .C2(new_n256), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n787), .A2(new_n825), .B1(new_n944), .B2(new_n779), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT52), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n784), .C1(new_n831), .C2(new_n788), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n792), .A2(new_n208), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n935), .A2(new_n567), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n369), .B1(new_n830), .B2(new_n768), .C1(new_n771), .C2(new_n1019), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n935), .A2(new_n441), .ZN(new_n1073));
  INV_X1    g0873(.A(G159), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n787), .A2(new_n1074), .B1(new_n836), .B2(new_n779), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT51), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n930), .A2(G50), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n330), .B1(new_n236), .B2(new_n768), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G77), .B2(new_n791), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n824), .B1(G143), .B2(new_n772), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1073), .B(new_n1082), .C1(new_n1076), .C2(new_n1075), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n764), .B1(new_n1072), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1064), .A2(new_n1065), .A3(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1063), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1059), .A2(new_n1086), .ZN(G390));
  NAND3_X1  g0887(.A1(new_n856), .A2(G330), .A3(new_n858), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n816), .A2(KEYINPUT99), .A3(new_n906), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n911), .B1(new_n1089), .B2(new_n907), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n901), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n900), .A2(new_n902), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n718), .A2(new_n685), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n906), .B1(new_n1093), .B2(new_n819), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n911), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n893), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n745), .A2(G330), .A3(new_n815), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n911), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n879), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT39), .B1(new_n885), .B2(new_n892), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n901), .B1(new_n910), .B2(new_n911), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1096), .B(new_n1101), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n960), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n755), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n844), .A2(new_n441), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n840), .B1(new_n567), .B2(new_n771), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT116), .Z(new_n1112));
  NOR2_X1   g0912(.A1(new_n787), .A2(new_n208), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n769), .B1(G77), .B2(new_n791), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n830), .B2(new_n779), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n369), .B1(new_n536), .B2(new_n788), .C1(new_n935), .C2(new_n217), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n783), .A2(G50), .B1(new_n786), .B2(G132), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1118), .B1(new_n835), .B2(new_n788), .C1(new_n935), .C2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(G125), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n771), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n804), .A2(G150), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n317), .B1(new_n792), .B2(new_n1074), .C1(new_n779), .C2(new_n1126), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n764), .B1(new_n1117), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1109), .A2(new_n752), .A3(new_n1110), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1101), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1094), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n858), .A2(G330), .A3(new_n815), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n1100), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(new_n1088), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n910), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT115), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n858), .A2(G330), .A3(new_n455), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT114), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n858), .A2(new_n455), .A3(KEYINPUT114), .A4(G330), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1140), .B1(new_n1145), .B2(new_n916), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n722), .A2(new_n455), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1147), .A2(new_n1148), .A3(KEYINPUT115), .A4(new_n649), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1139), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n706), .B1(new_n1151), .B2(new_n1107), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1107), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1108), .B(new_n1130), .C1(new_n1153), .C2(new_n1154), .ZN(G378));
  NAND2_X1  g0955(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1107), .B2(new_n1139), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT119), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(KEYINPUT119), .B(new_n1156), .C1(new_n1107), .C2(new_n1139), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n856), .A2(new_n858), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n885), .B2(new_n879), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n894), .B(G330), .C1(new_n1162), .C2(KEYINPUT40), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  NOR2_X1   g0964(.A1(new_n454), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n454), .A2(new_n1164), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n444), .B2(new_n862), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n862), .A2(new_n444), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1169), .A2(new_n1170), .A3(new_n1165), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(KEYINPUT118), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n889), .A2(new_n1175), .A3(G330), .A4(new_n894), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1174), .A2(new_n913), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n913), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1159), .A2(new_n1160), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT120), .B1(new_n1180), .B2(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n706), .B1(new_n1180), .B2(KEYINPUT57), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1181), .A2(new_n1182), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1172), .A2(new_n756), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n285), .B1(new_n261), .B2(new_n263), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n206), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n788), .A2(new_n217), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n780), .A2(G116), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n786), .A2(G107), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n330), .A2(G41), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n933), .A4(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1194), .B(new_n1198), .C1(new_n420), .C2(new_n777), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n772), .A2(G283), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n783), .A2(G58), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1199), .A2(new_n1035), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT58), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n792), .A2(new_n836), .B1(new_n768), .B2(new_n1120), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n935), .A2(new_n835), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(G132), .C2(new_n930), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1122), .B2(new_n779), .C1(new_n1126), .C2(new_n787), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1208));
  XOR2_X1   g1008(.A(new_n1207), .B(new_n1208), .Z(new_n1209));
  AOI21_X1  g1009(.A(G41), .B1(new_n772), .B2(G124), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n783), .A2(G159), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1210), .A2(new_n258), .A3(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1193), .B(new_n1203), .C1(new_n1209), .C2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(new_n764), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n845), .A2(G50), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1191), .A2(new_n822), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1184), .B2(new_n960), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1190), .A2(new_n1217), .ZN(G375));
  INV_X1    g1018(.A(new_n1139), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1156), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n984), .A3(new_n1150), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n911), .A2(new_n756), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n764), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n937), .A2(new_n317), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT121), .Z(new_n1225));
  NOR2_X1   g1025(.A1(new_n787), .A2(new_n830), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1032), .B1(new_n771), .B2(new_n831), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n935), .A2(new_n536), .B1(new_n208), .B2(new_n788), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n217), .B2(new_n768), .C1(new_n567), .C2(new_n779), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n935), .A2(new_n836), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1201), .B1(new_n1074), .B2(new_n768), .C1(new_n835), .C2(new_n787), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n930), .C2(new_n1119), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n780), .A2(G132), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n791), .A2(G50), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n332), .B1(new_n772), .B2(G128), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1223), .B1(new_n1230), .B2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n845), .A2(G68), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1222), .A2(new_n1238), .A3(new_n822), .A4(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1139), .B2(new_n960), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1221), .A2(new_n1241), .ZN(G381));
  XNOR2_X1  g1042(.A(G375), .B(KEYINPUT122), .ZN(new_n1243));
  INV_X1    g1043(.A(G378), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1044), .A2(new_n1047), .A3(new_n810), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(G381), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G387), .A2(G390), .ZN(new_n1249));
  INV_X1    g1049(.A(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1248), .A2(new_n1251), .ZN(G407));
  INV_X1    g1052(.A(G213), .ZN(new_n1253));
  INV_X1    g1053(.A(G343), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1251), .B2(new_n1248), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n1190), .A2(G378), .A3(new_n1217), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n984), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1217), .B1(new_n1186), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1244), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1253), .A2(G343), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n706), .B1(new_n1220), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n1150), .C1(new_n1265), .C2(new_n1220), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1241), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT123), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(G384), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1250), .A2(KEYINPUT123), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(G384), .A2(new_n1269), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1267), .A2(new_n1271), .A3(new_n1241), .A4(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(G2897), .A3(new_n1262), .A4(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT125), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(G2897), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(G2897), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1262), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1264), .A2(new_n1275), .A3(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1261), .A2(new_n1263), .A3(new_n1276), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT62), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1261), .A2(new_n1286), .A3(new_n1263), .A4(new_n1276), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1282), .A2(new_n1284), .A3(new_n1285), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1246), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(G387), .A2(G390), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1249), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n983), .A2(new_n984), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n959), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1003), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1296), .A2(new_n958), .A3(new_n1086), .A4(new_n1059), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1298), .A3(new_n1290), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1293), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1288), .A2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1261), .A2(new_n1263), .A3(new_n1276), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1302), .B2(KEYINPUT63), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1283), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1285), .A3(new_n1282), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1301), .A2(new_n1306), .ZN(G405));
  AND3_X1   g1107(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1299), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT127), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G375), .A2(new_n1244), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1257), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1257), .B(new_n1311), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1276), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1315), .A2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1313), .A2(new_n1314), .A3(new_n1316), .A4(new_n1276), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


