//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  AND2_X1   g031(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n457));
  NOR2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  OAI21_X1  g033(.A(G137), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(G101), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n463), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n457), .A2(new_n458), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT68), .Z(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(G2105), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n476), .A2(G136), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G138), .B(new_n462), .C1(new_n457), .C2(new_n458), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n462), .B2(G114), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n490), .A2(new_n492), .A3(new_n493), .A4(G2104), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n457), .C2(new_n458), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n488), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n499), .A2(new_n501), .A3(G50), .A4(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n499), .B(new_n501), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G88), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(new_n502), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n503), .A2(new_n504), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n508), .A2(new_n517), .B1(G651), .B2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n514), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI221_X1 g105(.A(new_n527), .B1(new_n505), .B2(new_n528), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n525), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n519), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n498), .B1(new_n535), .B2(KEYINPUT72), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n536), .B1(KEYINPUT72), .B2(new_n535), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n529), .A2(new_n538), .B1(new_n505), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n537), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n498), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT73), .B(G81), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n529), .A2(new_n546), .B1(new_n505), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n545), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n529), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n499), .A2(new_n501), .A3(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(G53), .ZN(new_n566));
  INV_X1    g141(.A(new_n505), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n563), .A2(new_n566), .B1(G91), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n519), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n572), .A2(KEYINPUT76), .A3(G651), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT76), .B1(new_n572), .B2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(G168), .ZN(G286));
  NAND2_X1  g153(.A1(new_n521), .A2(G651), .ZN(new_n579));
  INV_X1    g154(.A(new_n517), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n516), .B1(new_n515), .B2(new_n502), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(G303));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n505), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT77), .A4(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n511), .A2(new_n588), .A3(new_n512), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n514), .A2(G49), .A3(G543), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G288));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n529), .A2(new_n594), .B1(new_n505), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n513), .A2(G61), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT78), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n498), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n498), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n529), .A2(new_n605), .B1(new_n505), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n564), .A2(G54), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n498), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT79), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n567), .A2(G92), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT10), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(new_n618), .B2(G868), .ZN(G284));
  XOR2_X1   g194(.A(G284), .B(KEYINPUT80), .Z(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n576), .ZN(G297));
  XOR2_X1   g197(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n618), .B1(new_n624), .B2(G860), .ZN(G148));
  NOR2_X1   g200(.A1(new_n617), .A2(G559), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n555), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT11), .Z(G282));
  INV_X1    g206(.A(new_n630), .ZN(G323));
  NAND2_X1  g207(.A1(new_n476), .A2(G2104), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  INV_X1    g210(.A(G2100), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n476), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n473), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT82), .B(G2096), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n638), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XOR2_X1   g224(.A(G2427), .B(G2430), .Z(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  OAI221_X1 g247(.A(new_n667), .B1(new_n666), .B2(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n667), .A2(new_n669), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n636), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n682), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(KEYINPUT87), .ZN(new_n692));
  AOI211_X1 g267(.A(new_n687), .B(new_n689), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT88), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n693), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  INV_X1    g273(.A(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(G229));
  XOR2_X1   g276(.A(KEYINPUT31), .B(G11), .Z(new_n702));
  INV_X1    g277(.A(G28), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n703), .B2(KEYINPUT30), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n476), .A2(G141), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n473), .A2(G129), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT26), .Z(new_n712));
  NAND3_X1  g287(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n709), .A2(new_n710), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n708), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT27), .B(G1996), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n706), .B1(new_n707), .B2(new_n643), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G162), .A2(new_n707), .ZN(new_n718));
  AND3_X1   g293(.A1(new_n707), .A2(KEYINPUT95), .A3(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(KEYINPUT95), .B1(new_n707), .B2(G35), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT29), .B(G2090), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  NOR2_X1   g299(.A1(G164), .A2(new_n707), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G27), .B2(new_n707), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n723), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1966), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NOR2_X1   g304(.A1(G168), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n729), .B2(G21), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n717), .B(new_n727), .C1(new_n728), .C2(new_n731), .ZN(new_n732));
  AND2_X1   g307(.A1(KEYINPUT24), .A2(G34), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n707), .B1(KEYINPUT24), .B2(G34), .ZN(new_n734));
  OAI22_X1  g309(.A1(G160), .A2(new_n707), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2084), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n486), .A2(G127), .ZN(new_n737));
  AND2_X1   g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  OAI21_X1  g313(.A(G2105), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT25), .ZN(new_n740));
  NAND2_X1  g315(.A1(G103), .A2(G2104), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G2105), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n476), .A2(G139), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G29), .ZN(new_n747));
  NOR2_X1   g322(.A1(G29), .A2(G33), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2072), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n736), .B(new_n752), .C1(new_n715), .C2(new_n716), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n555), .A2(new_n729), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n729), .B2(G19), .ZN(new_n755));
  INV_X1    g330(.A(G1341), .ZN(new_n756));
  NOR2_X1   g331(.A1(G5), .A2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G171), .B2(G16), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n755), .A2(new_n756), .B1(new_n759), .B2(G1961), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n707), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n476), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n473), .A2(G128), .ZN(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  INV_X1    g343(.A(G2067), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n721), .A2(new_n722), .B1(new_n728), .B2(new_n731), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n770), .B(new_n771), .C1(new_n724), .C2(new_n726), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n732), .A2(new_n753), .A3(new_n760), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n729), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n618), .B2(new_n729), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1348), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n729), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT97), .B(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  INV_X1    g359(.A(new_n775), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n750), .A2(new_n751), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n787), .B1(G1961), .B2(new_n759), .C1(new_n755), .C2(new_n756), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n773), .A2(new_n776), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n590), .A2(new_n591), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n585), .B2(new_n586), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n729), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n729), .B2(G23), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n729), .A2(G6), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n601), .B2(new_n729), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n729), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n729), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT90), .B(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n793), .A2(new_n794), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n800), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n729), .A2(G24), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n608), .B2(new_n729), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(new_n699), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT89), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n476), .A2(G131), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n473), .A2(G119), .ZN(new_n817));
  NOR2_X1   g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n816), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G25), .B(new_n820), .S(G29), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n826));
  NOR4_X1   g401(.A1(new_n814), .A2(new_n815), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n809), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n825), .A2(KEYINPUT91), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n789), .A2(new_n830), .A3(new_n831), .ZN(G150));
  INV_X1    g407(.A(G150), .ZN(G311));
  NOR2_X1   g408(.A1(new_n617), .A2(new_n624), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT102), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n834), .B(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n498), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT100), .B(G55), .Z(new_n840));
  INV_X1    g415(.A(G93), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n529), .A2(new_n840), .B1(new_n505), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n550), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n554), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT101), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT101), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(new_n844), .C1(new_n554), .C2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n837), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT103), .Z(new_n854));
  INV_X1    g429(.A(new_n843), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n714), .B(new_n767), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n494), .A2(KEYINPUT105), .A3(new_n495), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT105), .B1(new_n494), .B2(new_n495), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n488), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n859), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n746), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n866));
  INV_X1    g441(.A(new_n745), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(KEYINPUT106), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n476), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n473), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n634), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n820), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(KEYINPUT107), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n880), .A2(new_n870), .A3(new_n869), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT104), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n643), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n871), .A2(new_n888), .A3(new_n880), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n880), .B1(new_n869), .B2(new_n870), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT108), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(new_n881), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n887), .B(KEYINPUT40), .C1(new_n893), .C2(new_n884), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n884), .B1(new_n892), .B2(new_n881), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n885), .A2(new_n886), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n894), .A2(new_n898), .ZN(G395));
  NAND2_X1  g474(.A1(new_n855), .A2(new_n628), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n849), .B(new_n626), .ZN(new_n901));
  XNOR2_X1  g476(.A(G299), .B(new_n617), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n618), .A2(G299), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n617), .A2(new_n576), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n904), .B1(new_n911), .B2(new_n901), .ZN(new_n912));
  XNOR2_X1  g487(.A(G166), .B(G288), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n608), .B(new_n601), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  XOR2_X1   g490(.A(new_n915), .B(KEYINPUT42), .Z(new_n916));
  XNOR2_X1  g491(.A(new_n912), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n900), .B1(new_n917), .B2(new_n628), .ZN(G295));
  OAI21_X1  g493(.A(new_n900), .B1(new_n917), .B2(new_n628), .ZN(G331));
  XNOR2_X1  g494(.A(G168), .B(KEYINPUT109), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G301), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n846), .A4(new_n848), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(G171), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  XNOR2_X1  g500(.A(G168), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G301), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n846), .A2(new_n924), .A3(new_n927), .A4(new_n848), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n927), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n849), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n923), .A2(new_n929), .A3(new_n903), .A4(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n915), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n910), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n915), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n932), .A2(KEYINPUT111), .A3(new_n935), .A4(new_n933), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n938), .A2(new_n940), .A3(new_n886), .A4(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n931), .A2(new_n903), .A3(new_n928), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n923), .A2(new_n931), .A3(new_n929), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(new_n911), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n915), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n936), .B2(new_n937), .ZN(new_n949));
  AND4_X1   g524(.A1(KEYINPUT43), .A2(new_n948), .A3(new_n949), .A4(new_n941), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n943), .A4(new_n941), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n496), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n485), .A3(new_n487), .A4(new_n860), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n463), .A2(G40), .A3(new_n470), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n714), .B(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n767), .B(new_n769), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n820), .A2(new_n823), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n820), .A2(new_n823), .ZN(new_n971));
  OR3_X1    g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n608), .B(new_n699), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n965), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(KEYINPUT45), .B(new_n961), .C1(new_n488), .C2(new_n496), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n463), .A2(G40), .A3(new_n470), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n728), .B1(new_n962), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT116), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n728), .C1(new_n962), .C2(new_n977), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n982));
  NAND3_X1  g557(.A1(new_n960), .A2(new_n961), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n961), .B1(new_n488), .B2(new_n496), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n964), .B1(new_n984), .B2(KEYINPUT50), .ZN(new_n985));
  INV_X1    g560(.A(G2084), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n988), .A2(G8), .A3(G168), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n960), .A2(new_n961), .A3(new_n976), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT113), .B1(new_n791), .B2(G1976), .ZN(new_n991));
  AND4_X1   g566(.A1(KEYINPUT113), .A2(new_n587), .A3(G1976), .A4(new_n592), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n990), .B(G8), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(G288), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n791), .A2(KEYINPUT113), .A3(G1976), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(G8), .A3(new_n990), .A4(new_n995), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G288), .A2(new_n994), .A3(new_n999), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR3_X1   g581(.A1(G166), .A2(KEYINPUT55), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(G303), .B2(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G2090), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n983), .A2(new_n985), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n960), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n964), .B1(new_n984), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1971), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1010), .B(G8), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G305), .A2(G1981), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n601), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n990), .A4(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1005), .A2(new_n1017), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n982), .B1(new_n960), .B2(new_n961), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n961), .C1(new_n488), .C2(new_n496), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n976), .ZN(new_n1031));
  NOR3_X1   g606(.A1(new_n1028), .A2(G2090), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1027), .B1(new_n1032), .B2(new_n1016), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n982), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n863), .B2(G1384), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1030), .A2(new_n976), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1011), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(KEYINPUT115), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1033), .A2(new_n1041), .A3(G8), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1010), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n989), .A2(new_n1026), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n989), .A2(new_n1026), .A3(new_n1044), .A4(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1046), .A2(new_n1052), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1047), .B1(new_n1054), .B2(new_n1043), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n989), .A2(new_n1026), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1053), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n569), .B2(new_n575), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n568), .B(KEYINPUT57), .C1(new_n574), .C2(new_n573), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1013), .A2(new_n1015), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n983), .A2(new_n985), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n784), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n990), .A2(G2067), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n617), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1074), .B(new_n617), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1348), .B1(new_n983), .B2(new_n985), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1078), .A2(new_n1069), .A3(new_n1076), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n618), .B1(new_n1079), .B2(KEYINPUT120), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(KEYINPUT120), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1059), .A2(new_n1065), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(new_n1066), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT61), .B1(new_n1072), .B2(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n990), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1034), .B2(G1996), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n555), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT59), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n1095), .A3(new_n555), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1096), .B1(KEYINPUT61), .B2(new_n1066), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1089), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1073), .B1(new_n1083), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n1073), .C1(new_n1083), .C2(new_n1098), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n988), .A2(G8), .A3(G286), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n988), .A2(G8), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n988), .A2(KEYINPUT123), .A3(G8), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G286), .A2(G8), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1109), .B(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1105), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1104), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1013), .A2(new_n1015), .A3(new_n724), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n964), .A2(new_n1121), .A3(G2078), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n963), .A2(new_n1123), .A3(new_n1013), .ZN(new_n1124));
  INV_X1    g699(.A(G1961), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1067), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1127), .B2(G171), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1120), .A2(new_n1121), .B1(new_n1067), .B2(new_n1125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n963), .A2(new_n975), .A3(new_n1123), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(G301), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1128), .A2(KEYINPUT124), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1127), .A2(G171), .ZN(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1119), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1026), .A3(new_n1044), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1100), .A2(new_n1102), .A3(new_n1118), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n990), .A2(G8), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1025), .A2(new_n999), .A3(new_n791), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1142), .B2(new_n1020), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1017), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1005), .A2(new_n1025), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1057), .A2(new_n1140), .A3(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1026), .A2(new_n1044), .A3(new_n1136), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1117), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT62), .B(new_n1104), .C1(new_n1113), .C2(new_n1116), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT125), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1153), .A2(new_n1107), .B1(KEYINPUT51), .B2(new_n1115), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT62), .B1(new_n1154), .B2(new_n1104), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1117), .A2(new_n1149), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .A4(new_n1148), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1152), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n974), .B1(new_n1147), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT46), .ZN(new_n1161));
  INV_X1    g736(.A(new_n965), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(G1996), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n965), .A2(KEYINPUT46), .A3(new_n966), .ZN(new_n1164));
  INV_X1    g739(.A(new_n968), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n965), .B1(new_n1165), .B2(new_n714), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT127), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT47), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n972), .A2(new_n965), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G290), .A2(G1986), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n965), .A2(KEYINPUT48), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT48), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1173), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n1162), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n767), .A2(G2067), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n965), .A2(new_n969), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1179), .B1(new_n1180), .B2(new_n970), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1181), .A2(KEYINPUT126), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n965), .B1(new_n1181), .B2(KEYINPUT126), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1178), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1170), .A2(new_n1171), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1160), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g761(.A1(new_n679), .A2(G319), .ZN(new_n1188));
  NOR3_X1   g762(.A1(G229), .A2(new_n1188), .A3(new_n663), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n1189), .B1(new_n896), .B2(new_n897), .ZN(new_n1190));
  AOI21_X1  g764(.A(new_n1190), .B1(new_n952), .B2(new_n953), .ZN(G308));
  OAI211_X1 g765(.A(new_n954), .B(new_n1189), .C1(new_n896), .C2(new_n897), .ZN(G225));
endmodule


