//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NOR2_X1   g0012(.A1(G58), .A2(G68), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n214), .A2(G50), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n207), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT66), .B(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n202), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G107), .A2(G264), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n223), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT5), .B(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G274), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n258), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n255), .B2(new_n253), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n262), .B2(G270), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT82), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G303), .ZN(new_n270));
  INV_X1    g0070(.A(G264), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT68), .B(G1698), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G257), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT76), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(new_n267), .B2(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n265), .A2(KEYINPUT76), .A3(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(new_n268), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n264), .B(new_n270), .C1(new_n275), .C2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n257), .B1(new_n219), .B2(new_n220), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n272), .A2(KEYINPUT68), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(G257), .ZN(new_n287));
  INV_X1    g0087(.A(new_n273), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n277), .A2(new_n268), .A3(new_n278), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n264), .B1(new_n291), .B2(new_n270), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n263), .B1(new_n283), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT83), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(KEYINPUT83), .B(new_n263), .C1(new_n283), .C2(new_n292), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n298));
  INV_X1    g0098(.A(new_n220), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n218), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT84), .A2(KEYINPUT20), .ZN(new_n302));
  AOI21_X1  g0102(.A(G20), .B1(G33), .B2(G283), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n267), .A2(G97), .ZN(new_n304));
  INV_X1    g0104(.A(G116), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n304), .B1(G20), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n302), .B1(new_n301), .B2(new_n306), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n305), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n299), .A2(new_n310), .A3(new_n218), .A4(new_n300), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n267), .A2(G1), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n311), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n297), .B1(new_n309), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n295), .A2(KEYINPUT21), .A3(new_n296), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT85), .ZN(new_n318));
  OAI211_X1 g0118(.A(G179), .B(new_n263), .C1(new_n283), .C2(new_n292), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n309), .A2(new_n315), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n317), .B2(new_n321), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n295), .A2(new_n296), .A3(new_n316), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT86), .B(KEYINPUT21), .Z(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n322), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT72), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G20), .A2(G33), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G150), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n267), .A2(G20), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n329), .B(new_n331), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n310), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n301), .B1(new_n246), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n312), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n206), .A2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G50), .A3(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n337), .A2(KEYINPUT9), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT9), .B1(new_n337), .B2(new_n340), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n258), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  XOR2_X1   g0146(.A(KEYINPUT67), .B(G226), .Z(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G41), .ZN(new_n349));
  AOI21_X1  g0149(.A(G1), .B1(new_n349), .B2(new_n254), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(new_n258), .A3(G274), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT3), .B(G33), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(new_n274), .A3(G222), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(G223), .A3(G1698), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n269), .A2(G77), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT69), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT69), .A4(new_n357), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n282), .ZN(new_n363));
  OAI211_X1 g0163(.A(G190), .B(new_n353), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n343), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  INV_X1    g0166(.A(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n352), .B1(new_n367), .B2(new_n360), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n328), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n353), .B1(new_n361), .B2(new_n363), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT10), .B1(new_n372), .B2(G200), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT72), .A3(new_n343), .A4(new_n364), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n342), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n337), .A2(KEYINPUT9), .A3(new_n340), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n364), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n372), .A2(G200), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n343), .B2(new_n364), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT10), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n351), .B1(new_n235), .B2(new_n345), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n274), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n386));
  INV_X1    g0186(.A(G87), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n386), .A2(new_n279), .B1(new_n267), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n388), .B2(new_n282), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G179), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n297), .B2(new_n389), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n207), .B1(new_n203), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR3_X1   g0195(.A1(new_n395), .A2(G20), .A3(G33), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n393), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n398), .B2(new_n213), .ZN(new_n399));
  INV_X1    g0199(.A(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n279), .A2(new_n403), .A3(new_n207), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n279), .B2(new_n207), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n402), .B(KEYINPUT16), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n403), .B1(new_n354), .B2(G20), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n202), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n399), .A2(new_n400), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n301), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n334), .B1(new_n206), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n338), .A2(new_n415), .B1(new_n336), .B2(new_n334), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n391), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n391), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G226), .A2(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n284), .A2(new_n286), .ZN(new_n423));
  INV_X1    g0223(.A(G223), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n290), .B1(G33), .B2(G87), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n281), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n427), .B2(new_n385), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n389), .A2(G190), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n414), .A2(new_n428), .A3(new_n416), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n389), .A2(new_n369), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n434), .B(new_n385), .C1(new_n388), .C2(new_n282), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .A3(new_n416), .A4(new_n414), .ZN(new_n437));
  AND4_X1   g0237(.A1(new_n419), .A2(new_n421), .A3(new_n432), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n372), .A2(new_n297), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n337), .A2(new_n340), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(G179), .C2(new_n372), .ZN(new_n441));
  INV_X1    g0241(.A(G244), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n351), .B1(new_n442), .B2(new_n345), .ZN(new_n443));
  OAI221_X1 g0243(.A(new_n354), .B1(new_n224), .B2(new_n272), .C1(new_n235), .C2(new_n423), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n354), .A2(G107), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n281), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G179), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n447), .A2(G169), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n339), .A2(G77), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n312), .A2(new_n451), .B1(G77), .B2(new_n310), .ZN(new_n452));
  XOR2_X1   g0252(.A(KEYINPUT15), .B(G87), .Z(new_n453));
  INV_X1    g0253(.A(KEYINPUT70), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT15), .B(G87), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n457), .A3(new_n332), .ZN(new_n458));
  INV_X1    g0258(.A(new_n334), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n459), .A2(new_n330), .B1(G20), .B2(G77), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n452), .B1(new_n461), .B2(new_n301), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n449), .A2(new_n450), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n447), .A2(G190), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n301), .ZN(new_n466));
  INV_X1    g0266(.A(new_n452), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n466), .B(new_n467), .C1(new_n369), .C2(new_n447), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n468), .B2(KEYINPUT71), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT71), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n462), .B(new_n470), .C1(new_n369), .C2(new_n447), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n463), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n384), .A2(new_n438), .A3(new_n441), .A4(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n330), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n474));
  INV_X1    g0274(.A(G77), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n333), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT11), .B1(new_n476), .B2(new_n301), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n310), .A2(G68), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT12), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(KEYINPUT11), .A3(new_n301), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n338), .A2(G68), .A3(new_n339), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G238), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n351), .B1(new_n485), .B2(new_n345), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT74), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n235), .A2(new_n272), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n274), .B2(G226), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n491), .B2(new_n269), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n492), .B2(new_n282), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n284), .A2(new_n286), .A3(G226), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n269), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n489), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n488), .B(new_n282), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n487), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT13), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n282), .B1(new_n496), .B2(new_n497), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n498), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT13), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n487), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n297), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT14), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n504), .B2(new_n487), .ZN(new_n509));
  AOI211_X1 g0309(.A(KEYINPUT13), .B(new_n486), .C1(new_n503), .C2(new_n498), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n507), .A2(new_n508), .B1(new_n511), .B2(G179), .ZN(new_n512));
  OAI21_X1  g0312(.A(G169), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT14), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n484), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(G190), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n501), .A2(new_n506), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n516), .A2(new_n518), .A3(new_n484), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT75), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n501), .A2(G179), .A3(new_n506), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n513), .B2(KEYINPUT14), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n508), .B1(new_n517), .B2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n483), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n516), .A2(new_n518), .A3(new_n484), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n473), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n295), .A2(G200), .A3(new_n296), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n320), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n434), .B1(new_n295), .B2(new_n296), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT87), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n295), .A2(new_n296), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G190), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT87), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n320), .A4(new_n529), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n284), .A2(new_n286), .A3(G244), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT4), .B1(new_n290), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n266), .A2(new_n268), .A3(G250), .A4(G1698), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n266), .A2(new_n268), .A3(new_n284), .A4(new_n286), .ZN(new_n543));
  NAND2_X1  g0343(.A1(KEYINPUT4), .A2(G244), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n541), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n282), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n260), .B1(new_n262), .B2(G257), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n369), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT79), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n548), .A2(new_n549), .B1(new_n550), .B2(new_n434), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n310), .A2(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n314), .B2(G97), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n409), .A2(new_n410), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT78), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n354), .A2(new_n403), .A3(G20), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT7), .B1(new_n269), .B2(new_n207), .ZN(new_n560));
  OAI211_X1 g0360(.A(KEYINPUT78), .B(G107), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  INV_X1    g0362(.A(G97), .ZN(new_n563));
  INV_X1    g0363(.A(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n564), .A2(KEYINPUT6), .A3(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n330), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n558), .A2(new_n561), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n554), .B1(new_n571), .B2(new_n301), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n256), .A2(new_n258), .ZN(new_n573));
  INV_X1    g0373(.A(G257), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n573), .A2(new_n574), .B1(new_n256), .B2(new_n259), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n279), .B2(new_n538), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n354), .A2(new_n274), .A3(KEYINPUT4), .A4(G244), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n541), .A3(new_n542), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n575), .B1(new_n579), .B2(new_n282), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(KEYINPUT79), .A3(G190), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n551), .A2(new_n572), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(G169), .B1(new_n546), .B2(new_n547), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT80), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(new_n550), .B2(G179), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n580), .A2(KEYINPUT80), .A3(new_n448), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n561), .A2(new_n570), .ZN(new_n587));
  AOI21_X1  g0387(.A(KEYINPUT78), .B1(new_n555), .B2(G107), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n301), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n553), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n267), .A2(new_n305), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G244), .A2(G1698), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n423), .B2(new_n485), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n290), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n258), .A2(G274), .A3(new_n255), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n206), .A2(G45), .ZN(new_n597));
  AND2_X1   g0397(.A1(G33), .A2(G41), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G1), .A2(G13), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(G250), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT81), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n595), .A2(new_n281), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(G200), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n207), .B1(new_n489), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n566), .A2(new_n387), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n606), .A2(new_n607), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n277), .A2(new_n278), .A3(new_n207), .A4(new_n268), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n609), .B1(new_n202), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n301), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n455), .A2(new_n457), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n336), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n314), .A2(G87), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n274), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n279), .B1(new_n267), .B2(new_n305), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n282), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n596), .A2(new_n600), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n596), .A2(KEYINPUT81), .A3(new_n600), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(G190), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n604), .A2(new_n616), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n603), .A2(new_n297), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n619), .A2(new_n448), .A3(new_n624), .ZN(new_n628));
  INV_X1    g0428(.A(new_n314), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n612), .B(new_n614), .C1(new_n629), .C2(new_n613), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n582), .A2(new_n591), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n284), .A2(new_n286), .A3(G250), .ZN(new_n635));
  NAND2_X1  g0435(.A1(G257), .A2(G1698), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n290), .ZN(new_n638));
  NAND2_X1  g0438(.A1(G33), .A2(G294), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n281), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n573), .A2(new_n271), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n634), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n260), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n262), .A2(G264), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n637), .A2(new_n290), .B1(G33), .B2(G294), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT90), .B(new_n644), .C1(new_n645), .C2(new_n281), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n642), .A2(G179), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n281), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G169), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G1), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(G20), .A3(new_n564), .ZN(new_n653));
  AND2_X1   g0453(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(KEYINPUT89), .A2(KEYINPUT25), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AOI211_X1 g0457(.A(new_n655), .B(new_n657), .C1(G107), .C2(new_n314), .ZN(new_n658));
  NAND2_X1  g0458(.A1(KEYINPUT22), .A2(G87), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n610), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT22), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n207), .A2(G87), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n269), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT23), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n207), .B2(G107), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n564), .A2(KEYINPUT23), .A3(G20), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n592), .B2(new_n207), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n661), .A2(KEYINPUT88), .A3(new_n664), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT88), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n660), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n669), .A2(new_n672), .A3(KEYINPUT24), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n301), .B1(new_n672), .B2(KEYINPUT24), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n658), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n650), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n648), .A2(G190), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n369), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n633), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  AND4_X1   g0482(.A1(new_n327), .A2(new_n528), .A3(new_n537), .A4(new_n682), .ZN(G372));
  NAND2_X1  g0483(.A1(new_n437), .A2(new_n432), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n526), .A2(new_n463), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n524), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n419), .A2(new_n421), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n384), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n441), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n528), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n324), .A2(new_n325), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n676), .A3(new_n321), .A4(new_n317), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT91), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n633), .A2(new_n681), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n317), .A2(new_n321), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(KEYINPUT91), .A3(new_n693), .A4(new_n676), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n631), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT26), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n626), .A2(new_n631), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n591), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n702), .B1(new_n591), .B2(new_n703), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n691), .B1(new_n692), .B2(new_n709), .ZN(G369));
  NAND2_X1  g0510(.A1(new_n652), .A2(new_n207), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT92), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G343), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n537), .B(new_n327), .C1(new_n320), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n320), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n317), .A2(new_n321), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n326), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n676), .A2(new_n718), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n675), .A2(new_n718), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n680), .B2(new_n675), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(new_n676), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(G330), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n327), .A2(new_n718), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n725), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n210), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n607), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n737), .A2(KEYINPUT93), .B1(new_n216), .B2(new_n735), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(KEYINPUT93), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  INV_X1    g0540(.A(KEYINPUT29), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n708), .A2(new_n741), .A3(new_n719), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT26), .B1(new_n743), .B2(new_n632), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n631), .B1(new_n744), .B2(new_n704), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n722), .A2(KEYINPUT85), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n324), .A2(new_n325), .B1(new_n650), .B2(new_n675), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n697), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT95), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n749), .A2(new_n697), .A3(KEYINPUT95), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n718), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n742), .B1(new_n754), .B2(new_n741), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n537), .A2(new_n327), .A3(new_n682), .A4(new_n719), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT30), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n618), .A2(new_n282), .B1(new_n622), .B2(new_n623), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n642), .A2(new_n580), .A3(new_n646), .A4(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n759), .B2(new_n319), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n642), .A2(new_n646), .ZN(new_n761));
  INV_X1    g0561(.A(new_n319), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n550), .A2(new_n603), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT30), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n679), .A2(new_n448), .A3(new_n550), .A4(new_n603), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n760), .B(new_n764), .C1(new_n533), .C2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT31), .B1(new_n766), .B2(new_n718), .ZN(new_n768));
  OAI21_X1  g0568(.A(KEYINPUT94), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n766), .A2(new_n718), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT31), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT94), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n756), .A2(new_n769), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n755), .B1(G330), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n740), .B1(new_n777), .B2(G1), .ZN(G364));
  NOR2_X1   g0578(.A1(new_n651), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n206), .B1(new_n779), .B2(G45), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n734), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT97), .B1(new_n724), .B2(G330), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT97), .ZN(new_n785));
  INV_X1    g0585(.A(G330), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n785), .B(new_n786), .C1(new_n720), .C2(new_n723), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT96), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n724), .B2(G330), .ZN(new_n790));
  INV_X1    g0590(.A(new_n724), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(KEYINPUT96), .A3(new_n786), .ZN(new_n792));
  AND4_X1   g0592(.A1(new_n783), .A2(new_n788), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT98), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n221), .B1(G20), .B2(new_n297), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT100), .Z(new_n800));
  NOR2_X1   g0600(.A1(new_n733), .A2(new_n269), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G355), .B1(new_n305), .B2(new_n733), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n733), .A2(new_n290), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G45), .B2(new_n216), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n251), .A2(new_n254), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n800), .B1(new_n806), .B2(KEYINPUT99), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(KEYINPUT99), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n207), .A2(new_n448), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n810), .A2(new_n369), .A3(G190), .ZN(new_n811));
  INV_X1    g0611(.A(G317), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n812), .A2(KEYINPUT33), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n809), .A2(G190), .A3(G200), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT101), .B(G326), .Z(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n434), .A2(G179), .A3(G200), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n207), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n818), .C2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n810), .A2(new_n434), .A3(G200), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n207), .A2(G179), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(new_n434), .A3(new_n369), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(G322), .B1(G329), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G311), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n810), .A2(G190), .A3(G200), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n826), .B(new_n269), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n823), .A2(new_n434), .A3(G200), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n823), .A2(G190), .A3(G200), .ZN(new_n833));
  INV_X1    g0633(.A(G303), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n831), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n821), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n822), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n354), .B1(new_n829), .B2(new_n475), .C1(new_n201), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT32), .B1(new_n824), .B2(new_n395), .ZN(new_n839));
  INV_X1    g0639(.A(new_n811), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n839), .B1(new_n246), .B2(new_n816), .C1(new_n840), .C2(new_n202), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n824), .A2(KEYINPUT32), .A3(new_n395), .ZN(new_n842));
  INV_X1    g0642(.A(new_n820), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G97), .ZN(new_n844));
  INV_X1    g0644(.A(new_n833), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(G87), .ZN(new_n846));
  INV_X1    g0646(.A(new_n832), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(G107), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n842), .A2(new_n844), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n838), .A2(new_n841), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n795), .B1(new_n836), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n808), .A2(new_n851), .A3(new_n782), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n791), .B2(new_n798), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n794), .A2(new_n853), .ZN(G396));
  NAND2_X1  g0654(.A1(new_n466), .A2(new_n467), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n718), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT103), .B1(new_n472), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n447), .A2(new_n369), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT71), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(new_n471), .A3(new_n464), .ZN(new_n860));
  INV_X1    g0660(.A(new_n463), .ZN(new_n861));
  AND4_X1   g0661(.A1(KEYINPUT103), .A2(new_n860), .A3(new_n861), .A4(new_n856), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n719), .ZN(new_n863));
  NOR3_X1   g0663(.A1(new_n857), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n709), .B2(new_n718), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n857), .A2(new_n862), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n708), .A2(new_n719), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n776), .A2(G330), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n782), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n795), .A2(new_n796), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n782), .B1(new_n874), .B2(G77), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n816), .A2(new_n834), .B1(new_n833), .B2(new_n564), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(G87), .B2(new_n847), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n354), .B1(new_n822), .B2(G294), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n828), .A2(G116), .B1(G311), .B2(new_n825), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G283), .A2(new_n811), .B1(new_n843), .B2(G97), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(G143), .A2(new_n822), .B1(new_n828), .B2(G159), .ZN(new_n882));
  INV_X1    g0682(.A(G137), .ZN(new_n883));
  INV_X1    g0683(.A(G150), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n882), .B1(new_n883), .B2(new_n816), .C1(new_n884), .C2(new_n840), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT34), .Z(new_n886));
  NAND2_X1  g0686(.A1(new_n847), .A2(G68), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n246), .B2(new_n833), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n843), .A2(G58), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n279), .B1(new_n825), .B2(G132), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n881), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n875), .B1(new_n895), .B2(new_n795), .ZN(new_n896));
  INV_X1    g0696(.A(new_n864), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n797), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n872), .A2(new_n898), .ZN(G384));
  NAND4_X1  g0699(.A1(new_n419), .A2(new_n421), .A3(new_n432), .A4(new_n437), .ZN(new_n900));
  INV_X1    g0700(.A(new_n716), .ZN(new_n901));
  INV_X1    g0701(.A(new_n301), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(new_n903), .B2(new_n408), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n407), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g0706(.A(KEYINPUT106), .B(new_n902), .C1(new_n903), .C2(new_n408), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n416), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n901), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(new_n430), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n908), .B2(new_n391), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n901), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n417), .A2(new_n901), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n418), .A2(new_n915), .A3(new_n910), .A4(new_n430), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT38), .B(new_n909), .C1(new_n914), .C2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n900), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n418), .A2(new_n915), .A3(new_n430), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT37), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n916), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT105), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n524), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n719), .A2(new_n484), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n519), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT105), .B(new_n483), .C1(new_n522), .C2(new_n523), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n526), .A2(new_n514), .A3(new_n512), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n930), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n767), .A2(new_n768), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n756), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n927), .A2(new_n936), .A3(new_n938), .A4(new_n897), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT40), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n909), .B1(new_n914), .B2(new_n917), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n925), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n918), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n864), .B1(new_n933), .B2(new_n935), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n938), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n528), .A2(new_n938), .ZN(new_n948));
  OAI21_X1  g0748(.A(G330), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT107), .Z(new_n951));
  NOR2_X1   g0751(.A1(new_n861), .A2(new_n718), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n868), .A2(new_n953), .B1(new_n935), .B2(new_n933), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT39), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n927), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n942), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n718), .B1(new_n929), .B2(new_n932), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n688), .A2(new_n716), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n690), .B1(new_n755), .B2(new_n528), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n951), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n951), .A2(new_n964), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n206), .B2(new_n779), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n967), .B2(KEYINPUT108), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(KEYINPUT108), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n393), .A2(G77), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n247), .B1(new_n216), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(G1), .A3(new_n651), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n973), .A2(G116), .A3(new_n222), .A4(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT104), .B(KEYINPUT36), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n969), .A2(new_n972), .A3(new_n977), .ZN(G367));
  OR2_X1    g0778(.A1(new_n719), .A2(new_n616), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(new_n631), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n632), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT43), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n582), .A2(new_n591), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n590), .A2(new_n718), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT109), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n591), .B1(new_n992), .B2(new_n676), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n743), .A2(new_n718), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n728), .A3(new_n730), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n993), .A2(new_n719), .B1(new_n996), .B2(KEYINPUT42), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n985), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n985), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n989), .A2(new_n994), .A3(new_n991), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n729), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1004), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n734), .B(KEYINPUT41), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n724), .A2(G330), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n730), .A2(new_n728), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n746), .A2(new_n747), .A3(new_n693), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n728), .A2(new_n1011), .A3(new_n719), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(new_n788), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n725), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1022), .B2(new_n1005), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1026));
  NAND3_X1  g0826(.A1(new_n1022), .A2(new_n1005), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n731), .B2(new_n995), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1025), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n729), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1025), .A2(new_n729), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1019), .A2(new_n1032), .A3(new_n777), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1008), .B1(new_n1034), .B2(new_n777), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n780), .B1(new_n1035), .B2(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1037), .B(new_n1008), .C1(new_n1034), .C2(new_n777), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1007), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n803), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1040), .A2(new_n241), .B1(new_n210), .B2(new_n613), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n837), .A2(new_n884), .B1(new_n829), .B2(new_n246), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n269), .B(new_n1042), .C1(G137), .C2(new_n825), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n816), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(G143), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n843), .A2(G68), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n832), .A2(new_n475), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n811), .B2(G159), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n201), .B2(new_n833), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n833), .A2(new_n305), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT46), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n820), .A2(new_n564), .B1(new_n832), .B2(new_n563), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G294), .B2(new_n811), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n822), .A2(G303), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT113), .B(G317), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n828), .A2(G283), .B1(new_n825), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n290), .B1(new_n1044), .B2(G311), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1047), .A2(new_n1050), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT47), .Z(new_n1061));
  INV_X1    g0861(.A(new_n795), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n782), .B1(new_n800), .B2(new_n1041), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT114), .Z(new_n1064));
  INV_X1    g0864(.A(new_n798), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n982), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1039), .A2(new_n1066), .ZN(G387));
  NAND2_X1  g0867(.A1(new_n1019), .A2(new_n781), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n728), .A2(new_n1065), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1056), .A2(new_n822), .B1(new_n828), .B2(G303), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1044), .A2(G322), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n827), .C2(new_n840), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n843), .A2(G283), .B1(new_n845), .B2(G294), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n279), .B1(new_n832), .B2(new_n305), .C1(new_n817), .C2(new_n824), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n837), .A2(new_n246), .B1(new_n824), .B2(new_n884), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G68), .B2(new_n828), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n816), .A2(new_n395), .B1(new_n833), .B2(new_n475), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n459), .B2(new_n811), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n613), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n843), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n279), .B1(new_n847), .B2(G97), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1084), .A2(new_n1086), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1062), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n736), .ZN(new_n1092));
  AOI211_X1 g0892(.A(G45), .B(new_n1092), .C1(G68), .C2(G77), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n334), .A2(G50), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT50), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1040), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n238), .B2(new_n254), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n801), .A2(new_n1092), .B1(new_n564), .B2(new_n733), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(KEYINPUT115), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT115), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1100), .A2(new_n800), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n783), .B(new_n1091), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT116), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1019), .A2(new_n777), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n734), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1019), .A2(new_n777), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1068), .B1(new_n1069), .B2(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(G393));
  OAI22_X1  g0907(.A1(new_n1040), .A2(new_n245), .B1(new_n563), .B2(new_n210), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n782), .B1(new_n800), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n822), .A2(G159), .B1(new_n1044), .B2(G150), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT51), .Z(new_n1111));
  AOI21_X1  g0911(.A(new_n279), .B1(new_n825), .B2(G143), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n845), .A2(G68), .B1(new_n847), .B2(G87), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n820), .A2(new_n475), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n459), .B2(new_n828), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n246), .B2(new_n840), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n822), .A2(G311), .B1(new_n1044), .B2(G317), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT52), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n354), .B1(new_n825), .B2(G322), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n829), .B2(new_n818), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n848), .B1(new_n840), .B2(new_n834), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n820), .A2(new_n305), .B1(new_n833), .B2(new_n831), .ZN(new_n1124));
  OR3_X1    g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1114), .A2(new_n1118), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1109), .B1(new_n1126), .B2(new_n795), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n995), .B2(new_n1065), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n780), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1034), .A2(new_n734), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1104), .A2(new_n1129), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(G390));
  NOR2_X1   g0934(.A1(new_n864), .A2(new_n786), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n936), .A2(new_n938), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n959), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n927), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n750), .A2(new_n751), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1140), .A2(new_n707), .A3(new_n753), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1141), .A2(new_n719), .A3(new_n867), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n953), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1139), .B1(new_n1143), .B2(new_n936), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n718), .B(new_n866), .C1(new_n700), .C2(new_n707), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n936), .B1(new_n1145), .B2(new_n952), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n1138), .B1(new_n957), .B2(new_n958), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1137), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1139), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n952), .B1(new_n754), .B2(new_n867), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n936), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n957), .A2(new_n958), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n954), .B2(new_n959), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n776), .A2(new_n936), .A3(G330), .A4(new_n897), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1148), .A2(new_n781), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n782), .B1(new_n874), .B2(new_n459), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n837), .A2(new_n305), .B1(new_n824), .B2(new_n818), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n354), .B(new_n1159), .C1(G97), .C2(new_n828), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n816), .A2(new_n831), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1161), .B(new_n1115), .C1(G107), .C2(new_n811), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1160), .A2(new_n1162), .A3(new_n846), .A4(new_n887), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n354), .B1(new_n832), .B2(new_n246), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT121), .ZN(new_n1165));
  INV_X1    g0965(.A(G132), .ZN(new_n1166));
  INV_X1    g0966(.A(G125), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n837), .A2(new_n1166), .B1(new_n824), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n828), .B2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n840), .A2(new_n883), .B1(new_n395), .B2(new_n820), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G128), .B2(new_n1044), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n833), .A2(new_n884), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT53), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1163), .B1(new_n1165), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1158), .B1(new_n1177), .B2(new_n795), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1153), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n797), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1157), .A2(KEYINPUT122), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT122), .B1(new_n1157), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1152), .A2(new_n1155), .A3(new_n1154), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1136), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n528), .A2(new_n938), .A3(G330), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT118), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT118), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n528), .A2(new_n938), .A3(new_n1189), .A4(G330), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n741), .B1(new_n1141), .B2(new_n719), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n742), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n528), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n691), .A3(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1145), .A2(new_n952), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n776), .A2(G330), .A3(new_n897), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1151), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1198), .B2(new_n1136), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n938), .A2(new_n1135), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1151), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1150), .A2(new_n1202), .A3(new_n1155), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1195), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT120), .B1(new_n1186), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1150), .A2(new_n1202), .A3(new_n1155), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n963), .B(new_n1191), .C1(new_n1208), .C2(new_n1199), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n734), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT119), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1204), .A2(KEYINPUT119), .A3(new_n1156), .A4(new_n1148), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1183), .B1(new_n1211), .B2(new_n1215), .ZN(G378));
  NAND2_X1  g1016(.A1(new_n384), .A2(new_n441), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1217), .A2(new_n440), .A3(new_n901), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n901), .A2(new_n440), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n384), .A2(new_n441), .A3(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n947), .B2(G330), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n786), .B(new_n1224), .C1(new_n940), .C2(new_n946), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n962), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n962), .ZN(new_n1229));
  AND4_X1   g1029(.A1(new_n945), .A2(new_n936), .A3(new_n897), .A4(new_n938), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1230), .A2(new_n943), .B1(new_n939), .B2(KEYINPUT40), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1224), .B1(new_n1231), .B2(new_n786), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n947), .A2(G330), .A3(new_n1225), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n781), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1224), .A2(new_n796), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n782), .B1(new_n874), .B2(G50), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n840), .A2(new_n1166), .B1(new_n816), .B2(new_n1167), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(G128), .A2(new_n822), .B1(new_n828), .B2(G137), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n833), .B2(new_n1169), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G150), .C2(new_n843), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n847), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n279), .A2(new_n349), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1046), .B1(new_n831), .B2(new_n824), .C1(new_n837), .C2(new_n564), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n1087), .C2(new_n828), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n832), .A2(new_n201), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G77), .B2(new_n845), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n811), .A2(G97), .B1(new_n1044), .B2(G116), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT58), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1248), .B(new_n246), .C1(G33), .C2(G41), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1247), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1237), .B1(new_n1259), .B2(new_n795), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1236), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1235), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1195), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT119), .B1(new_n1186), .B2(new_n1204), .ZN(new_n1264));
  NOR3_X1   g1064(.A1(new_n1206), .A2(new_n1209), .A3(new_n1212), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n962), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1232), .A2(new_n1229), .A3(new_n1233), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT57), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n735), .B1(new_n1266), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT57), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1195), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1262), .B1(new_n1272), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(G375));
  NAND2_X1  g1078(.A1(new_n1200), .A2(new_n1203), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n781), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1151), .A2(new_n796), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT123), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n783), .B1(new_n873), .B2(new_n202), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n828), .A2(G150), .B1(G128), .B2(new_n825), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n883), .B2(new_n837), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1285), .A2(new_n279), .A3(new_n1251), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(G132), .A2(new_n1044), .B1(new_n845), .B2(G159), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n843), .A2(G50), .B1(new_n811), .B2(new_n1170), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n816), .A2(new_n818), .B1(new_n833), .B2(new_n563), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1048), .B(new_n1290), .C1(G116), .C2(new_n811), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n354), .B1(new_n828), .B2(G107), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n822), .A2(G283), .B1(G303), .B2(new_n825), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1291), .A2(new_n1088), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n1282), .B(new_n1283), .C1(new_n1062), .C2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1280), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1279), .A2(new_n1263), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1008), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1209), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1298), .B1(new_n1299), .B2(new_n1301), .ZN(G381));
  OR2_X1    g1102(.A1(G396), .A2(G393), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1133), .A2(new_n872), .A3(new_n898), .ZN(new_n1304));
  NOR4_X1   g1104(.A1(G387), .A2(new_n1303), .A3(G381), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1306), .A2(new_n734), .A3(new_n1205), .A4(new_n1210), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1157), .A2(new_n1180), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1305), .A2(new_n1307), .A3(new_n1308), .A4(new_n1277), .ZN(G407));
  OAI21_X1  g1109(.A(new_n1308), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n717), .A2(G213), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G407), .B(G213), .C1(G375), .C2(new_n1312), .ZN(G409));
  AOI22_X1  g1113(.A1(new_n1269), .A2(new_n781), .B1(new_n1236), .B2(new_n1260), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT57), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n734), .B1(new_n1274), .B2(new_n1270), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G378), .B(new_n1314), .C1(new_n1315), .C2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1269), .A2(new_n1300), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1262), .B1(new_n1266), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT124), .B1(new_n1320), .B2(new_n1310), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1314), .B1(new_n1274), .B2(new_n1318), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT124), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1322), .A2(new_n1307), .A3(new_n1323), .A4(new_n1308), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1317), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1209), .A2(KEYINPUT60), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1326), .A2(new_n1299), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n735), .B1(new_n1326), .B2(new_n1299), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1298), .ZN(new_n1330));
  OR2_X1    g1130(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1329), .A2(new_n1298), .A3(new_n1331), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1325), .A2(new_n1311), .A3(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT62), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1325), .A2(new_n1311), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n717), .A2(G213), .A3(G2897), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1297), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1333), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1335), .B(new_n1340), .C1(new_n1341), .C2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1340), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1339), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1325), .A2(new_n1349), .A3(new_n1311), .A4(new_n1336), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1338), .A2(new_n1347), .A3(new_n1348), .A4(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G387), .A2(new_n1133), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT126), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(G396), .B(G393), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1039), .A2(new_n1066), .A3(G390), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(KEYINPUT126), .ZN(new_n1358));
  AOI22_X1  g1158(.A1(new_n1358), .A2(new_n1354), .B1(new_n1352), .B2(new_n1355), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1357), .A2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1351), .A2(new_n1360), .ZN(new_n1361));
  AOI21_X1  g1161(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1346), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1337), .A2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1358), .A2(new_n1354), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1352), .A2(new_n1355), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1356), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1325), .A2(KEYINPUT63), .A3(new_n1311), .A4(new_n1336), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1362), .A2(new_n1364), .A3(new_n1368), .A4(new_n1369), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1361), .A2(new_n1370), .ZN(G405));
  INV_X1    g1171(.A(KEYINPUT127), .ZN(new_n1372));
  OAI211_X1 g1172(.A(new_n1317), .B(new_n1372), .C1(new_n1277), .C2(new_n1310), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1360), .A2(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1373), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1368), .A2(new_n1375), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1374), .A2(new_n1376), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1317), .B1(new_n1277), .B2(new_n1310), .ZN(new_n1378));
  AND2_X1   g1178(.A1(new_n1378), .A2(KEYINPUT127), .ZN(new_n1379));
  OR2_X1    g1179(.A1(new_n1379), .A2(new_n1336), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1377), .A2(new_n1380), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1379), .A2(new_n1336), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1382), .A2(new_n1374), .A3(new_n1376), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1381), .A2(new_n1383), .ZN(G402));
endmodule


