//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  OR2_X1    g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n206), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT68), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n208), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT0), .B(G128), .Z(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n215), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT81), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  AOI21_X1  g045(.A(G101), .B1(new_n221), .B2(G107), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G101), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT82), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n221), .B2(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(KEYINPUT82), .A3(G104), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT81), .B(G107), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(new_n241), .C1(new_n242), .C2(G104), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(G104), .B2(new_n223), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n242), .B2(new_n222), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n243), .A2(G101), .B1(new_n246), .B2(new_n232), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n248), .A2(new_n206), .A3(new_n208), .A4(G128), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n238), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(KEYINPUT83), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n260), .B(KEYINPUT1), .C1(new_n207), .C2(G146), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(G128), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n249), .B1(new_n262), .B2(new_n216), .ZN(new_n263));
  AOI21_X1  g077(.A(G104), .B1(new_n224), .B2(new_n226), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n240), .A2(new_n241), .ZN(new_n265));
  OAI21_X1  g079(.A(G101), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n233), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT84), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(G128), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n260), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n216), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n250), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n233), .A4(new_n266), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT10), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n258), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(KEYINPUT85), .B(KEYINPUT10), .C1(new_n268), .C2(new_n274), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n204), .B(new_n257), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT86), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n263), .A2(new_n267), .A3(KEYINPUT84), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n273), .B1(new_n247), .B2(new_n272), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n275), .A2(new_n258), .A3(new_n276), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n287), .A2(KEYINPUT86), .A3(new_n204), .A4(new_n257), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n249), .B1(new_n216), .B2(new_n252), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n267), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n275), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT12), .B1(new_n292), .B2(new_n203), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n204), .C1(new_n275), .C2(new_n291), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G227), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT80), .ZN(new_n301));
  XNOR2_X1  g115(.A(G110), .B(G140), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n281), .B2(new_n288), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n287), .A2(new_n257), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n203), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n298), .A2(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n192), .B1(new_n307), .B2(G469), .ZN(new_n308));
  INV_X1    g122(.A(new_n303), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n289), .B2(new_n306), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n303), .B(new_n296), .C1(new_n281), .C2(new_n288), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n190), .B(new_n191), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n189), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT66), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n317), .A3(G116), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n318), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n323), .A3(G119), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n318), .A2(new_n324), .A3(KEYINPUT5), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT89), .B1(new_n318), .B2(KEYINPUT5), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n319), .A2(G113), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n318), .A3(new_n324), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n330), .A3(new_n247), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n324), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n328), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(new_n330), .B1(new_n230), .B2(new_n236), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n334), .A2(new_n234), .A3(KEYINPUT88), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT88), .B1(new_n334), .B2(new_n234), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G122), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n331), .C1(new_n335), .C2(new_n336), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n340), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(KEYINPUT6), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT88), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n345));
  INV_X1    g159(.A(new_n330), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n329), .B1(new_n318), .B2(new_n324), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n237), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n344), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(new_n234), .A3(KEYINPUT88), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n338), .B1(new_n351), .B2(new_n331), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n337), .A2(new_n354), .A3(new_n339), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n342), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n211), .A2(new_n212), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(G125), .B2(new_n254), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n299), .A2(G224), .ZN(new_n362));
  XOR2_X1   g176(.A(new_n362), .B(KEYINPUT91), .Z(new_n363));
  XOR2_X1   g177(.A(new_n361), .B(new_n363), .Z(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n360), .A2(KEYINPUT93), .B1(KEYINPUT7), .B2(new_n362), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(new_n361), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n361), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n341), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n338), .B(KEYINPUT8), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n319), .A2(G113), .A3(new_n326), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n372), .A2(KEYINPUT92), .ZN(new_n373));
  INV_X1    g187(.A(new_n325), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n374), .B1(new_n372), .B2(KEYINPUT92), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n346), .B(new_n267), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n247), .B1(new_n327), .B2(new_n330), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n191), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G210), .B1(G237), .B2(G902), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n366), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n356), .B(new_n355), .C1(new_n343), .C2(new_n352), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n364), .B1(new_n385), .B2(new_n342), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n380), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G214), .B1(G237), .B2(G902), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT87), .Z(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n221), .ZN(new_n394));
  NOR2_X1   g208(.A1(G237), .A2(G953), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G214), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n207), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT94), .B1(new_n400), .B2(new_n205), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n400), .A2(new_n205), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G125), .ZN(new_n406));
  INV_X1    g220(.A(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G140), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n408), .A3(KEYINPUT16), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n407), .A2(KEYINPUT16), .A3(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(G146), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT74), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n396), .A2(new_n207), .ZN(new_n413));
  AOI21_X1  g227(.A(G143), .B1(new_n395), .B2(G214), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT17), .B(G131), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n205), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n410), .A3(new_n418), .A4(G146), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n412), .A2(new_n415), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n397), .A2(G131), .ZN(new_n422));
  OR3_X1    g236(.A1(new_n413), .A2(G131), .A3(new_n414), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI22_X1  g238(.A1(new_n420), .A2(new_n421), .B1(new_n424), .B2(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n421), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n394), .B(new_n404), .C1(new_n425), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT76), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n411), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n407), .A2(KEYINPUT16), .A3(G140), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n400), .B2(KEYINPUT16), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT76), .A3(G146), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n400), .B(KEYINPUT19), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n205), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n424), .A2(new_n430), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n404), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n394), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n428), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(G475), .A2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n392), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n392), .A3(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n404), .B1(new_n425), .B2(new_n427), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n438), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n428), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n191), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n443), .A2(new_n444), .B1(new_n448), .B2(G475), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n207), .A2(G128), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n207), .A2(KEYINPUT96), .A3(G128), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT96), .B1(new_n207), .B2(G128), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G134), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT96), .ZN(new_n456));
  INV_X1    g270(.A(G128), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(G143), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n207), .A2(KEYINPUT96), .A3(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n194), .A3(new_n451), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n320), .A2(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT67), .B(G116), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(G122), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n455), .A2(new_n461), .B1(new_n242), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n462), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n321), .A2(new_n323), .A3(G122), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(KEYINPUT14), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(KEYINPUT14), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT98), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT98), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n471), .A3(KEYINPUT14), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n465), .B1(new_n473), .B2(new_n223), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n450), .B1(new_n460), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n460), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n476), .A2(KEYINPUT97), .B1(KEYINPUT13), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT97), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT13), .B1(new_n458), .B2(new_n459), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n450), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n194), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n467), .A2(new_n466), .ZN(new_n483));
  INV_X1    g297(.A(new_n242), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n461), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n474), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G217), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n187), .A2(new_n488), .A3(G953), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n474), .B(new_n489), .C1(new_n482), .C2(new_n486), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n191), .ZN(new_n494));
  INV_X1    g308(.A(G478), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n494), .B(new_n496), .Z(new_n497));
  NAND2_X1  g311(.A1(new_n299), .A2(G952), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(G234), .B2(G237), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n191), .B(new_n299), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n449), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n391), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT22), .B(G137), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n417), .A2(new_n419), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n418), .B1(new_n432), .B2(G146), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT72), .B1(new_n314), .B2(G128), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT66), .B(G119), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(G128), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n515));
  AND4_X1   g329(.A1(new_n515), .A2(new_n315), .A3(new_n317), .A4(G128), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT24), .B(G110), .ZN(new_n518));
  OAI22_X1  g332(.A1(new_n510), .A2(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n513), .B2(G128), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(G128), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n457), .A2(KEYINPUT23), .A3(G119), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT73), .B1(new_n524), .B2(G110), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(KEYINPUT73), .A3(G110), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n400), .A2(new_n205), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n433), .A2(new_n430), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G110), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n521), .A2(new_n531), .A3(new_n522), .A4(new_n523), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n532), .A2(KEYINPUT75), .B1(new_n517), .B2(new_n518), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n509), .B1(new_n528), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  INV_X1    g351(.A(new_n530), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n517), .A2(new_n518), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n412), .A2(new_n417), .A3(new_n419), .ZN(new_n541));
  INV_X1    g355(.A(new_n527), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n525), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n543), .A3(new_n508), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n544), .A3(new_n191), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n488), .B1(G234), .B2(new_n191), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT25), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n550), .A2(G902), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n536), .A2(new_n544), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n536), .B2(new_n544), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n395), .A2(G210), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT27), .Z(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT28), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT64), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n196), .A2(G134), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n198), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(G131), .ZN(new_n567));
  AOI211_X1 g381(.A(KEYINPUT64), .B(new_n201), .C1(new_n565), .C2(new_n198), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n202), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT65), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n290), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT65), .B(new_n202), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n359), .B1(new_n202), .B2(new_n200), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n333), .A2(new_n330), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT69), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n569), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT69), .B(new_n202), .C1(new_n567), .C2(new_n568), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n254), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n203), .A2(new_n213), .A3(new_n219), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n330), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n563), .B1(new_n578), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n563), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n562), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT30), .B(new_n574), .C1(new_n571), .C2(new_n572), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n582), .B2(new_n583), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n577), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n562), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n587), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT31), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n582), .A2(new_n583), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n586), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(G134), .B(G137), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT64), .B1(new_n603), .B2(new_n201), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n566), .A2(new_n564), .A3(G131), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n201), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n254), .B1(new_n607), .B2(KEYINPUT65), .ZN(new_n608));
  INV_X1    g422(.A(new_n572), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n575), .B(new_n593), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n290), .B1(new_n569), .B2(new_n579), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n611), .A2(new_n581), .B1(new_n220), .B2(new_n203), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n612), .B2(new_n593), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n602), .B1(new_n613), .B2(new_n577), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT31), .B1(new_n614), .B2(new_n596), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n591), .B1(new_n599), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT32), .ZN(new_n617));
  NOR2_X1   g431(.A1(G472), .A2(G902), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n573), .A2(new_n575), .B1(new_n333), .B2(new_n330), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT28), .B1(new_n602), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n596), .B1(new_n621), .B2(new_n589), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n597), .A2(new_n598), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n614), .A2(KEYINPUT31), .A3(new_n596), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n618), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT32), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT71), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT29), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n562), .B1(new_n587), .B2(new_n563), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n588), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n614), .A2(new_n596), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT29), .B1(new_n621), .B2(new_n631), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(KEYINPUT71), .C1(new_n596), .C2(new_n614), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n600), .A2(new_n601), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n563), .B1(new_n638), .B2(new_n587), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n632), .A2(new_n639), .A3(new_n630), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n635), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(G472), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n558), .B1(new_n628), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n313), .A2(new_n505), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  NAND2_X1  g460(.A1(new_n298), .A2(new_n303), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n304), .A2(new_n306), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(G469), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n192), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n312), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n616), .B2(new_n191), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n625), .A2(new_n626), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n653), .A2(new_n558), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n189), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT99), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n313), .A2(KEYINPUT99), .A3(new_n655), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n389), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n383), .B2(new_n387), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n503), .ZN(new_n664));
  AOI21_X1  g478(.A(G478), .B1(new_n493), .B2(new_n191), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT33), .B1(new_n491), .B2(new_n492), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT33), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n487), .B2(new_n490), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n492), .A2(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n476), .A2(KEYINPUT97), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n477), .A2(KEYINPUT13), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n481), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G134), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n461), .A3(new_n485), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n674), .A2(new_n675), .A3(new_n474), .A4(new_n489), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n668), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n668), .A2(new_n669), .A3(new_n676), .A4(KEYINPUT101), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n666), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n495), .A2(G902), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n665), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n444), .ZN(new_n685));
  INV_X1    g499(.A(G475), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n446), .B2(new_n428), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n685), .A2(new_n442), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n684), .A2(KEYINPUT102), .A3(new_n688), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n664), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n661), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT34), .B(G104), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G6));
  NAND2_X1  g510(.A1(new_n388), .A2(new_n389), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n497), .A2(new_n688), .A3(new_n502), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n661), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT35), .B(G107), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G9));
  INV_X1    g517(.A(new_n553), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n539), .A2(new_n543), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT104), .B1(new_n509), .B2(KEYINPUT36), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT36), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n508), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n706), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n707), .A2(new_n706), .A3(new_n710), .ZN(new_n712));
  OR3_X1    g526(.A1(new_n705), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n705), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n704), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n550), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n716), .B1(new_n547), .B2(new_n548), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n715), .B1(new_n717), .B2(new_n551), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n653), .A2(new_n654), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n313), .A2(new_n505), .A3(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT37), .B(G110), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G12));
  INV_X1    g536(.A(G900), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n499), .B1(new_n500), .B2(new_n723), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n497), .A2(new_n688), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n651), .A2(new_n656), .A3(new_n725), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n627), .A2(new_n619), .B1(new_n642), .B2(G472), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n727), .A2(new_n697), .A3(new_n718), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G128), .ZN(G30));
  INV_X1    g544(.A(new_n597), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n596), .B1(new_n638), .B2(new_n587), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n191), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(G472), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n628), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n449), .A2(new_n497), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT38), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n382), .B1(new_n366), .B2(new_n381), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n386), .A2(new_n380), .A3(new_n384), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n383), .A2(new_n387), .A3(KEYINPUT38), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n718), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n737), .A2(new_n743), .A3(new_n662), .A4(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n724), .B(KEYINPUT39), .Z(new_n746));
  NAND2_X1  g560(.A1(new_n313), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT40), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT40), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n313), .A2(new_n749), .A3(new_n746), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G143), .ZN(G45));
  NOR3_X1   g566(.A1(new_n683), .A2(new_n449), .A3(new_n724), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n651), .A2(new_n656), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n728), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G146), .ZN(G48));
  AOI21_X1  g571(.A(new_n256), .B1(new_n285), .B2(new_n286), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT86), .B1(new_n758), .B2(new_n204), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n279), .A2(new_n280), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n306), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n761), .A2(new_n303), .B1(new_n304), .B2(new_n297), .ZN(new_n762));
  OAI21_X1  g576(.A(G469), .B1(new_n762), .B2(G902), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n188), .A3(new_n312), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n693), .A2(new_n644), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT41), .B(G113), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G15));
  NAND3_X1  g581(.A1(new_n764), .A2(new_n644), .A3(new_n700), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT105), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n764), .A2(KEYINPUT105), .A3(new_n700), .A4(new_n644), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  INV_X1    g587(.A(new_n504), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n728), .A2(new_n774), .A3(new_n764), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G119), .ZN(G21));
  NAND2_X1  g590(.A1(new_n623), .A2(new_n624), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n562), .B1(new_n639), .B2(new_n590), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n626), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(G472), .B1(new_n625), .B2(G902), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT106), .B(G472), .C1(new_n625), .C2(G902), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n558), .B(new_n779), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n736), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n697), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n764), .A3(new_n503), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G122), .ZN(G24));
  NAND2_X1  g602(.A1(new_n782), .A2(new_n783), .ZN(new_n789));
  INV_X1    g603(.A(new_n779), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n744), .A3(new_n753), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n763), .A2(new_n663), .A3(new_n188), .A4(new_n312), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G125), .ZN(G27));
  NAND4_X1  g610(.A1(new_n383), .A2(new_n387), .A3(new_n188), .A4(new_n389), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n644), .A2(new_n651), .A3(new_n753), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n797), .B1(new_n308), .B2(new_n312), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT42), .A3(new_n644), .A4(new_n753), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  AND3_X1   g619(.A1(new_n802), .A2(new_n644), .A3(new_n725), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n194), .ZN(G36));
  AND3_X1   g621(.A1(new_n647), .A2(KEYINPUT45), .A3(new_n648), .ZN(new_n808));
  OAI21_X1  g622(.A(G469), .B1(new_n307), .B2(KEYINPUT45), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n808), .B1(new_n809), .B2(KEYINPUT107), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT107), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(G469), .C1(new_n307), .C2(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n192), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n312), .B1(new_n813), .B2(KEYINPUT46), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n812), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n815), .A2(KEYINPUT46), .A3(new_n650), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n388), .A2(new_n662), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n653), .A2(new_n654), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n718), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n683), .B2(new_n688), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT108), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT43), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n682), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n666), .B(new_n828), .C1(new_n679), .C2(new_n680), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n449), .B(new_n827), .C1(new_n829), .C2(new_n665), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT44), .B1(new_n821), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n821), .A2(KEYINPUT44), .A3(new_n831), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT109), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n821), .A2(new_n835), .A3(KEYINPUT44), .A4(new_n831), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n819), .B(new_n832), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n817), .A2(new_n837), .A3(new_n188), .A4(new_n746), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G137), .ZN(G39));
  NAND4_X1  g653(.A1(new_n818), .A2(new_n727), .A3(new_n558), .A4(new_n753), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n188), .B1(new_n814), .B2(new_n816), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT47), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT47), .B(new_n188), .C1(new_n814), .C2(new_n816), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n840), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n405), .ZN(G42));
  INV_X1    g660(.A(G952), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n299), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT111), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n651), .A2(new_n798), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n791), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n718), .B(new_n779), .C1(new_n782), .C2(new_n783), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT111), .A3(new_n753), .A4(new_n802), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n628), .A2(new_n643), .ZN(new_n854));
  INV_X1    g668(.A(new_n724), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n449), .A2(new_n497), .A3(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n854), .A2(new_n818), .A3(new_n744), .A4(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n851), .A2(new_n853), .B1(new_n313), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n806), .B1(new_n801), .B2(new_n803), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g674(.A(KEYINPUT110), .B(new_n390), .C1(new_n739), .C2(new_n740), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n497), .A2(new_n688), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n861), .A2(new_n699), .B1(KEYINPUT110), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n689), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT110), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n391), .B2(new_n502), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n659), .A2(new_n864), .A3(new_n660), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n558), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n763), .A2(new_n188), .A3(new_n312), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT105), .B1(new_n871), .B2(new_n700), .ZN(new_n872));
  INV_X1    g686(.A(new_n771), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n867), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n313), .B(new_n505), .C1(new_n644), .C2(new_n719), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n765), .A2(new_n775), .A3(new_n787), .A4(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n860), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n792), .A2(new_n794), .B1(new_n726), .B2(new_n728), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n855), .A2(new_n188), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n881), .B(new_n715), .C1(new_n717), .C2(new_n551), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n388), .A2(new_n389), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n312), .B2(new_n308), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n785), .B1(new_n628), .B2(new_n734), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n755), .A2(new_n728), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n879), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n854), .A2(new_n663), .A3(new_n744), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n651), .A2(new_n656), .A3(new_n725), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n888), .A2(new_n889), .B1(new_n791), .B2(new_n793), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n651), .A2(new_n663), .A3(new_n882), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n888), .A2(new_n754), .B1(new_n891), .B2(new_n737), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT112), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n878), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n880), .A2(new_n886), .A3(new_n879), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT112), .B1(new_n890), .B2(new_n892), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT52), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n894), .A4(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT113), .ZN(new_n899));
  INV_X1    g713(.A(new_n866), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n689), .B2(new_n863), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n661), .A2(new_n901), .B1(new_n770), .B2(new_n771), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n765), .A2(new_n775), .A3(new_n787), .A4(new_n875), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n859), .A4(new_n858), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT52), .B1(new_n895), .B2(new_n896), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT53), .A4(new_n897), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT52), .B1(new_n890), .B2(new_n892), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n877), .A2(new_n894), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n899), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n874), .A2(new_n876), .ZN(new_n915));
  INV_X1    g729(.A(new_n860), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n894), .A2(new_n897), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n911), .ZN(new_n918));
  XOR2_X1   g732(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n919));
  NAND4_X1  g733(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n894), .A4(new_n909), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n819), .A2(new_n870), .ZN(new_n923));
  INV_X1    g737(.A(new_n499), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n824), .B2(new_n830), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n644), .A3(new_n925), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT48), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n691), .A2(new_n692), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n558), .A2(new_n924), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n628), .A2(new_n929), .A3(new_n734), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n923), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n847), .A2(G953), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n784), .A2(new_n925), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n931), .B(new_n932), .C1(new_n793), .C2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n763), .A2(new_n312), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n189), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n843), .A2(new_n844), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n933), .A2(new_n819), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n852), .A2(new_n764), .A3(new_n818), .A4(new_n925), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n684), .A2(new_n688), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n764), .A2(new_n930), .A3(new_n818), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n868), .A2(new_n944), .A3(new_n743), .A4(new_n925), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n763), .A2(new_n188), .A3(new_n312), .A4(new_n662), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(KEYINPUT115), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(KEYINPUT115), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n943), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT50), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n945), .B(new_n951), .C1(new_n947), .C2(new_n948), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n950), .A2(KEYINPUT51), .A3(new_n952), .ZN(new_n953));
  AOI211_X1 g767(.A(new_n927), .B(new_n934), .C1(new_n939), .C2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT117), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n956));
  INV_X1    g770(.A(new_n943), .ZN(new_n957));
  AND4_X1   g771(.A1(KEYINPUT116), .A2(new_n956), .A3(new_n952), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT116), .B1(new_n950), .B2(new_n952), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n939), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT51), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(KEYINPUT117), .B(KEYINPUT51), .C1(new_n939), .C2(new_n960), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n954), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n848), .B1(new_n922), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n935), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT49), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT49), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n868), .A2(new_n656), .A3(new_n390), .ZN(new_n970));
  NOR4_X1   g784(.A1(new_n735), .A2(new_n970), .A3(new_n688), .A4(new_n683), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n968), .A2(new_n743), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n966), .A2(new_n972), .ZN(G75));
  NAND2_X1  g787(.A1(new_n847), .A2(G953), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT118), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n918), .A2(new_n920), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(G210), .A3(G902), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT56), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n358), .B(new_n365), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT55), .Z(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n982), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n978), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n983), .B2(new_n985), .ZN(G51));
  XNOR2_X1  g800(.A(new_n192), .B(KEYINPUT57), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n762), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n815), .B(KEYINPUT119), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n977), .A2(G902), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n976), .B1(new_n992), .B2(new_n994), .ZN(G54));
  NAND4_X1  g809(.A1(new_n977), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n440), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n440), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n976), .B1(new_n997), .B2(new_n998), .ZN(G60));
  INV_X1    g813(.A(new_n681), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G478), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT59), .Z(new_n1002));
  NOR2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n988), .B2(new_n989), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n975), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1002), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT54), .ZN(new_n1007));
  AOI22_X1  g821(.A1(new_n898), .A2(KEYINPUT113), .B1(new_n910), .B2(new_n911), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1007), .B1(new_n1008), .B2(new_n908), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n1009), .B2(new_n988), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1005), .B1(new_n1000), .B2(new_n1010), .ZN(G63));
  NAND2_X1  g825(.A1(new_n713), .A2(new_n714), .ZN(new_n1012));
  NAND2_X1  g826(.A1(G217), .A2(G902), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT60), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n977), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n555), .A2(new_n556), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1014), .B1(new_n918), .B2(new_n920), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1016), .B(new_n975), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1018), .A2(new_n1017), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1023), .A2(new_n975), .A3(new_n1016), .A4(new_n1020), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(G66));
  NOR2_X1   g839(.A1(new_n915), .A2(G953), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT121), .ZN(new_n1027));
  INV_X1    g841(.A(G224), .ZN(new_n1028));
  OAI21_X1  g842(.A(G953), .B1(new_n501), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n385), .B(new_n342), .C1(G898), .C2(new_n299), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT122), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1030), .B(new_n1032), .ZN(G69));
  XNOR2_X1  g847(.A(new_n613), .B(new_n434), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n862), .B1(new_n684), .B2(new_n688), .ZN(new_n1035));
  OR4_X1    g849(.A1(new_n869), .A2(new_n747), .A3(new_n819), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n880), .A2(new_n756), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1038), .A2(new_n1039), .A3(new_n751), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n838), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n845), .ZN(new_n1042));
  INV_X1    g856(.A(new_n751), .ZN(new_n1043));
  OAI21_X1  g857(.A(KEYINPUT62), .B1(new_n1043), .B2(new_n1037), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(KEYINPUT123), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT123), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1046), .B(KEYINPUT62), .C1(new_n1043), .C2(new_n1037), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1041), .A2(new_n1042), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1034), .B1(new_n1049), .B2(new_n299), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1034), .B1(new_n723), .B2(new_n299), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n786), .A2(new_n644), .ZN(new_n1052));
  NAND4_X1  g866(.A1(new_n817), .A2(new_n188), .A3(new_n746), .A4(new_n1052), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n838), .A2(new_n1053), .A3(new_n859), .A4(new_n1038), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n1054), .A2(new_n845), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1051), .B1(new_n1055), .B2(new_n299), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n1050), .A2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g871(.A(KEYINPUT124), .B(KEYINPUT125), .Z(new_n1058));
  AOI21_X1  g872(.A(new_n299), .B1(G227), .B2(G900), .ZN(new_n1059));
  XNOR2_X1  g873(.A(new_n1058), .B(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g874(.A(new_n1057), .B(new_n1060), .ZN(G72));
  NAND4_X1  g875(.A1(new_n1041), .A2(new_n1042), .A3(new_n1048), .A4(new_n915), .ZN(new_n1062));
  NAND2_X1  g876(.A1(G472), .A2(G902), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1063), .B(KEYINPUT63), .Z(new_n1064));
  NAND2_X1  g878(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g879(.A(new_n614), .B(KEYINPUT126), .ZN(new_n1066));
  INV_X1    g880(.A(new_n1066), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n1067), .A2(new_n562), .ZN(new_n1068));
  AOI21_X1  g882(.A(KEYINPUT127), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g883(.A(KEYINPUT127), .ZN(new_n1070));
  INV_X1    g884(.A(new_n1068), .ZN(new_n1071));
  AOI211_X1 g885(.A(new_n1070), .B(new_n1071), .C1(new_n1062), .C2(new_n1064), .ZN(new_n1072));
  NOR2_X1   g886(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g887(.A(new_n913), .B(new_n1064), .C1(new_n634), .C2(new_n731), .ZN(new_n1074));
  INV_X1    g888(.A(new_n915), .ZN(new_n1075));
  NOR3_X1   g889(.A1(new_n1054), .A2(new_n845), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g890(.A(new_n1064), .ZN(new_n1077));
  OAI211_X1 g891(.A(new_n562), .B(new_n1067), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n1074), .A2(new_n975), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g893(.A1(new_n1073), .A2(new_n1079), .ZN(G57));
endmodule


