//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G58), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n204), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n228), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G50), .B(G68), .Z(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1698), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n252), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(G1698), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n254), .B1(new_n255), .B2(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G274), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT64), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT64), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n264), .A2(new_n266), .A3(new_n269), .A4(G274), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n260), .A2(new_n264), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n268), .A2(new_n270), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g0074(.A(KEYINPUT65), .B(G179), .Z(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(KEYINPUT66), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n217), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n221), .B1(new_n208), .B2(G20), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(new_n282), .B1(new_n221), .B2(new_n278), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n209), .B1(new_n201), .B2(new_n221), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n250), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI211_X1 g0089(.A(new_n284), .B(new_n288), .C1(G150), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n280), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n283), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n276), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n274), .A2(new_n275), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT66), .B1(new_n274), .B2(G169), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n273), .B2(G200), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n261), .A2(G190), .A3(new_n272), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT69), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n274), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n299), .A2(new_n307), .A3(new_n301), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n296), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n278), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT12), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n287), .B2(new_n255), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(KEYINPUT11), .A3(new_n280), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n208), .A2(G20), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n281), .A2(G68), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT11), .B1(new_n314), .B2(new_n280), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT13), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n268), .A2(new_n270), .B1(G238), .B2(new_n271), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n228), .A2(G1698), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  OAI221_X1 g0125(.A(new_n323), .B1(G226), .B2(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT71), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(new_n266), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n326), .A2(KEYINPUT71), .A3(new_n327), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n321), .B(new_n322), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(G190), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n330), .A2(new_n328), .A3(new_n266), .ZN(new_n333));
  INV_X1    g0133(.A(new_n322), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT13), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n320), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n331), .A3(KEYINPUT72), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(KEYINPUT13), .C1(new_n333), .C2(new_n334), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(G200), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(G169), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n337), .A2(new_n345), .A3(G169), .A4(new_n339), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n335), .A2(new_n331), .A3(G179), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n342), .B1(new_n348), .B2(new_n320), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n350));
  AOI21_X1  g0150(.A(new_n285), .B1(new_n208), .B2(G20), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n281), .B1(new_n278), .B2(new_n285), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n251), .A2(new_n209), .A3(new_n252), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n252), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT73), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(G68), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n227), .A2(new_n310), .ZN(new_n362));
  OAI21_X1  g0162(.A(G20), .B1(new_n362), .B2(new_n201), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n289), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT16), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n324), .A2(new_n325), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT7), .B1(new_n368), .B2(new_n209), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n369), .B2(new_n359), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n366), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n280), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n352), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n222), .A2(G1698), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(G223), .B2(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G87), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n375), .A2(new_n368), .B1(new_n250), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(new_n260), .B1(G232), .B2(new_n271), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n268), .A2(new_n270), .ZN(new_n379));
  AOI21_X1  g0179(.A(G200), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n350), .B1(new_n373), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n361), .A2(new_n366), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n355), .A2(new_n357), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n365), .B1(new_n388), .B2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n291), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n382), .B2(G200), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n391), .A2(new_n393), .A3(new_n352), .A4(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n384), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n352), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n387), .B2(new_n390), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n378), .A2(new_n379), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G169), .ZN(new_n402));
  INV_X1    g0202(.A(new_n275), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n378), .A2(new_n379), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(KEYINPUT18), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n404), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n373), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n398), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n271), .A2(G244), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n379), .A2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n253), .A2(G232), .B1(new_n368), .B2(G107), .ZN(new_n414));
  INV_X1    g0214(.A(G238), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n258), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n260), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n403), .ZN(new_n419));
  INV_X1    g0219(.A(G169), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n418), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT67), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n286), .ZN(new_n425));
  INV_X1    g0225(.A(new_n285), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n426), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n291), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n281), .A2(G77), .A3(new_n316), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G77), .B2(new_n277), .ZN(new_n430));
  OR3_X1    g0230(.A1(new_n428), .A2(KEYINPUT68), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT68), .B1(new_n428), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n421), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n413), .A2(new_n417), .A3(G190), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n418), .A2(G200), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n431), .A2(new_n432), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n309), .A2(new_n349), .A3(new_n411), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n209), .B(G87), .C1(new_n324), .C2(new_n325), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT22), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT22), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n256), .A2(new_n443), .A3(new_n209), .A4(G87), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT78), .B(G116), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n209), .A4(G33), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT78), .A2(G116), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT78), .A2(G116), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n209), .B(G33), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n209), .B2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n451), .A2(KEYINPUT83), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT24), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n454), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n458), .A2(new_n448), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n445), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n291), .B1(new_n457), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n250), .A2(G1), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n278), .A2(new_n280), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT25), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n277), .A2(new_n466), .A3(G107), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n277), .B2(G107), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n465), .A2(G107), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT84), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n461), .B1(new_n460), .B2(new_n445), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n461), .A2(new_n445), .A3(new_n448), .A4(new_n455), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n280), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT84), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n470), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n253), .A2(G250), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT85), .B(G294), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n260), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n263), .A2(G1), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n484), .A2(new_n266), .A3(G274), .A4(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n266), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G169), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n482), .A2(new_n260), .B1(new_n491), .B2(G264), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G179), .A3(new_n486), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n472), .A2(new_n477), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G190), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n493), .A2(G200), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n500), .A2(new_n475), .A3(new_n470), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(G33), .B1(new_n449), .B2(new_n450), .ZN(new_n504));
  INV_X1    g0304(.A(G244), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G1698), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G238), .B2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n507), .B2(new_n368), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n260), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n208), .A2(G45), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G250), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT77), .B1(new_n260), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n266), .A2(new_n513), .A3(G250), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G274), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n260), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n485), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT79), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT79), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n509), .A2(new_n515), .A3(new_n521), .A4(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(G190), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G200), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n520), .A2(KEYINPUT81), .A3(G190), .A4(new_n522), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n287), .B2(new_n204), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n256), .A2(new_n209), .A3(G68), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n209), .B1(new_n327), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G87), .B2(new_n206), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n280), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n422), .B(KEYINPUT67), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n278), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G87), .B2(new_n465), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n525), .A2(new_n527), .A3(new_n528), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n526), .A2(new_n420), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n424), .A2(new_n465), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n535), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n543), .A2(KEYINPUT80), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(KEYINPUT80), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n520), .A2(new_n275), .A3(new_n522), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n446), .A2(new_n277), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n465), .B2(G116), .ZN(new_n550));
  OR3_X1    g0350(.A1(new_n449), .A2(new_n450), .A3(new_n209), .ZN(new_n551));
  AOI21_X1  g0351(.A(G20), .B1(G33), .B2(G283), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n250), .A2(G97), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n552), .A2(new_n553), .B1(new_n279), .B2(new_n217), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n551), .A2(KEYINPUT20), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n486), .B1(new_n490), .B2(new_n224), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n486), .B(new_n560), .C1(new_n490), .C2(new_n224), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n562));
  INV_X1    g0362(.A(G1698), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n256), .A2(G257), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n368), .A2(G303), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n260), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n568), .B2(G200), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n381), .B2(new_n568), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .A4(new_n557), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n559), .A2(new_n561), .A3(new_n567), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G179), .A3(new_n557), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT21), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n557), .A2(G169), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n570), .A2(new_n571), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G244), .B(new_n563), .C1(new_n324), .C2(new_n325), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n563), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G283), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n260), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n486), .B1(new_n490), .B2(new_n229), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n420), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n584), .B2(new_n260), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n275), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT75), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(KEYINPUT6), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n593), .A2(new_n595), .B1(new_n204), .B2(G107), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(KEYINPUT6), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n206), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(G20), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n289), .A2(G77), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(KEYINPUT76), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT76), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n358), .A2(G107), .A3(new_n360), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n291), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n465), .A2(G97), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G97), .B2(new_n277), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n589), .B(new_n591), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n601), .A2(new_n602), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT76), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n601), .A2(KEYINPUT76), .A3(new_n602), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(new_n280), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n588), .A2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n590), .A2(G190), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n577), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n440), .A2(new_n503), .A3(new_n548), .A4(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n589), .A2(new_n591), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n540), .A2(new_n624), .A3(new_n547), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n519), .A2(G200), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n525), .A2(new_n528), .A3(new_n539), .A4(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n519), .A2(new_n420), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n628), .A2(new_n624), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n576), .A2(new_n571), .A3(new_n573), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n475), .A2(new_n470), .B1(new_n494), .B2(new_n496), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n610), .B(new_n619), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n628), .A2(new_n502), .A3(new_n631), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n440), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n410), .ZN(new_n641));
  INV_X1    g0441(.A(new_n434), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n348), .A2(new_n320), .B1(new_n341), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n398), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n306), .A2(new_n308), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n296), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(G369));
  INV_X1    g0447(.A(new_n634), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n557), .A2(new_n654), .ZN(new_n655));
  MUX2_X1   g0455(.A(new_n648), .B(new_n577), .S(new_n655), .Z(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n472), .A2(new_n477), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n654), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n503), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n498), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n648), .A2(new_n654), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n503), .A2(new_n666), .B1(new_n635), .B2(new_n662), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(G399));
  NOR3_X1   g0468(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  INV_X1    g0470(.A(new_n212), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n670), .A2(new_n208), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n216), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  NAND4_X1  g0475(.A1(new_n621), .A2(new_n503), .A3(new_n548), .A4(new_n662), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n572), .A2(G179), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n520), .A2(new_n495), .A3(new_n590), .A4(new_n522), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n499), .A2(new_n590), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n275), .A3(new_n519), .A4(new_n568), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n677), .B2(new_n678), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n654), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n654), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n676), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n620), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n628), .A2(new_n631), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n648), .A2(new_n498), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n693), .A2(new_n502), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n548), .A2(new_n629), .A3(new_n624), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT26), .B1(new_n694), .B2(new_n610), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n698), .A2(new_n631), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n654), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n639), .A2(new_n662), .ZN(new_n703));
  XNOR2_X1  g0503(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n691), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n675), .B1(new_n706), .B2(G1), .ZN(G364));
  INV_X1    g0507(.A(G13), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G20), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n208), .B1(new_n709), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n672), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n659), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(G330), .B2(new_n657), .ZN(new_n714));
  INV_X1    g0514(.A(new_n712), .ZN(new_n715));
  OR2_X1    g0515(.A1(G355), .A2(KEYINPUT90), .ZN(new_n716));
  NAND2_X1  g0516(.A1(G355), .A2(KEYINPUT90), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n212), .A3(new_n256), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n671), .A2(new_n256), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G45), .B2(new_n215), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n244), .A2(new_n263), .ZN(new_n721));
  OAI221_X1 g0521(.A(new_n718), .B1(G116), .B2(new_n212), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n217), .B1(G20), .B2(new_n420), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n715), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n209), .A2(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n381), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n256), .B1(new_n731), .B2(G283), .ZN(new_n732));
  INV_X1    g0532(.A(G303), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n480), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n381), .A2(G179), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n209), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n732), .B1(new_n733), .B2(new_n734), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n275), .A2(new_n209), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n381), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT92), .B(G326), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n740), .A2(G190), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT33), .B(G317), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n738), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n729), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT91), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G322), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n381), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n739), .A2(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n739), .A2(new_n748), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n757), .B1(G311), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n752), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  INV_X1    g0563(.A(new_n745), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n221), .A2(new_n742), .B1(new_n764), .B2(new_n310), .ZN(new_n765));
  INV_X1    g0565(.A(new_n734), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n766), .A2(G87), .B1(new_n731), .B2(G107), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n767), .B(new_n256), .C1(new_n204), .C2(new_n737), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n227), .A2(new_n756), .B1(new_n758), .B2(new_n255), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n747), .A2(new_n760), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n726), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n728), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  INV_X1    g0574(.A(new_n725), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n657), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n714), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(G396));
  NOR2_X1   g0578(.A1(new_n726), .A2(new_n723), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n715), .B1(new_n255), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n730), .A2(new_n376), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G107), .B2(new_n766), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n782), .B(new_n368), .C1(new_n204), .C2(new_n737), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(G283), .B2(new_n745), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n733), .B2(new_n742), .ZN(new_n785));
  INV_X1    g0585(.A(new_n752), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G311), .B1(new_n446), .B2(new_n759), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n756), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n756), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G159), .A2(new_n759), .B1(new_n791), .B2(G143), .ZN(new_n792));
  INV_X1    g0592(.A(G137), .ZN(new_n793));
  INV_X1    g0593(.A(G150), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n742), .B2(new_n793), .C1(new_n794), .C2(new_n764), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT34), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n256), .B1(new_n734), .B2(new_n221), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n737), .A2(new_n227), .B1(new_n730), .B2(new_n310), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(new_n786), .C2(G132), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n790), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n433), .A2(new_n654), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(new_n437), .B1(new_n433), .B2(new_n421), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n421), .A2(new_n433), .A3(new_n662), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n780), .B1(new_n800), .B2(new_n772), .C1(new_n805), .C2(new_n724), .ZN(new_n806));
  INV_X1    g0606(.A(new_n805), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n703), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n662), .B(new_n805), .C1(new_n633), .C2(new_n638), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(KEYINPUT94), .A3(new_n690), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n811), .B(new_n715), .C1(new_n690), .C2(new_n810), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT94), .B1(new_n810), .B2(new_n690), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n806), .B1(new_n812), .B2(new_n813), .ZN(G384));
  NOR2_X1   g0614(.A1(new_n709), .A2(new_n208), .ZN(new_n815));
  INV_X1    g0615(.A(G330), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT101), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n348), .A2(new_n320), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n320), .A2(new_n654), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n818), .A2(new_n341), .A3(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n320), .B(new_n654), .C1(new_n348), .C2(new_n342), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(new_n689), .A3(new_n805), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n389), .A2(KEYINPUT16), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n352), .B1(new_n372), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n652), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n398), .B2(new_n410), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n400), .A2(new_n393), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n825), .B1(new_n407), .B2(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n373), .A2(new_n407), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n373), .A2(new_n826), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n829), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n828), .A2(KEYINPUT38), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT97), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n828), .A2(new_n837), .A3(KEYINPUT97), .A4(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n828), .A2(new_n837), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n840), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n840), .A2(new_n844), .A3(KEYINPUT98), .A4(new_n841), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n823), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n817), .B1(new_n849), .B2(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(new_n823), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT38), .B1(new_n828), .B2(new_n837), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n839), .B2(new_n838), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT98), .B1(new_n853), .B2(new_n841), .ZN(new_n854));
  INV_X1    g0654(.A(new_n848), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(KEYINPUT101), .A3(new_n857), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n829), .A2(new_n833), .A3(new_n834), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n398), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n384), .A2(new_n397), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n641), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n834), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n859), .A2(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT38), .ZN(new_n871));
  INV_X1    g0671(.A(new_n838), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT40), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n850), .A2(new_n858), .B1(new_n851), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n440), .A2(new_n689), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n816), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n879), .B(new_n838), .C1(new_n870), .C2(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n818), .A2(new_n654), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n803), .B(KEYINPUT96), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n809), .A2(new_n885), .B1(new_n820), .B2(new_n821), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n854), .B2(new_n855), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n410), .A2(new_n652), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n702), .A2(new_n440), .A3(new_n705), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n646), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n889), .B(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n815), .B1(new_n878), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n892), .B2(new_n878), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n596), .A2(KEYINPUT35), .A3(new_n600), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(G116), .A3(new_n218), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT35), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n596), .A2(new_n600), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n899), .A2(KEYINPUT36), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(KEYINPUT36), .ZN(new_n901));
  OAI21_X1  g0701(.A(G77), .B1(new_n227), .B2(new_n310), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n215), .A2(new_n902), .B1(G50), .B2(new_n310), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n708), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT95), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n894), .A2(new_n900), .A3(new_n901), .A4(new_n905), .ZN(G367));
  OAI21_X1  g0706(.A(new_n654), .B1(new_n607), .B2(new_n609), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n693), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n624), .A2(new_n654), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n503), .A2(new_n666), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT42), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n908), .A2(new_n498), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n662), .B1(new_n914), .B2(new_n624), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n911), .A2(KEYINPUT42), .A3(new_n912), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT43), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n539), .A2(new_n662), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n631), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n695), .B2(new_n919), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT102), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n916), .A2(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n918), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n665), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n910), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n672), .B(KEYINPUT41), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n910), .A2(new_n667), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT45), .Z(new_n931));
  NOR2_X1   g0731(.A1(new_n910), .A2(new_n667), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n926), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n926), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n912), .B1(new_n664), .B2(new_n666), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n658), .B2(KEYINPUT103), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n940), .B(new_n941), .Z(new_n942));
  NAND3_X1  g0742(.A1(new_n938), .A2(new_n706), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(new_n943), .B2(new_n706), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n710), .B1(new_n944), .B2(KEYINPUT104), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n928), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n922), .A2(new_n725), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n786), .A2(G317), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n756), .A2(new_n733), .ZN(new_n950));
  INV_X1    g0750(.A(G283), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n758), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT46), .B1(new_n766), .B2(new_n446), .ZN(new_n953));
  NOR4_X1   g0753(.A1(new_n949), .A2(new_n950), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n368), .B1(new_n737), .B2(new_n205), .ZN(new_n955));
  NAND2_X1  g0755(.A1(KEYINPUT46), .A2(G116), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n730), .A2(new_n204), .B1(new_n734), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(KEYINPUT105), .B(G311), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n955), .B(new_n957), .C1(new_n741), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n954), .B(new_n960), .C1(new_n735), .C2(new_n764), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n737), .A2(new_n310), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G77), .B2(new_n731), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n963), .B(new_n256), .C1(new_n227), .C2(new_n734), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G159), .B2(new_n745), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n752), .A2(new_n793), .B1(new_n794), .B2(new_n756), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G50), .B2(new_n759), .ZN(new_n967));
  INV_X1    g0767(.A(G143), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n965), .B(new_n967), .C1(new_n968), .C2(new_n742), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n726), .ZN(new_n972));
  INV_X1    g0772(.A(new_n719), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n727), .B1(new_n212), .B2(new_n536), .C1(new_n973), .C2(new_n240), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n948), .A2(new_n712), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n947), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT106), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(G387));
  NAND2_X1  g0778(.A1(new_n942), .A2(new_n711), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n664), .A2(new_n775), .ZN(new_n980));
  INV_X1    g0780(.A(new_n737), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n981), .A2(G283), .B1(new_n766), .B2(new_n480), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G303), .A2(new_n759), .B1(new_n791), .B2(G317), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n742), .B2(new_n754), .C1(new_n764), .C2(new_n958), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT48), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT49), .Z(new_n990));
  INV_X1    g0790(.A(new_n446), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n368), .B1(new_n991), .B2(new_n730), .C1(new_n752), .C2(new_n743), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n256), .B1(new_n730), .B2(new_n204), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G77), .B2(new_n766), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n742), .B2(new_n761), .C1(new_n285), .C2(new_n764), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n424), .A2(new_n981), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT109), .B(G150), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n752), .B2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n221), .A2(new_n756), .B1(new_n758), .B2(new_n310), .ZN(new_n1000));
  NOR3_X1   g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n726), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n670), .A2(new_n212), .A3(new_n256), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(G107), .B2(new_n212), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT107), .ZN(new_n1005));
  AOI211_X1 g0805(.A(G45), .B(new_n670), .C1(G68), .C2(G77), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n285), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n719), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n237), .A2(G45), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1005), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n715), .B1(new_n1013), .B2(new_n727), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1002), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n942), .A2(new_n706), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n672), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n942), .A2(new_n706), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n979), .B1(new_n980), .B2(new_n1015), .C1(new_n1017), .C2(new_n1018), .ZN(G393));
  OAI21_X1  g0819(.A(new_n1016), .B1(new_n936), .B2(new_n937), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n943), .A2(new_n672), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n911), .A2(new_n725), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n727), .B1(new_n204), .B2(new_n212), .C1(new_n973), .C2(new_n247), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n712), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n741), .A2(G317), .B1(new_n791), .B2(G311), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n759), .A2(G294), .B1(new_n446), .B2(new_n981), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n733), .C2(new_n764), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n256), .B1(new_n731), .B2(G107), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n951), .B2(new_n734), .C1(new_n752), .C2(new_n754), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  AOI22_X1  g0831(.A1(new_n741), .A2(G150), .B1(new_n791), .B2(G159), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT51), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n752), .A2(new_n968), .B1(new_n310), .B2(new_n734), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n745), .A2(G50), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n759), .A2(new_n426), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n737), .A2(new_n255), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1038), .A2(new_n781), .A3(new_n368), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1028), .A2(new_n1031), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1024), .B1(new_n1041), .B2(new_n726), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n938), .A2(new_n711), .B1(new_n1022), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1021), .A2(new_n1043), .ZN(G390));
  NAND2_X1  g0844(.A1(new_n809), .A2(new_n885), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n822), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n883), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(KEYINPUT113), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT113), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n886), .B2(new_n883), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1048), .A2(new_n1050), .A3(new_n881), .A4(new_n880), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n863), .A2(new_n859), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n410), .B1(KEYINPUT100), .B2(new_n866), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n834), .B1(new_n1053), .B2(new_n865), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n843), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n883), .B1(new_n1055), .B2(new_n838), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n802), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n804), .B1(new_n701), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n822), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1051), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n691), .A2(new_n805), .A3(new_n822), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1051), .A2(new_n1062), .A3(new_n1060), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n691), .A2(new_n440), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n890), .A2(new_n646), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1059), .B1(new_n690), .B2(new_n807), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n1045), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1062), .A2(new_n1058), .A3(new_n1069), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1064), .A2(new_n1065), .A3(new_n1073), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1075), .A2(new_n672), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n779), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n712), .B1(new_n1078), .B2(new_n426), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n998), .A2(new_n734), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT53), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G137), .B2(new_n745), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n791), .A2(G132), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT54), .B(G143), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n786), .A2(G125), .B1(new_n759), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n256), .B1(new_n730), .B2(new_n221), .C1(new_n737), .C2(new_n761), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n741), .B2(G128), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n752), .A2(new_n788), .B1(new_n310), .B2(new_n730), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT114), .Z(new_n1090));
  AOI22_X1  g0890(.A1(G107), .A2(new_n745), .B1(new_n741), .B2(G283), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n256), .B(new_n1038), .C1(G87), .C2(new_n766), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G97), .A2(new_n759), .B1(new_n791), .B2(G116), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1088), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1079), .B1(new_n1095), .B2(new_n726), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n882), .B2(new_n724), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1066), .B2(new_n710), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1077), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G378));
  INV_X1    g0900(.A(new_n889), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT120), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n889), .A2(KEYINPUT120), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n292), .A2(new_n826), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n309), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n309), .A2(new_n1105), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n850), .A2(new_n858), .ZN(new_n1113));
  OAI21_X1  g0913(.A(G330), .B1(new_n873), .B2(new_n823), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1111), .B(new_n1114), .C1(new_n850), .C2(new_n858), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1103), .B(new_n1104), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT101), .B1(new_n856), .B2(new_n857), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n849), .A2(new_n817), .A3(KEYINPUT40), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1111), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1113), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n1102), .A3(new_n1123), .A4(new_n1101), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT57), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1068), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1076), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1051), .A2(new_n1062), .A3(new_n1060), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1062), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1068), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n889), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1135), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1122), .A2(new_n1123), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1133), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n672), .B(new_n1128), .C1(new_n1139), .C2(KEYINPUT57), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n731), .A2(G58), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT115), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n742), .B2(new_n223), .C1(new_n204), .C2(new_n764), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n368), .A2(new_n262), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1144), .B(new_n962), .C1(G77), .C2(new_n766), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1145), .B1(new_n951), .B2(new_n752), .C1(new_n536), .C2(new_n758), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n791), .A2(G107), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT116), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT117), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(KEYINPUT58), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1144), .B(new_n221), .C1(G33), .C2(G41), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n766), .A2(new_n1084), .ZN(new_n1153));
  INV_X1    g0953(.A(G128), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1153), .B1(new_n794), .B2(new_n737), .C1(new_n756), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n741), .A2(G125), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n764), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1155), .B(new_n1158), .C1(G137), .C2(new_n759), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1160), .A2(KEYINPUT59), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n731), .C2(G159), .ZN(new_n1162));
  INV_X1    g0962(.A(G124), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n752), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT118), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT59), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1159), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1151), .B(new_n1152), .C1(new_n1161), .C2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1150), .A2(KEYINPUT58), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n726), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n715), .B1(new_n221), .B2(new_n779), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1170), .B(new_n1171), .C1(new_n1111), .C2(new_n724), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n711), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1140), .A2(new_n1175), .ZN(G375));
  NAND2_X1  g0976(.A1(new_n1059), .A2(new_n723), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n712), .B1(new_n1078), .B2(G68), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n752), .A2(new_n1154), .B1(new_n794), .B2(new_n758), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G137), .B2(new_n791), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n256), .B1(new_n737), .B2(new_n221), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G159), .B2(new_n766), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G132), .A2(new_n741), .B1(new_n745), .B2(new_n1084), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1142), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n741), .A2(G294), .B1(new_n759), .B2(G107), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n991), .B2(new_n764), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT122), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n997), .B1(new_n951), .B2(new_n756), .C1(new_n752), .C2(new_n733), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n368), .B1(new_n730), .B2(new_n255), .C1(new_n204), .C2(new_n734), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1178), .B1(new_n1191), .B2(new_n726), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1132), .A2(new_n711), .B1(new_n1177), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n929), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1074), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1071), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT121), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1071), .A2(new_n1068), .A3(KEYINPUT121), .A4(new_n1072), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1193), .B1(new_n1195), .B2(new_n1200), .ZN(G381));
  INV_X1    g1001(.A(G375), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(G393), .A2(G396), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1204), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n977), .A2(new_n1099), .A3(new_n1202), .A4(new_n1205), .ZN(G407));
  NAND2_X1  g1006(.A1(new_n653), .A2(G213), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1202), .A2(new_n1099), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(G407), .A2(G213), .A3(new_n1209), .ZN(G409));
  INV_X1    g1010(.A(KEYINPUT60), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1073), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n672), .B1(new_n1200), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1071), .A2(new_n1068), .A3(KEYINPUT60), .A4(new_n1072), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT124), .ZN(new_n1215));
  OAI21_X1  g1015(.A(KEYINPUT125), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT124), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1214), .B(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1198), .B(new_n1199), .C1(new_n1211), .C2(new_n1073), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT125), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n672), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT126), .ZN(new_n1223));
  OR2_X1    g1023(.A1(G384), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1193), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(G384), .A2(new_n1223), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1225), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1228), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1076), .A2(new_n1126), .ZN(new_n1234));
  NOR3_X1   g1034(.A1(new_n1116), .A2(new_n1117), .A3(new_n1135), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1137), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1194), .B(new_n1234), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1118), .A2(new_n1124), .A3(new_n711), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1172), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1099), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1140), .A2(G378), .A3(new_n1175), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1240), .B1(new_n1239), .B2(new_n1099), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1207), .B(new_n1233), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT62), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1239), .A2(new_n1099), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT123), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1250), .A2(KEYINPUT62), .A3(new_n1207), .A4(new_n1233), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1207), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1229), .A2(new_n1232), .B1(G2897), .B2(new_n1208), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1225), .B(new_n1228), .C1(new_n1216), .C2(new_n1221), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1208), .A2(G2897), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1254), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1252), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT127), .ZN(new_n1262));
  AND2_X1   g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  OAI21_X1  g1063(.A(G390), .B1(new_n1263), .B2(new_n1203), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1203), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT106), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(G390), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n976), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1252), .A2(new_n1260), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1245), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(KEYINPUT63), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(KEYINPUT63), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(new_n1268), .A3(new_n1275), .A4(new_n1260), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G375), .A2(new_n1099), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1242), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1279), .B(new_n1233), .Z(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1268), .ZN(G402));
endmodule


