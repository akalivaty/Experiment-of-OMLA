

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744;

  NOR2_X1 U372 ( .A1(n560), .A2(n589), .ZN(n704) );
  XNOR2_X2 U373 ( .A(n349), .B(n405), .ZN(n459) );
  XNOR2_X2 U374 ( .A(n404), .B(G110), .ZN(n349) );
  NOR2_X1 U375 ( .A1(n566), .A2(n513), .ZN(n703) );
  BUF_X1 U376 ( .A(G104), .Z(n675) );
  NAND2_X1 U377 ( .A1(n693), .A2(n709), .ZN(n371) );
  AND2_X2 U378 ( .A1(n492), .A2(n600), .ZN(n382) );
  XNOR2_X2 U379 ( .A(n420), .B(n419), .ZN(n559) );
  OR2_X2 U380 ( .A1(n649), .A2(n644), .ZN(n420) );
  NOR2_X2 U381 ( .A1(n744), .A2(n743), .ZN(n549) );
  NAND2_X2 U382 ( .A1(n594), .A2(n357), .ZN(n378) );
  XNOR2_X2 U383 ( .A(n379), .B(n362), .ZN(n594) );
  XNOR2_X2 U384 ( .A(n555), .B(n421), .ZN(n537) );
  XNOR2_X1 U385 ( .A(n544), .B(KEYINPUT1), .ZN(n495) );
  XNOR2_X1 U386 ( .A(n424), .B(n423), .ZN(n483) );
  INV_X1 U387 ( .A(KEYINPUT64), .ZN(n411) );
  OR2_X1 U388 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  AND2_X1 U389 ( .A1(n579), .A2(n703), .ZN(n539) );
  OR2_X1 U390 ( .A1(n546), .A2(n560), .ZN(n547) );
  XNOR2_X1 U391 ( .A(n616), .B(n615), .ZN(n709) );
  INV_X1 U392 ( .A(n495), .ZN(n600) );
  AND2_X1 U393 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U394 ( .A(n394), .B(n393), .ZN(n727) );
  XNOR2_X1 U395 ( .A(n732), .B(n460), .ZN(n718) );
  XNOR2_X1 U396 ( .A(n431), .B(n415), .ZN(n455) );
  XNOR2_X1 U397 ( .A(n411), .B(G953), .ZN(n456) );
  NOR2_X2 U398 ( .A1(n536), .A2(n535), .ZN(n568) );
  XNOR2_X1 U399 ( .A(n604), .B(n603), .ZN(n350) );
  XNOR2_X1 U400 ( .A(n604), .B(n603), .ZN(n678) );
  NAND2_X1 U401 ( .A1(n380), .A2(n602), .ZN(n604) );
  INV_X1 U402 ( .A(n397), .ZN(n351) );
  XNOR2_X2 U403 ( .A(n472), .B(n353), .ZN(n732) );
  OR2_X1 U404 ( .A1(n611), .A2(n360), .ZN(n693) );
  INV_X1 U405 ( .A(KEYINPUT79), .ZN(n391) );
  XNOR2_X1 U406 ( .A(n389), .B(KEYINPUT77), .ZN(n388) );
  NAND2_X1 U407 ( .A1(n701), .A2(n570), .ZN(n389) );
  NAND2_X1 U408 ( .A1(n371), .A2(n354), .ZN(n370) );
  NAND2_X1 U409 ( .A1(n461), .A2(G902), .ZN(n375) );
  XNOR2_X1 U410 ( .A(n383), .B(G140), .ZN(n479) );
  INV_X1 U411 ( .A(G137), .ZN(n383) );
  XNOR2_X1 U412 ( .A(n412), .B(n413), .ZN(n368) );
  XNOR2_X1 U413 ( .A(n459), .B(n407), .ZN(n364) );
  XOR2_X1 U414 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n481) );
  XOR2_X1 U415 ( .A(G122), .B(G107), .Z(n426) );
  XNOR2_X1 U416 ( .A(n448), .B(n447), .ZN(n686) );
  XNOR2_X1 U417 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U418 ( .A1(n384), .A2(n545), .ZN(n560) );
  XNOR2_X1 U419 ( .A(n385), .B(KEYINPUT28), .ZN(n384) );
  AND2_X1 U420 ( .A1(n550), .A2(n612), .ZN(n385) );
  XNOR2_X1 U421 ( .A(n487), .B(KEYINPUT25), .ZN(n488) );
  BUF_X1 U422 ( .A(n456), .Z(n735) );
  INV_X1 U423 ( .A(KEYINPUT78), .ZN(n386) );
  NAND2_X1 U424 ( .A1(n397), .A2(n356), .ZN(n396) );
  XNOR2_X1 U425 ( .A(n370), .B(n617), .ZN(n622) );
  XNOR2_X1 U426 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U427 ( .A(G143), .B(G140), .ZN(n443) );
  NAND2_X2 U428 ( .A1(n374), .A2(n372), .ZN(n544) );
  NAND2_X1 U429 ( .A1(G469), .A2(n473), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n455), .B(n454), .ZN(n472) );
  INV_X1 U431 ( .A(KEYINPUT82), .ZN(n639) );
  XNOR2_X1 U432 ( .A(n366), .B(n455), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n367), .B(n414), .ZN(n366) );
  XNOR2_X1 U434 ( .A(n451), .B(n450), .ZN(n566) );
  XNOR2_X1 U435 ( .A(n449), .B(G475), .ZN(n450) );
  XNOR2_X1 U436 ( .A(n598), .B(n597), .ZN(n607) );
  XNOR2_X1 U437 ( .A(n369), .B(KEYINPUT93), .ZN(n611) );
  XNOR2_X1 U438 ( .A(n484), .B(n355), .ZN(n394) );
  XNOR2_X1 U439 ( .A(n482), .B(n731), .ZN(n393) );
  XNOR2_X1 U440 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U441 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U442 ( .A(KEYINPUT88), .B(n654), .Z(n715) );
  AND2_X1 U443 ( .A1(n697), .A2(KEYINPUT44), .ZN(n352) );
  XNOR2_X1 U444 ( .A(n359), .B(n488), .ZN(n497) );
  XOR2_X1 U445 ( .A(n479), .B(KEYINPUT94), .Z(n353) );
  XOR2_X1 U446 ( .A(n569), .B(KEYINPUT80), .Z(n354) );
  XOR2_X1 U447 ( .A(n481), .B(n480), .Z(n355) );
  AND2_X1 U448 ( .A1(n350), .A2(n352), .ZN(n356) );
  XOR2_X1 U449 ( .A(n593), .B(KEYINPUT92), .Z(n357) );
  NOR2_X1 U450 ( .A1(n591), .A2(n668), .ZN(n358) );
  NOR2_X1 U451 ( .A1(n727), .A2(G902), .ZN(n359) );
  OR2_X1 U452 ( .A1(n613), .A2(n612), .ZN(n360) );
  XOR2_X1 U453 ( .A(KEYINPUT87), .B(KEYINPUT33), .Z(n361) );
  XOR2_X1 U454 ( .A(KEYINPUT75), .B(KEYINPUT19), .Z(n362) );
  XNOR2_X1 U455 ( .A(n364), .B(n469), .ZN(n667) );
  AND2_X1 U456 ( .A1(n401), .A2(n399), .ZN(n398) );
  BUF_X1 U457 ( .A(n722), .Z(n726) );
  BUF_X1 U458 ( .A(n607), .Z(n363) );
  BUF_X1 U459 ( .A(n638), .Z(n662) );
  INV_X1 U460 ( .A(KEYINPUT44), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n667), .B(n365), .ZN(n649) );
  INV_X1 U462 ( .A(n368), .ZN(n367) );
  NAND2_X1 U463 ( .A1(n369), .A2(n614), .ZN(n616) );
  NAND2_X1 U464 ( .A1(n369), .A2(n596), .ZN(n598) );
  XNOR2_X2 U465 ( .A(n378), .B(n595), .ZN(n369) );
  INV_X1 U466 ( .A(n676), .ZN(n397) );
  NAND2_X1 U467 ( .A1(n676), .A2(n402), .ZN(n401) );
  XNOR2_X2 U468 ( .A(n403), .B(KEYINPUT35), .ZN(n676) );
  OR2_X1 U469 ( .A1(n718), .A2(n373), .ZN(n372) );
  NAND2_X1 U470 ( .A1(n718), .A2(n461), .ZN(n376) );
  XNOR2_X2 U471 ( .A(n377), .B(G128), .ZN(n431) );
  XNOR2_X2 U472 ( .A(KEYINPUT65), .B(G143), .ZN(n377) );
  NAND2_X1 U473 ( .A1(n559), .A2(n558), .ZN(n379) );
  NAND2_X1 U474 ( .A1(n380), .A2(n618), .ZN(n620) );
  AND2_X2 U475 ( .A1(n607), .A2(n599), .ZN(n380) );
  XNOR2_X1 U476 ( .A(n381), .B(KEYINPUT34), .ZN(n610) );
  NOR2_X2 U477 ( .A1(n608), .A2(n611), .ZN(n381) );
  XNOR2_X2 U478 ( .A(n382), .B(n361), .ZN(n608) );
  XNOR2_X1 U479 ( .A(n387), .B(n386), .ZN(n571) );
  NAND2_X1 U480 ( .A1(n390), .A2(n388), .ZN(n387) );
  XNOR2_X1 U481 ( .A(n392), .B(n391), .ZN(n390) );
  NAND2_X1 U482 ( .A1(n564), .A2(KEYINPUT47), .ZN(n392) );
  INV_X1 U483 ( .A(n594), .ZN(n589) );
  NAND2_X1 U484 ( .A1(n398), .A2(n396), .ZN(n626) );
  NAND2_X1 U485 ( .A1(n400), .A2(n402), .ZN(n399) );
  NAND2_X1 U486 ( .A1(n678), .A2(n697), .ZN(n400) );
  NAND2_X1 U487 ( .A1(n610), .A2(n609), .ZN(n403) );
  XNOR2_X1 U488 ( .A(n628), .B(n627), .ZN(n638) );
  XNOR2_X2 U489 ( .A(n476), .B(n475), .ZN(n612) );
  BUF_X1 U490 ( .A(n649), .Z(n651) );
  INV_X1 U491 ( .A(KEYINPUT69), .ZN(n573) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U493 ( .A(KEYINPUT8), .ZN(n423) );
  NOR2_X1 U494 ( .A1(n580), .A2(n582), .ZN(n556) );
  BUF_X1 U495 ( .A(n495), .Z(n618) );
  INV_X1 U496 ( .A(KEYINPUT56), .ZN(n656) );
  XNOR2_X2 U497 ( .A(G107), .B(G104), .ZN(n404) );
  XNOR2_X1 U498 ( .A(G101), .B(KEYINPUT74), .ZN(n405) );
  XNOR2_X1 U499 ( .A(KEYINPUT72), .B(KEYINPUT16), .ZN(n406) );
  XNOR2_X1 U500 ( .A(n406), .B(G122), .ZN(n407) );
  XNOR2_X1 U501 ( .A(G116), .B(G113), .ZN(n408) );
  XNOR2_X1 U502 ( .A(n408), .B(KEYINPUT3), .ZN(n410) );
  XOR2_X1 U503 ( .A(KEYINPUT71), .B(G119), .Z(n409) );
  XNOR2_X1 U504 ( .A(n410), .B(n409), .ZN(n469) );
  XOR2_X1 U505 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n413) );
  NAND2_X1 U506 ( .A1(n456), .A2(G224), .ZN(n412) );
  XNOR2_X1 U507 ( .A(G146), .B(G125), .ZN(n441) );
  XNOR2_X1 U508 ( .A(n441), .B(KEYINPUT17), .ZN(n414) );
  XNOR2_X1 U509 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n415) );
  XNOR2_X1 U510 ( .A(G902), .B(KEYINPUT15), .ZN(n485) );
  INV_X1 U511 ( .A(n485), .ZN(n644) );
  INV_X1 U512 ( .A(G902), .ZN(n473) );
  INV_X1 U513 ( .A(G237), .ZN(n416) );
  NAND2_X1 U514 ( .A1(n473), .A2(n416), .ZN(n422) );
  NAND2_X1 U515 ( .A1(n422), .A2(G210), .ZN(n418) );
  INV_X1 U516 ( .A(KEYINPUT90), .ZN(n417) );
  XNOR2_X1 U517 ( .A(n418), .B(n417), .ZN(n419) );
  BUF_X1 U518 ( .A(n559), .Z(n555) );
  XNOR2_X1 U519 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n421) );
  NAND2_X1 U520 ( .A1(n422), .A2(G214), .ZN(n558) );
  NAND2_X1 U521 ( .A1(n537), .A2(n558), .ZN(n514) );
  NAND2_X1 U522 ( .A1(n456), .A2(G234), .ZN(n424) );
  NAND2_X1 U523 ( .A1(G217), .A2(n483), .ZN(n430) );
  XNOR2_X1 U524 ( .A(G116), .B(G134), .ZN(n425) );
  XNOR2_X1 U525 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U526 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n427) );
  XNOR2_X1 U527 ( .A(n432), .B(n431), .ZN(n724) );
  NAND2_X1 U528 ( .A1(n724), .A2(n473), .ZN(n434) );
  XNOR2_X1 U529 ( .A(KEYINPUT103), .B(G478), .ZN(n433) );
  XNOR2_X1 U530 ( .A(n434), .B(n433), .ZN(n565) );
  XOR2_X1 U531 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n436) );
  XNOR2_X1 U532 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n435) );
  XNOR2_X1 U533 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U534 ( .A(G113), .B(G131), .Z(n438) );
  INV_X1 U535 ( .A(KEYINPUT102), .ZN(n437) );
  XNOR2_X1 U536 ( .A(KEYINPUT10), .B(n441), .ZN(n731) );
  XNOR2_X1 U537 ( .A(n442), .B(n731), .ZN(n448) );
  XOR2_X1 U538 ( .A(G122), .B(n675), .Z(n444) );
  XNOR2_X1 U539 ( .A(n444), .B(n443), .ZN(n446) );
  NOR2_X1 U540 ( .A1(G953), .A2(G237), .ZN(n462) );
  NAND2_X1 U541 ( .A1(G214), .A2(n462), .ZN(n445) );
  NOR2_X1 U542 ( .A1(G902), .A2(n686), .ZN(n451) );
  INV_X1 U543 ( .A(KEYINPUT13), .ZN(n449) );
  AND2_X1 U544 ( .A1(n565), .A2(n566), .ZN(n587) );
  INV_X1 U545 ( .A(n587), .ZN(n512) );
  NOR2_X1 U546 ( .A1(n514), .A2(n512), .ZN(n453) );
  XNOR2_X1 U547 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n453), .B(n452), .ZN(n546) );
  BUF_X1 U549 ( .A(n546), .Z(n510) );
  XNOR2_X1 U550 ( .A(G134), .B(G131), .ZN(n454) );
  NAND2_X1 U551 ( .A1(n735), .A2(G227), .ZN(n457) );
  XNOR2_X1 U552 ( .A(n457), .B(G146), .ZN(n458) );
  XNOR2_X1 U553 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U554 ( .A(G469), .ZN(n461) );
  XOR2_X1 U555 ( .A(KEYINPUT98), .B(G137), .Z(n464) );
  NAND2_X1 U556 ( .A1(n462), .A2(G210), .ZN(n463) );
  XNOR2_X1 U557 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U558 ( .A(G101), .B(G146), .Z(n466) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n465) );
  XNOR2_X1 U560 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U561 ( .A(n468), .B(n467), .Z(n470) );
  XNOR2_X1 U562 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U563 ( .A(n472), .B(n471), .ZN(n680) );
  NAND2_X1 U564 ( .A1(n680), .A2(n473), .ZN(n476) );
  INV_X1 U565 ( .A(KEYINPUT99), .ZN(n474) );
  XNOR2_X1 U566 ( .A(n474), .B(G472), .ZN(n475) );
  XNOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT6), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n612), .B(n477), .ZN(n599) );
  XNOR2_X1 U569 ( .A(G119), .B(G128), .ZN(n478) );
  XNOR2_X1 U570 ( .A(n479), .B(n478), .ZN(n482) );
  XNOR2_X1 U571 ( .A(G110), .B(KEYINPUT95), .ZN(n480) );
  NAND2_X1 U572 ( .A1(G221), .A2(n483), .ZN(n484) );
  NAND2_X1 U573 ( .A1(n485), .A2(G234), .ZN(n486) );
  XNOR2_X1 U574 ( .A(n486), .B(KEYINPUT20), .ZN(n489) );
  NAND2_X1 U575 ( .A1(G217), .A2(n489), .ZN(n487) );
  NAND2_X1 U576 ( .A1(n489), .A2(G221), .ZN(n491) );
  XOR2_X1 U577 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n490) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n586) );
  AND2_X1 U579 ( .A1(n497), .A2(n586), .ZN(n504) );
  INV_X1 U580 ( .A(n504), .ZN(n523) );
  NOR2_X1 U581 ( .A1(n599), .A2(n523), .ZN(n492) );
  NOR2_X1 U582 ( .A1(n510), .A2(n608), .ZN(n493) );
  NOR2_X1 U583 ( .A1(n493), .A2(G953), .ZN(n635) );
  NAND2_X1 U584 ( .A1(G234), .A2(G237), .ZN(n494) );
  XNOR2_X1 U585 ( .A(n494), .B(KEYINPUT14), .ZN(n525) );
  NAND2_X1 U586 ( .A1(G952), .A2(n525), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n618), .A2(n523), .ZN(n496) );
  XNOR2_X1 U588 ( .A(n496), .B(KEYINPUT50), .ZN(n503) );
  INV_X1 U589 ( .A(n497), .ZN(n601) );
  NOR2_X1 U590 ( .A1(n586), .A2(n497), .ZN(n498) );
  XNOR2_X1 U591 ( .A(n498), .B(KEYINPUT49), .ZN(n500) );
  INV_X1 U592 ( .A(n612), .ZN(n499) );
  NAND2_X1 U593 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U594 ( .A(KEYINPUT121), .B(n501), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n503), .A2(n502), .ZN(n507) );
  AND2_X1 U596 ( .A1(n612), .A2(n504), .ZN(n505) );
  AND2_X1 U597 ( .A1(n600), .A2(n505), .ZN(n614) );
  INV_X1 U598 ( .A(n614), .ZN(n506) );
  NAND2_X1 U599 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U600 ( .A(KEYINPUT51), .B(n508), .ZN(n509) );
  NOR2_X1 U601 ( .A1(n510), .A2(n509), .ZN(n520) );
  NOR2_X1 U602 ( .A1(n537), .A2(n558), .ZN(n511) );
  NOR2_X1 U603 ( .A1(n512), .A2(n511), .ZN(n516) );
  INV_X1 U604 ( .A(n565), .ZN(n513) );
  AND2_X1 U605 ( .A1(n566), .A2(n513), .ZN(n692) );
  XNOR2_X1 U606 ( .A(n692), .B(KEYINPUT104), .ZN(n578) );
  NOR2_X1 U607 ( .A1(n578), .A2(n703), .ZN(n569) );
  NOR2_X1 U608 ( .A1(n569), .A2(n514), .ZN(n515) );
  NOR2_X1 U609 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U610 ( .A(n517), .B(KEYINPUT122), .ZN(n518) );
  NOR2_X1 U611 ( .A1(n518), .A2(n608), .ZN(n519) );
  NOR2_X1 U612 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U613 ( .A(n521), .B(KEYINPUT52), .ZN(n522) );
  NOR2_X1 U614 ( .A1(n529), .A2(n522), .ZN(n633) );
  OR2_X2 U615 ( .A1(n523), .A2(n544), .ZN(n613) );
  XNOR2_X1 U616 ( .A(KEYINPUT110), .B(n613), .ZN(n536) );
  NAND2_X1 U617 ( .A1(n612), .A2(n558), .ZN(n524) );
  XOR2_X1 U618 ( .A(KEYINPUT30), .B(n524), .Z(n534) );
  NAND2_X1 U619 ( .A1(G902), .A2(n525), .ZN(n591) );
  NOR2_X1 U620 ( .A1(G900), .A2(n591), .ZN(n527) );
  INV_X1 U621 ( .A(n735), .ZN(n526) );
  NAND2_X1 U622 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U623 ( .A(KEYINPUT109), .B(n528), .ZN(n531) );
  NOR2_X1 U624 ( .A1(G953), .A2(n529), .ZN(n530) );
  XOR2_X1 U625 ( .A(KEYINPUT91), .B(n530), .Z(n592) );
  NOR2_X1 U626 ( .A1(n531), .A2(n592), .ZN(n532) );
  XNOR2_X1 U627 ( .A(n532), .B(KEYINPUT76), .ZN(n540) );
  INV_X1 U628 ( .A(n540), .ZN(n533) );
  NAND2_X1 U629 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U630 ( .A1(n568), .A2(n537), .ZN(n538) );
  XNOR2_X1 U631 ( .A(n538), .B(KEYINPUT39), .ZN(n579) );
  XNOR2_X1 U632 ( .A(KEYINPUT40), .B(n539), .ZN(n744) );
  INV_X1 U633 ( .A(n586), .ZN(n541) );
  NOR2_X1 U634 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(n542), .Z(n543) );
  NOR2_X1 U636 ( .A1(n497), .A2(n543), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n544), .B(KEYINPUT111), .ZN(n545) );
  XNOR2_X1 U638 ( .A(KEYINPUT113), .B(n547), .ZN(n548) );
  XNOR2_X1 U639 ( .A(KEYINPUT42), .B(n548), .ZN(n743) );
  XNOR2_X1 U640 ( .A(n549), .B(KEYINPUT46), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n703), .A2(n550), .ZN(n552) );
  INV_X1 U642 ( .A(n558), .ZN(n551) );
  NOR2_X1 U643 ( .A1(n552), .A2(n551), .ZN(n554) );
  INV_X1 U644 ( .A(n599), .ZN(n553) );
  NAND2_X1 U645 ( .A1(n554), .A2(n553), .ZN(n580) );
  INV_X1 U646 ( .A(n555), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n556), .B(KEYINPUT36), .ZN(n557) );
  NAND2_X1 U648 ( .A1(n557), .A2(n600), .ZN(n712) );
  XNOR2_X1 U649 ( .A(KEYINPUT85), .B(n712), .ZN(n563) );
  NAND2_X1 U650 ( .A1(n354), .A2(n704), .ZN(n561) );
  NOR2_X1 U651 ( .A1(KEYINPUT47), .A2(n561), .ZN(n562) );
  NOR2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n572) );
  INV_X1 U653 ( .A(n704), .ZN(n564) );
  NOR2_X1 U654 ( .A1(n566), .A2(n565), .ZN(n609) );
  AND2_X1 U655 ( .A1(n555), .A2(n609), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n568), .A2(n567), .ZN(n701) );
  NAND2_X1 U657 ( .A1(KEYINPUT47), .A2(n569), .ZN(n570) );
  AND2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U659 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U660 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U661 ( .A(n577), .B(KEYINPUT48), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n579), .A2(n578), .ZN(n714) );
  OR2_X1 U663 ( .A1(n580), .A2(n600), .ZN(n581) );
  XNOR2_X1 U664 ( .A(n581), .B(KEYINPUT43), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n583), .A2(n582), .ZN(n660) );
  NAND2_X1 U666 ( .A1(n714), .A2(n660), .ZN(n584) );
  NOR2_X2 U667 ( .A1(n585), .A2(n584), .ZN(n734) );
  NAND2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U669 ( .A(n588), .B(KEYINPUT107), .ZN(n596) );
  INV_X1 U670 ( .A(G898), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n590), .A2(G953), .ZN(n668) );
  NOR2_X1 U672 ( .A1(n592), .A2(n358), .ZN(n593) );
  INV_X1 U673 ( .A(KEYINPUT0), .ZN(n595) );
  INV_X1 U674 ( .A(KEYINPUT22), .ZN(n597) );
  AND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U676 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n612), .A2(n497), .ZN(n605) );
  AND2_X1 U678 ( .A1(n618), .A2(n605), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n363), .A2(n606), .ZN(n697) );
  INV_X1 U680 ( .A(KEYINPUT31), .ZN(n615) );
  INV_X1 U681 ( .A(KEYINPUT105), .ZN(n617) );
  INV_X1 U682 ( .A(KEYINPUT86), .ZN(n619) );
  XNOR2_X1 U683 ( .A(n620), .B(n619), .ZN(n621) );
  NAND2_X1 U684 ( .A1(n621), .A2(n497), .ZN(n677) );
  NAND2_X1 U685 ( .A1(n622), .A2(n677), .ZN(n624) );
  INV_X1 U686 ( .A(KEYINPUT108), .ZN(n623) );
  XNOR2_X1 U687 ( .A(n624), .B(n623), .ZN(n625) );
  NAND2_X1 U688 ( .A1(n626), .A2(n625), .ZN(n628) );
  XNOR2_X1 U689 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n627) );
  AND2_X1 U690 ( .A1(n734), .A2(n662), .ZN(n629) );
  NAND2_X1 U691 ( .A1(n629), .A2(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U692 ( .A1(n630), .A2(n647), .ZN(n631) );
  XNOR2_X1 U693 ( .A(KEYINPUT83), .B(n631), .ZN(n632) );
  NOR2_X1 U694 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U695 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U696 ( .A(KEYINPUT53), .B(n636), .ZN(n637) );
  INV_X1 U697 ( .A(n637), .ZN(G75) );
  NAND2_X1 U698 ( .A1(n638), .A2(n644), .ZN(n640) );
  XNOR2_X1 U699 ( .A(n640), .B(n639), .ZN(n641) );
  NAND2_X1 U700 ( .A1(n641), .A2(n734), .ZN(n643) );
  INV_X1 U701 ( .A(KEYINPUT81), .ZN(n642) );
  XNOR2_X1 U702 ( .A(n643), .B(n642), .ZN(n646) );
  NAND2_X1 U703 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U704 ( .A1(n646), .A2(n645), .ZN(n648) );
  AND2_X2 U705 ( .A1(n648), .A2(n647), .ZN(n722) );
  NAND2_X1 U706 ( .A1(n722), .A2(G210), .ZN(n653) );
  XNOR2_X1 U707 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U708 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U709 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X1 U710 ( .A1(n735), .A2(G952), .ZN(n654) );
  NAND2_X1 U711 ( .A1(n655), .A2(n715), .ZN(n657) );
  XNOR2_X1 U712 ( .A(n657), .B(n656), .ZN(G51) );
  XOR2_X1 U713 ( .A(G113), .B(KEYINPUT119), .Z(n659) );
  INV_X1 U714 ( .A(n703), .ZN(n673) );
  NOR2_X1 U715 ( .A1(n709), .A2(n673), .ZN(n658) );
  XOR2_X1 U716 ( .A(n659), .B(n658), .Z(G15) );
  XNOR2_X1 U717 ( .A(n660), .B(G140), .ZN(G42) );
  INV_X1 U718 ( .A(G953), .ZN(n661) );
  NAND2_X1 U719 ( .A1(n662), .A2(n661), .ZN(n666) );
  NAND2_X1 U720 ( .A1(G953), .A2(G224), .ZN(n663) );
  XNOR2_X1 U721 ( .A(KEYINPUT61), .B(n663), .ZN(n664) );
  NAND2_X1 U722 ( .A1(n664), .A2(G898), .ZN(n665) );
  NAND2_X1 U723 ( .A1(n666), .A2(n665), .ZN(n672) );
  INV_X1 U724 ( .A(n667), .ZN(n669) );
  NAND2_X1 U725 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U726 ( .A(n670), .B(KEYINPUT125), .ZN(n671) );
  XNOR2_X1 U727 ( .A(n672), .B(n671), .ZN(G69) );
  NOR2_X1 U728 ( .A1(n693), .A2(n673), .ZN(n674) );
  XOR2_X1 U729 ( .A(n675), .B(n674), .Z(G6) );
  XOR2_X1 U730 ( .A(n351), .B(G122), .Z(G24) );
  XNOR2_X1 U731 ( .A(n677), .B(G101), .ZN(G3) );
  XNOR2_X1 U732 ( .A(n350), .B(G119), .ZN(G21) );
  NAND2_X1 U733 ( .A1(n722), .A2(G472), .ZN(n682) );
  XNOR2_X1 U734 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U736 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U737 ( .A1(n683), .A2(n715), .ZN(n684) );
  XNOR2_X1 U738 ( .A(n684), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U739 ( .A1(n722), .A2(G475), .ZN(n688) );
  XNOR2_X1 U740 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n685) );
  XNOR2_X1 U741 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n688), .B(n687), .ZN(n689) );
  NAND2_X1 U743 ( .A1(n689), .A2(n715), .ZN(n691) );
  XNOR2_X1 U744 ( .A(KEYINPUT67), .B(KEYINPUT60), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(G60) );
  XOR2_X1 U746 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n695) );
  INV_X1 U747 ( .A(n692), .ZN(n708) );
  NOR2_X1 U748 ( .A1(n693), .A2(n708), .ZN(n694) );
  XOR2_X1 U749 ( .A(n695), .B(n694), .Z(n696) );
  XNOR2_X1 U750 ( .A(G107), .B(n696), .ZN(G9) );
  XNOR2_X1 U751 ( .A(G110), .B(n697), .ZN(G12) );
  XOR2_X1 U752 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n699) );
  NAND2_X1 U753 ( .A1(n704), .A2(n692), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U755 ( .A(G128), .B(n700), .Z(G30) );
  XNOR2_X1 U756 ( .A(G143), .B(KEYINPUT116), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n702), .B(n701), .ZN(G45) );
  XOR2_X1 U758 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n706) );
  NAND2_X1 U759 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U761 ( .A(G146), .B(n707), .ZN(G48) );
  NOR2_X1 U762 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U763 ( .A(KEYINPUT120), .B(n710), .Z(n711) );
  XNOR2_X1 U764 ( .A(G116), .B(n711), .ZN(G18) );
  XOR2_X1 U765 ( .A(n712), .B(G125), .Z(n713) );
  XNOR2_X1 U766 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U767 ( .A(G134), .B(n714), .ZN(G36) );
  INV_X1 U768 ( .A(n715), .ZN(n730) );
  NAND2_X1 U769 ( .A1(n726), .A2(G469), .ZN(n720) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n716), .B(KEYINPUT57), .ZN(n717) );
  XNOR2_X1 U772 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U773 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U774 ( .A1(n730), .A2(n721), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n722), .A2(G478), .ZN(n723) );
  XOR2_X1 U776 ( .A(n724), .B(n723), .Z(n725) );
  NOR2_X1 U777 ( .A1(n730), .A2(n725), .ZN(G63) );
  NAND2_X1 U778 ( .A1(n726), .A2(G217), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(G66) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT126), .ZN(n733) );
  XOR2_X1 U782 ( .A(n733), .B(n732), .Z(n737) );
  XNOR2_X1 U783 ( .A(n734), .B(n737), .ZN(n736) );
  NAND2_X1 U784 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U785 ( .A(G227), .B(n737), .Z(n738) );
  NAND2_X1 U786 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U787 ( .A1(G953), .A2(n739), .ZN(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n742), .Z(G72) );
  XOR2_X1 U790 ( .A(G137), .B(n743), .Z(G39) );
  XOR2_X1 U791 ( .A(G131), .B(n744), .Z(G33) );
endmodule

