//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n206), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(KEYINPUT70), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(KEYINPUT10), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n218), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n210), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT67), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n256), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n201), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n210), .B1(new_n262), .B2(new_n202), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n210), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n254), .ZN(new_n267));
  INV_X1    g0067(.A(G50), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n209), .B2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(new_n269), .B1(new_n268), .B2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n264), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(G274), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT3), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n288));
  AND3_X1   g0088(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT66), .ZN(new_n289));
  AOI21_X1  g0089(.A(KEYINPUT66), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G222), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(G223), .A3(G1698), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n293), .B(new_n294), .C1(new_n228), .C2(new_n291), .ZN(new_n295));
  INV_X1    g0095(.A(new_n279), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n272), .A2(new_n274), .B1(new_n297), .B2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n252), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n251), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n271), .B1(new_n297), .B2(G169), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n297), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n298), .A2(new_n301), .A3(new_n251), .A4(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT18), .ZN(new_n313));
  OR2_X1    g0113(.A1(G223), .A2(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n281), .A2(G1698), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n286), .A2(new_n314), .A3(new_n288), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G87), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n296), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n280), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(KEYINPUT75), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n279), .B1(new_n316), .B2(new_n317), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n280), .A2(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n324), .A2(new_n325), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n327), .A2(new_n328), .B1(new_n307), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n222), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n332), .B2(new_n202), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n259), .A2(G159), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n286), .A2(new_n288), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n210), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(G68), .ZN(new_n339));
  AOI21_X1  g0139(.A(G20), .B1(new_n286), .B2(new_n288), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n337), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(KEYINPUT16), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n254), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT74), .B1(new_n285), .B2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n285), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n285), .A2(KEYINPUT74), .A3(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n210), .B1(new_n289), .B2(new_n290), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n337), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n335), .B1(new_n351), .B2(new_n222), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT16), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n257), .B1(new_n209), .B2(G20), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n267), .B1(new_n266), .B2(new_n257), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n313), .B(new_n330), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n254), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n333), .A2(new_n334), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n346), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n222), .B1(new_n340), .B2(new_n337), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n360), .B1(new_n366), .B2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n286), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n288), .A3(new_n348), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT66), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n362), .B2(new_n346), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT66), .ZN(new_n374));
  AOI21_X1  g0174(.A(G20), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n371), .B1(new_n375), .B2(KEYINPUT7), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n361), .B1(new_n376), .B2(G68), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n367), .B1(new_n377), .B2(KEYINPUT16), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n356), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n313), .B1(new_n379), .B2(new_n330), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n359), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT75), .B1(new_n319), .B2(new_n321), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n324), .A2(new_n325), .A3(new_n323), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n299), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n324), .A2(new_n325), .A3(G190), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n378), .A2(new_n387), .A3(new_n356), .ZN(new_n388));
  NOR2_X1   g0188(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n389));
  NAND2_X1  g0189(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n378), .A2(new_n387), .A3(new_n356), .A4(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n228), .B1(new_n209), .B2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n267), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n266), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n397), .B1(G77), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n257), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n255), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n399), .B1(new_n403), .B2(new_n254), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n291), .A2(G232), .A3(new_n292), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n291), .A2(G238), .A3(G1698), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n373), .A2(new_n374), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G107), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n296), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n280), .B1(new_n229), .B2(new_n283), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n404), .B1(new_n413), .B2(new_n328), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n409), .B2(new_n296), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n307), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT69), .B1(new_n415), .B2(new_n307), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(G190), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n404), .C1(new_n299), .C2(new_n415), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OR3_X1    g0221(.A1(new_n312), .A2(new_n395), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n259), .A2(G50), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT72), .B1(new_n210), .B2(G68), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n425), .B1(new_n426), .B2(new_n423), .C1(new_n256), .C2(new_n228), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT73), .B1(new_n427), .B2(new_n254), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT11), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT11), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n428), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n398), .A2(KEYINPUT12), .A3(G68), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT12), .B1(new_n398), .B2(G68), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n222), .B1(new_n209), .B2(G20), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n435), .A2(new_n436), .B1(new_n267), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n291), .A2(KEYINPUT71), .A3(G226), .A4(new_n292), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n373), .A2(G226), .A3(new_n292), .A4(new_n374), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G97), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n441), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n296), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n280), .B1(new_n223), .B2(new_n283), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT13), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT13), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n453), .A3(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n440), .B1(new_n455), .B2(G169), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n448), .B2(new_n450), .ZN(new_n457));
  AOI211_X1 g0257(.A(KEYINPUT13), .B(new_n449), .C1(new_n447), .C2(new_n296), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n440), .B(G169), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n452), .A2(G179), .A3(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n439), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n439), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(G190), .A3(new_n454), .ZN(new_n464));
  OAI21_X1  g0264(.A(G200), .B1(new_n457), .B2(new_n458), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n422), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n209), .A2(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NAND2_X1  g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n473), .A2(new_n296), .A3(new_n230), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n225), .A2(new_n292), .ZN(new_n475));
  INV_X1    g0275(.A(G257), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G1698), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n286), .A2(new_n475), .A3(new_n288), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G294), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n279), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  AND2_X1   g0281(.A1(G1), .A2(G13), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(new_n278), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n474), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(KEYINPUT84), .A3(G179), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT84), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(new_n470), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G264), .A3(new_n279), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n473), .A2(new_n483), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n478), .A2(new_n479), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n279), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n487), .B1(new_n494), .B2(new_n307), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n480), .A2(new_n484), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n328), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n486), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n486), .B(new_n500), .C1(new_n495), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT25), .B1(new_n266), .B2(new_n206), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n287), .A2(G1), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n266), .A2(new_n254), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n504), .A2(new_n505), .B1(new_n507), .B2(G107), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n286), .A2(new_n288), .A3(new_n210), .A4(G87), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT22), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n511), .B1(new_n510), .B2(KEYINPUT22), .ZN(new_n513));
  OR3_X1    g0313(.A1(new_n224), .A2(KEYINPUT22), .A3(G20), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n512), .A2(new_n513), .B1(new_n407), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n210), .B2(G107), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n517), .A2(new_n518), .B1(new_n520), .B2(new_n210), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT83), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(KEYINPUT24), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n524), .B1(new_n515), .B2(new_n521), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n360), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n509), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n502), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n529), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n494), .A2(new_n299), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G190), .B2(new_n494), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n532), .A2(new_n508), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT86), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(new_n534), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT86), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n537), .B(new_n538), .C1(new_n530), .C2(new_n502), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT20), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n210), .B1(new_n205), .B2(G33), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G283), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT77), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT77), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(G33), .A3(G283), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n253), .A2(new_n218), .B1(G20), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n540), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n543), .A2(new_n545), .ZN(new_n551));
  OAI211_X1 g0351(.A(KEYINPUT20), .B(new_n548), .C1(new_n551), .C2(new_n541), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n398), .A2(G116), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n507), .B2(G116), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n328), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(G303), .B1(new_n289), .B2(new_n290), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n230), .A2(G1698), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G257), .B2(G1698), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n559), .A2(new_n336), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n279), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n490), .A2(new_n279), .ZN(new_n562));
  INV_X1    g0362(.A(G270), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n492), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(KEYINPUT81), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n373), .B2(new_n374), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n559), .A2(new_n336), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n296), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n473), .A2(new_n296), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(G270), .B1(new_n483), .B2(new_n473), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n556), .A2(new_n565), .A3(KEYINPUT21), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n553), .A2(new_n555), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n575), .A2(G179), .A3(new_n569), .A4(new_n572), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n575), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n565), .A2(new_n573), .A3(G200), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT81), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n570), .B1(new_n569), .B2(new_n572), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G190), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n578), .B(new_n579), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n556), .A2(new_n565), .A3(new_n573), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n577), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n373), .A2(G250), .A3(G1698), .A4(new_n374), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n229), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n373), .A2(new_n292), .A3(new_n374), .A4(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n286), .A2(new_n288), .A3(G244), .A4(new_n292), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n590), .B1(new_n545), .B2(new_n543), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n589), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n296), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n571), .A2(G257), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(new_n492), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n398), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n507), .B2(G97), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT6), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n603), .A2(new_n205), .A3(G107), .ZN(new_n604));
  XNOR2_X1  g0404(.A(G97), .B(G107), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n606), .A2(new_n210), .B1(new_n228), .B2(new_n260), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n351), .B2(new_n206), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n602), .B1(new_n609), .B2(new_n254), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n595), .A2(new_n296), .B1(G257), .B2(new_n571), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(G190), .A3(new_n492), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n599), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n598), .A2(new_n328), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n607), .B1(new_n376), .B2(G107), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n601), .B1(new_n615), .B2(new_n360), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n307), .A3(new_n492), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n210), .B1(new_n446), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(G87), .B2(new_n207), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n286), .A2(new_n288), .A3(new_n210), .A4(G68), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT79), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(new_n620), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n624), .B2(new_n620), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n622), .B(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n254), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n402), .A2(new_n266), .ZN(new_n630));
  INV_X1    g0430(.A(new_n402), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n507), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n483), .A2(new_n489), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT78), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n636), .A2(new_n209), .A3(G45), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n635), .A2(G250), .A3(new_n279), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(G238), .A2(G1698), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n229), .B2(G1698), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n520), .B1(new_n363), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n634), .B(new_n638), .C1(new_n641), .C2(new_n279), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n328), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n638), .A2(new_n634), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n223), .A2(new_n292), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n229), .A2(G1698), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n286), .A2(new_n645), .A3(new_n288), .A4(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n279), .B1(new_n647), .B2(new_n519), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n307), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n633), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n648), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(G190), .A3(new_n634), .A4(new_n638), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n628), .A2(new_n254), .B1(new_n266), .B2(new_n402), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n507), .A2(G87), .ZN(new_n655));
  OAI21_X1  g0455(.A(G200), .B1(new_n644), .B2(new_n648), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n651), .A2(KEYINPUT80), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT80), .B1(new_n651), .B2(new_n657), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n588), .A2(new_n619), .A3(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n469), .A2(new_n536), .A3(new_n539), .A4(new_n661), .ZN(G372));
  AND2_X1   g0462(.A1(new_n613), .A2(new_n618), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n657), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n537), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n530), .A2(new_n498), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n577), .A2(new_n668), .A3(new_n587), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT21), .B1(new_n582), .B2(new_n556), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n574), .A2(new_n576), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT87), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT26), .B1(new_n660), .B2(new_n618), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n618), .A2(new_n664), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n651), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n469), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n310), .ZN(new_n681));
  INV_X1    g0481(.A(new_n418), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n457), .A2(new_n458), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT14), .B1(new_n683), .B2(new_n328), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n460), .A3(new_n459), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n467), .A2(new_n682), .B1(new_n685), .B2(new_n439), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n391), .A2(new_n389), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n352), .A2(new_n353), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n357), .B1(new_n688), .B2(new_n367), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n687), .B1(new_n689), .B2(new_n387), .ZN(new_n690));
  INV_X1    g0490(.A(new_n393), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n381), .B1(new_n686), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n304), .A2(new_n311), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n681), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n680), .A2(new_n695), .ZN(G369));
  INV_X1    g0496(.A(KEYINPUT88), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n588), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n575), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n588), .A2(new_n697), .ZN(new_n707));
  INV_X1    g0507(.A(new_n673), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n706), .A2(new_n707), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n704), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n536), .B(new_n539), .C1(new_n530), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n531), .A2(new_n704), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n667), .A2(new_n704), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n670), .A2(new_n671), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(new_n704), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n536), .A2(new_n539), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n716), .A2(new_n717), .A3(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n213), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT89), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n727), .B1(new_n216), .B2(new_n724), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n727), .B2(new_n726), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND4_X1  g0530(.A1(new_n536), .A2(new_n661), .A3(new_n539), .A4(new_n712), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n569), .A2(G179), .A3(new_n572), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT90), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n494), .A2(new_n642), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n569), .A2(KEYINPUT90), .A3(new_n572), .A4(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n734), .A2(new_n611), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n611), .A2(new_n735), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n734), .A4(new_n736), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n596), .A2(new_n492), .A3(new_n597), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n649), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n565), .A2(new_n573), .A3(new_n494), .A4(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n739), .B(new_n741), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n712), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT91), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n744), .B2(new_n742), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n485), .A2(G179), .A3(new_n649), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n582), .A2(KEYINPUT91), .A3(new_n598), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n739), .A2(new_n741), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n753), .B2(new_n704), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n710), .B1(new_n731), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n712), .B1(new_n674), .B2(new_n679), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT92), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n531), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n666), .B1(new_n761), .B2(new_n718), .ZN(new_n762));
  OR3_X1    g0562(.A1(new_n660), .A2(KEYINPUT26), .A3(new_n618), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT26), .B1(new_n618), .B2(new_n664), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n651), .A3(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT29), .B(new_n712), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n673), .A2(new_n667), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n535), .A2(new_n619), .A3(new_n664), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND3_X1   g0570(.A1(new_n675), .A2(new_n651), .A3(new_n678), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n704), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT92), .B1(new_n772), .B2(KEYINPUT29), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n756), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n730), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(new_n265), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n209), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n723), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n711), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n709), .A2(new_n710), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT95), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n709), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n291), .A2(G355), .A3(new_n213), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G116), .B2(new_n213), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n213), .A2(new_n336), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n276), .B2(new_n217), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n246), .A2(G45), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n218), .B1(G20), .B2(new_n328), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n786), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n779), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n583), .A2(new_n299), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n210), .A2(G179), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n407), .B1(new_n566), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  NAND2_X1  g0604(.A1(G20), .A2(G179), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n800), .ZN(new_n807));
  INV_X1    g0607(.A(G326), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n801), .A2(new_n583), .A3(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n801), .A2(new_n583), .A3(new_n299), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n811), .A2(G283), .B1(new_n813), .B2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(G294), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n583), .A2(G200), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n210), .B1(new_n816), .B2(new_n307), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n806), .A2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n809), .B(new_n818), .C1(G322), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n806), .A2(new_n583), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G200), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n299), .ZN(new_n824));
  XNOR2_X1  g0624(.A(KEYINPUT33), .B(G317), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT101), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G311), .A2(new_n823), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n804), .A2(new_n821), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n824), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n222), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n817), .B(KEYINPUT99), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n205), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n830), .B(new_n833), .C1(G77), .C2(new_n823), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n813), .A2(G159), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n820), .A2(G58), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n810), .A2(new_n206), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n802), .A2(new_n224), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n407), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT98), .ZN(new_n843));
  INV_X1    g0643(.A(new_n807), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n839), .B(new_n843), .C1(G50), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n828), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n799), .B1(new_n847), .B2(new_n796), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n787), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n782), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(G396));
  INV_X1    g0651(.A(KEYINPUT104), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n418), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n404), .A2(new_n712), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n420), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n414), .B(KEYINPUT104), .C1(new_n416), .C2(new_n417), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n772), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n682), .A2(new_n704), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n772), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n756), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n779), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n864), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n784), .A2(new_n796), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n779), .B1(new_n868), .B2(G77), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n833), .B1(G116), .B2(new_n823), .ZN(new_n870));
  INV_X1    g0670(.A(new_n802), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n811), .A2(G87), .B1(new_n871), .B2(G107), .ZN(new_n872));
  INV_X1    g0672(.A(G311), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(new_n812), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n815), .A2(new_n819), .B1(new_n807), .B2(new_n566), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n874), .A2(new_n291), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(G283), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n870), .B(new_n876), .C1(new_n877), .C2(new_n829), .ZN(new_n878));
  AOI22_X1  g0678(.A1(G137), .A2(new_n844), .B1(new_n820), .B2(G143), .ZN(new_n879));
  INV_X1    g0679(.A(new_n823), .ZN(new_n880));
  INV_X1    g0680(.A(G159), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .C1(new_n258), .C2(new_n829), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(new_n817), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G58), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n336), .B1(new_n871), .B2(G50), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n810), .A2(new_n222), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(G132), .B2(new_n813), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n883), .A2(KEYINPUT34), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n869), .B1(new_n892), .B2(new_n796), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT103), .Z(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n785), .B2(new_n862), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n866), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G384));
  NOR2_X1   g0697(.A1(new_n776), .A2(new_n209), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n366), .A2(KEYINPUT16), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n356), .B1(new_n343), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n702), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n381), .B2(new_n394), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n330), .B2(new_n901), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n388), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT107), .B1(new_n689), .B2(new_n702), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n379), .A2(new_n908), .A3(new_n901), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n330), .B1(new_n354), .B2(new_n357), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n904), .A3(new_n388), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n903), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n910), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n385), .B1(new_n327), .B2(new_n299), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n354), .A2(new_n917), .A3(new_n357), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT109), .B(new_n393), .C1(new_n918), .C2(new_n687), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n911), .A2(KEYINPUT18), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n358), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT109), .B1(new_n392), .B2(new_n393), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n911), .A2(new_n388), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT108), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n907), .B2(new_n909), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n904), .B2(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n910), .A2(new_n926), .A3(KEYINPUT37), .A4(new_n924), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n923), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI211_X1 g0730(.A(KEYINPUT39), .B(new_n915), .C1(new_n914), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n920), .A2(new_n358), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n901), .B(new_n900), .C1(new_n692), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n910), .A2(new_n912), .ZN(new_n935));
  INV_X1    g0735(.A(new_n906), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n937), .A3(KEYINPUT38), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n914), .B1(new_n903), .B2(new_n913), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT110), .B1(new_n931), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n930), .A2(new_n914), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(new_n932), .A3(new_n938), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT110), .ZN(new_n944));
  INV_X1    g0744(.A(new_n940), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n685), .A2(new_n439), .A3(new_n712), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n853), .A2(new_n856), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n704), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n772), .B2(new_n858), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n439), .A2(new_n704), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n462), .A2(new_n467), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n439), .B(new_n704), .C1(new_n685), .C2(new_n466), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n938), .A2(new_n939), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n959), .A2(new_n960), .B1(new_n933), .B2(new_n702), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n949), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n773), .A2(new_n469), .A3(new_n760), .A4(new_n766), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n695), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n915), .B1(new_n930), .B2(new_n914), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n754), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n731), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n957), .A2(new_n969), .A3(new_n862), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT40), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n861), .B1(new_n955), .B2(new_n956), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT40), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n960), .A4(new_n969), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n469), .A2(new_n969), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n978), .A2(new_n979), .A3(new_n710), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n898), .B1(new_n965), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n965), .B2(new_n981), .ZN(new_n983));
  INV_X1    g0783(.A(new_n606), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT35), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(KEYINPUT35), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n985), .A2(G116), .A3(new_n219), .A4(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n216), .A2(new_n228), .A3(new_n332), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n201), .A2(new_n222), .ZN(new_n992));
  OAI211_X1 g0792(.A(G1), .B(new_n265), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT106), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n983), .A2(new_n995), .ZN(G367));
  OAI21_X1  g0796(.A(new_n663), .B1(new_n610), .B2(new_n712), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(new_n761), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n704), .B1(new_n998), .B2(new_n618), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n618), .A2(new_n712), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n720), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT42), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n999), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n654), .A2(new_n655), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n704), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n665), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n651), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT111), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT43), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n999), .B(new_n1019), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1022), .A2(new_n1023), .B1(new_n716), .B2(new_n1002), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1010), .A2(new_n1018), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n716), .A2(new_n1002), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n1010), .C2(new_n1021), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n723), .B(KEYINPUT41), .Z(new_n1028));
  NAND3_X1  g0828(.A1(new_n720), .A2(new_n717), .A3(new_n1001), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT45), .Z(new_n1030));
  AOI21_X1  g0830(.A(new_n1001), .B1(new_n720), .B2(new_n717), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT44), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT113), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n716), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1030), .B(new_n1032), .C1(KEYINPUT113), .C2(new_n716), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n720), .B1(new_n715), .B2(new_n719), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(new_n711), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n774), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1028), .B1(new_n1040), .B2(new_n774), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1024), .B(new_n1027), .C1(new_n1041), .C2(new_n778), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n811), .A2(G77), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n331), .B2(new_n802), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n407), .B(new_n1044), .C1(G137), .C2(new_n813), .ZN(new_n1045));
  INV_X1    g0845(.A(G143), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n807), .C1(new_n258), .C2(new_n819), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n832), .A2(new_n222), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n201), .B2(new_n823), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n881), .B2(new_n829), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT114), .B1(new_n802), .B2(new_n547), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n844), .A2(G311), .B1(KEYINPUT46), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(KEYINPUT46), .B2(new_n1051), .C1(new_n566), .C2(new_n819), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n817), .A2(new_n206), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n336), .B1(new_n810), .B2(new_n205), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G317), .C2(new_n813), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n877), .B2(new_n880), .C1(new_n815), .C2(new_n829), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1047), .A2(new_n1050), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n796), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n779), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n791), .A2(new_n242), .B1(new_n722), .B2(new_n631), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n1062), .B2(new_n797), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n786), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1060), .B(new_n1063), .C1(new_n1064), .C2(new_n1014), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1042), .A2(new_n1065), .ZN(G387));
  AOI21_X1  g0866(.A(new_n724), .B1(new_n774), .B2(new_n1039), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n774), .B2(new_n1039), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n713), .A2(new_n714), .A3(new_n786), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n239), .A2(G45), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n291), .A2(new_n213), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1070), .A2(new_n792), .B1(new_n725), .B2(new_n1071), .ZN(new_n1072));
  OR3_X1    g0872(.A1(new_n257), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT50), .B1(new_n257), .B2(G50), .ZN(new_n1074));
  AOI21_X1  g0874(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1073), .A2(new_n725), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1072), .A2(new_n1076), .B1(new_n206), .B2(new_n722), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n779), .B1(new_n1077), .B2(new_n798), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n831), .A2(new_n631), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n880), .B2(new_n222), .C1(new_n257), .C2(new_n829), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n807), .A2(new_n881), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n819), .A2(new_n268), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n336), .B1(new_n811), .B2(G97), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n871), .A2(G77), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1083), .B(new_n1084), .C1(new_n258), .C2(new_n812), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT115), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n363), .B1(new_n811), .B2(G116), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n817), .A2(new_n877), .B1(new_n802), .B2(new_n815), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n820), .B1(new_n844), .B2(G322), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1090), .B1(new_n880), .B2(new_n566), .C1(new_n873), .C2(new_n829), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT48), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n1092), .B2(new_n1091), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT49), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1088), .B1(new_n808), .B2(new_n812), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1087), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1078), .B1(new_n1098), .B2(new_n796), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1039), .A2(new_n778), .B1(new_n1069), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1068), .A2(new_n1100), .ZN(G393));
  NAND2_X1  g0901(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1030), .A2(new_n716), .A3(new_n1032), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n774), .A2(new_n1039), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1040), .B(new_n723), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1001), .A2(new_n1064), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT116), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n840), .B1(G322), .B2(new_n813), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n877), .B2(new_n802), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n291), .B(new_n1110), .C1(G116), .C2(new_n885), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n815), .B2(new_n880), .C1(new_n566), .C2(new_n829), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G311), .A2(new_n820), .B1(new_n844), .B2(G317), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT52), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n258), .A2(new_n807), .B1(new_n819), .B2(new_n881), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT51), .Z(new_n1116));
  OAI22_X1  g0916(.A1(new_n1046), .A2(new_n812), .B1(new_n802), .B2(new_n222), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n336), .B(new_n1117), .C1(G87), .C2(new_n811), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n201), .A2(new_n824), .B1(new_n823), .B2(new_n400), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n831), .A2(G77), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1112), .A2(new_n1114), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n796), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n797), .B1(new_n205), .B2(new_n213), .C1(new_n792), .C2(new_n249), .ZN(new_n1124));
  AND4_X1   g0924(.A1(new_n779), .A2(new_n1108), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1104), .B2(new_n778), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT117), .B1(new_n1106), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1106), .A2(KEYINPUT117), .A3(new_n1126), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(G390));
  AOI21_X1  g0930(.A(new_n710), .B1(new_n731), .B2(new_n968), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n862), .A3(new_n957), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n756), .A2(new_n862), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n958), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT118), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n972), .A2(new_n1136), .A3(new_n1131), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n757), .A2(new_n857), .B1(new_n704), .B2(new_n951), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n712), .B1(new_n762), .B2(new_n765), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(new_n857), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(new_n952), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n756), .A2(new_n862), .A3(new_n957), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1131), .A2(new_n862), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1144), .C1(new_n957), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1140), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n469), .A2(new_n1131), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n963), .A2(new_n695), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n948), .B1(new_n1139), .B2(new_n957), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(KEYINPUT110), .B(new_n940), .C1(new_n966), .C2(new_n932), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n957), .B1(new_n1142), .B2(new_n952), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n966), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n947), .A3(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1156), .A2(new_n1159), .A3(new_n1144), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n972), .A2(new_n1136), .A3(new_n1131), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1136), .B1(new_n972), .B2(new_n1131), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1151), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1163), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1152), .B1(new_n941), .B2(new_n946), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1159), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1156), .A2(new_n1159), .A3(new_n1144), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1149), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n723), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n724), .B1(new_n1176), .B2(new_n1151), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(KEYINPUT119), .A3(new_n1172), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1169), .A2(new_n778), .A3(new_n1170), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n785), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n779), .B1(new_n868), .B2(new_n400), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1120), .B1(new_n880), .B2(new_n205), .C1(new_n206), .C2(new_n829), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G116), .A2(new_n820), .B1(new_n844), .B2(G283), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n841), .B(new_n888), .C1(G294), .C2(new_n813), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n407), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n871), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT53), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n802), .B2(new_n258), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n820), .A2(G132), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n844), .A2(G128), .ZN(new_n1192));
  INV_X1    g0992(.A(G125), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n262), .A2(new_n810), .B1(new_n1193), .B2(new_n812), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n407), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1191), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g0996(.A(KEYINPUT54), .B(G143), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n823), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n824), .A2(G137), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n832), .C2(new_n881), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1184), .A2(new_n1187), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1183), .B1(new_n1201), .B2(new_n796), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1182), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1180), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1179), .A2(new_n1205), .ZN(G378));
  NAND2_X1  g1006(.A1(new_n975), .A2(G330), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n271), .A2(new_n901), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n694), .A2(new_n310), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n312), .A2(new_n271), .A3(new_n901), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1207), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1214), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n975), .A2(G330), .A3(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1215), .A2(new_n949), .A3(new_n961), .A4(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n710), .B(new_n1214), .C1(new_n971), .C2(new_n974), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n975), .B2(G330), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n962), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n778), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n868), .A2(new_n201), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n363), .A2(G41), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G50), .B(new_n1225), .C1(new_n287), .C2(new_n275), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT120), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G97), .A2(new_n824), .B1(new_n823), .B2(new_n631), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT121), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n811), .A2(G58), .B1(new_n813), .B2(G283), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1084), .A3(new_n1225), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n819), .A2(new_n206), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n807), .A2(new_n547), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1048), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1229), .A2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT122), .Z(new_n1236));
  AOI21_X1  g1036(.A(new_n1227), .B1(new_n1236), .B2(KEYINPUT58), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n820), .A2(G128), .B1(new_n871), .B2(new_n1197), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT123), .Z(new_n1239));
  AOI22_X1  g1039(.A1(G132), .A2(new_n824), .B1(new_n823), .B2(G137), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n1193), .B2(new_n807), .C1(new_n258), .C2(new_n832), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT59), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(KEYINPUT124), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n287), .B(new_n275), .C1(new_n810), .C2(new_n881), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G124), .B2(new_n813), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT124), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1247), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1237), .B1(KEYINPUT58), .B2(new_n1236), .C1(new_n1245), .C2(new_n1249), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1061), .B(new_n1224), .C1(new_n1250), .C2(new_n796), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n785), .B2(new_n1216), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1223), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1172), .A2(new_n1150), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n723), .B1(new_n1255), .B2(KEYINPUT57), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1172), .A2(new_n1150), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1222), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1254), .B1(new_n1256), .B2(new_n1258), .ZN(G375));
  INV_X1    g1059(.A(new_n1028), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n957), .B1(new_n756), .B2(new_n862), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1161), .A2(new_n1162), .A3(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1149), .B(new_n1146), .C1(new_n1262), .C2(new_n953), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1151), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n958), .A2(new_n784), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n779), .B1(new_n868), .B2(G68), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1043), .B1(new_n566), .B2(new_n812), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n291), .B(new_n1267), .C1(G97), .C2(new_n871), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1268), .B1(new_n877), .B2(new_n819), .C1(new_n815), .C2(new_n807), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1079), .B1(new_n880), .B2(new_n206), .C1(new_n547), .C2(new_n829), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n844), .A2(G132), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n820), .A2(G137), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n336), .B1(new_n811), .B2(G58), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(G128), .A2(new_n813), .B1(new_n871), .B2(G159), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(G150), .A2(new_n823), .B1(new_n824), .B2(new_n1197), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n268), .B2(new_n832), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1269), .A2(new_n1270), .B1(new_n1275), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1266), .B1(new_n1278), .B2(new_n796), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1147), .A2(new_n778), .B1(new_n1265), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1264), .A2(new_n1280), .ZN(G381));
  NAND4_X1  g1081(.A1(new_n1128), .A2(new_n1042), .A3(new_n1065), .A4(new_n1129), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n896), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1282), .A2(G381), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1257), .A2(new_n1222), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT57), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n724), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1255), .A2(KEYINPUT57), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1253), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1204), .B1(new_n1177), .B2(new_n1172), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1290), .A3(new_n1291), .ZN(G407));
  NOR2_X1   g1092(.A1(new_n1285), .A2(new_n703), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1294));
  OAI21_X1  g1094(.A(G213), .B1(new_n1293), .B2(new_n1294), .ZN(G409));
  NOR2_X1   g1095(.A1(new_n1286), .A2(new_n1028), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1291), .B1(new_n1296), .B2(new_n1253), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1204), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(G375), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G213), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(G343), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1263), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1149), .A4(new_n1146), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1151), .A3(new_n723), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1280), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT125), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(KEYINPUT125), .A3(new_n1280), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(new_n896), .A3(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1307), .A2(new_n1308), .A3(G384), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1299), .A2(new_n1302), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT62), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT61), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1299), .A2(new_n1317), .A3(new_n1302), .A4(new_n1313), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1301), .A2(G2897), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1311), .A2(new_n1312), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1173), .A2(new_n1205), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1254), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1290), .B2(G378), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1322), .B1(new_n1326), .B2(new_n1301), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1315), .A2(new_n1316), .A3(new_n1318), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G390), .A2(G387), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n850), .B1(new_n1068), .B2(new_n1100), .ZN(new_n1330));
  OAI21_X1  g1130(.A(KEYINPUT127), .B1(new_n1283), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1329), .A2(new_n1282), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1283), .A2(new_n1330), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1333), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1333), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1329), .A2(new_n1282), .A3(new_n1331), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1328), .A2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT126), .B1(new_n1326), .B2(new_n1301), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT126), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1299), .A2(new_n1341), .A3(new_n1302), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1340), .A2(new_n1342), .A3(new_n1322), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT63), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1314), .A2(new_n1344), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1302), .A4(new_n1313), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1335), .A2(new_n1316), .A3(new_n1337), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1343), .A2(new_n1345), .A3(new_n1346), .A4(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1348), .ZN(G405));
  NAND2_X1  g1149(.A1(new_n1290), .A2(G378), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1291), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1352), .A2(new_n1312), .A3(new_n1311), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1350), .A2(new_n1313), .A3(new_n1351), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1338), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1355), .B(new_n1356), .ZN(G402));
endmodule


