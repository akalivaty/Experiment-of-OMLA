

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826;

  BUF_X1 U374 ( .A(n762), .Z(n792) );
  XOR2_X1 U375 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n400) );
  NOR2_X1 U376 ( .A1(n744), .A2(G902), .ZN(n541) );
  XNOR2_X1 U377 ( .A(G113), .B(G122), .ZN(n545) );
  XNOR2_X1 U378 ( .A(G140), .B(G137), .ZN(n517) );
  INV_X1 U379 ( .A(KEYINPUT8), .ZN(n480) );
  NAND2_X2 U380 ( .A1(n486), .A2(n484), .ZN(n357) );
  AND2_X1 U381 ( .A1(n732), .A2(n731), .ZN(n734) );
  NOR2_X4 U382 ( .A1(n394), .A2(n478), .ZN(n476) );
  AND2_X2 U383 ( .A1(n419), .A2(n488), .ZN(n374) );
  AND2_X2 U384 ( .A1(n497), .A2(n496), .ZN(n495) );
  NAND2_X1 U385 ( .A1(n656), .A2(n670), .ZN(n456) );
  XNOR2_X2 U386 ( .A(n652), .B(KEYINPUT0), .ZN(n670) );
  XNOR2_X2 U387 ( .A(n565), .B(n505), .ZN(n812) );
  XNOR2_X2 U388 ( .A(n574), .B(n504), .ZN(n565) );
  XNOR2_X2 U389 ( .A(G101), .B(KEYINPUT68), .ZN(n506) );
  XNOR2_X2 U390 ( .A(n506), .B(KEYINPUT67), .ZN(n539) );
  NAND2_X2 U391 ( .A1(n645), .A2(n633), .ZN(n533) );
  NAND2_X1 U392 ( .A1(n588), .A2(n395), .ZN(n589) );
  NAND2_X1 U393 ( .A1(n454), .A2(n453), .ZN(n441) );
  XNOR2_X2 U394 ( .A(G143), .B(G128), .ZN(n574) );
  NAND2_X1 U395 ( .A1(n353), .A2(n407), .ZN(n406) );
  NAND2_X1 U396 ( .A1(n409), .A2(n410), .ZN(n353) );
  XNOR2_X1 U397 ( .A(G143), .B(G128), .ZN(n423) );
  XNOR2_X1 U398 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n537) );
  XNOR2_X1 U399 ( .A(KEYINPUT100), .B(KEYINPUT101), .ZN(n552) );
  INV_X1 U400 ( .A(KEYINPUT15), .ZN(n520) );
  XOR2_X1 U401 ( .A(G116), .B(G137), .Z(n538) );
  INV_X1 U402 ( .A(G134), .ZN(n504) );
  INV_X1 U403 ( .A(G902), .ZN(n512) );
  XOR2_X1 U404 ( .A(G116), .B(G107), .Z(n566) );
  OR2_X1 U405 ( .A1(G237), .A2(G902), .ZN(n583) );
  XNOR2_X1 U406 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n354) );
  AND2_X2 U407 ( .A1(n389), .A2(n482), .ZN(n388) );
  NOR2_X2 U408 ( .A1(n782), .A2(n772), .ZN(n675) );
  XNOR2_X2 U409 ( .A(n671), .B(KEYINPUT31), .ZN(n782) );
  XNOR2_X2 U410 ( .A(n458), .B(KEYINPUT69), .ZN(n645) );
  INV_X1 U411 ( .A(n781), .ZN(n636) );
  NOR2_X2 U412 ( .A1(G953), .A2(G237), .ZN(n547) );
  XNOR2_X1 U413 ( .A(n746), .B(n367), .ZN(n366) );
  AND2_X1 U414 ( .A1(n387), .A2(KEYINPUT82), .ZN(n386) );
  OR2_X1 U415 ( .A1(n592), .A2(KEYINPUT81), .ZN(n485) );
  NAND2_X1 U416 ( .A1(n636), .A2(n770), .ZN(n704) );
  NAND2_X1 U417 ( .A1(n661), .A2(n692), .ZN(n458) );
  XNOR2_X1 U418 ( .A(n812), .B(G146), .ZN(n430) );
  INV_X1 U419 ( .A(n796), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n380), .B(n480), .ZN(n562) );
  INV_X1 U421 ( .A(G953), .ZN(n359) );
  INV_X1 U422 ( .A(KEYINPUT56), .ZN(n363) );
  NAND2_X1 U423 ( .A1(n366), .A2(n355), .ZN(n750) );
  AND2_X1 U424 ( .A1(n360), .A2(n359), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n723), .B(KEYINPUT119), .ZN(n360) );
  AND2_X1 U426 ( .A1(n361), .A2(n720), .ZN(n722) );
  INV_X1 U427 ( .A(n815), .ZN(n733) );
  NAND2_X1 U428 ( .A1(n500), .A2(n499), .ZN(n498) );
  NAND2_X1 U429 ( .A1(n494), .A2(n492), .ZN(n491) );
  OR2_X1 U430 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U431 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U432 ( .A1(n448), .A2(n446), .ZN(n625) );
  AND2_X1 U433 ( .A1(n450), .A2(n449), .ZN(n448) );
  INV_X2 U434 ( .A(n593), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n372), .B(KEYINPUT107), .ZN(n824) );
  NOR2_X1 U436 ( .A1(n682), .A2(n681), .ZN(n768) );
  NAND2_X1 U437 ( .A1(n374), .A2(n373), .ZN(n372) );
  NOR2_X1 U438 ( .A1(n634), .A2(n669), .ZN(n784) );
  NAND2_X1 U439 ( .A1(n375), .A2(n490), .ZN(n373) );
  AND2_X1 U440 ( .A1(n415), .A2(n398), .ZN(n411) );
  NOR2_X1 U441 ( .A1(n599), .A2(n598), .ZN(n466) );
  NOR2_X1 U442 ( .A1(n460), .A2(KEYINPUT106), .ZN(n490) );
  XNOR2_X1 U443 ( .A(n630), .B(n614), .ZN(n709) );
  BUF_X1 U444 ( .A(n690), .Z(n460) );
  INV_X1 U445 ( .A(n766), .ZN(n369) );
  XNOR2_X1 U446 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U447 ( .A1(n468), .A2(n467), .ZN(n394) );
  INV_X1 U448 ( .A(n745), .ZN(n367) );
  XNOR2_X1 U449 ( .A(n532), .B(KEYINPUT21), .ZN(n594) );
  NOR2_X1 U450 ( .A1(n647), .A2(n816), .ZN(n472) );
  NAND2_X1 U451 ( .A1(n562), .A2(G221), .ZN(n376) );
  XNOR2_X1 U452 ( .A(n578), .B(KEYINPUT16), .ZN(n580) );
  XNOR2_X1 U453 ( .A(n465), .B(G119), .ZN(n578) );
  XNOR2_X1 U454 ( .A(G113), .B(KEYINPUT3), .ZN(n465) );
  INV_X1 U455 ( .A(G210), .ZN(n584) );
  NAND2_X2 U456 ( .A1(G234), .A2(G237), .ZN(n534) );
  XNOR2_X1 U457 ( .A(G143), .B(G131), .ZN(n555) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(G131), .ZN(n505) );
  XNOR2_X2 U459 ( .A(KEYINPUT97), .B(KEYINPUT20), .ZN(n522) );
  NAND2_X1 U460 ( .A1(n357), .A2(n607), .ZN(n389) );
  INV_X1 U461 ( .A(n357), .ZN(n385) );
  XNOR2_X1 U462 ( .A(n791), .B(n790), .ZN(n362) );
  NAND2_X1 U463 ( .A1(n740), .A2(n688), .ZN(n361) );
  NOR2_X1 U464 ( .A1(n362), .A2(n796), .ZN(G54) );
  XNOR2_X1 U465 ( .A(n364), .B(n363), .ZN(G51) );
  NAND2_X1 U466 ( .A1(n368), .A2(n355), .ZN(n364) );
  XNOR2_X1 U467 ( .A(n365), .B(n354), .ZN(G60) );
  NAND2_X1 U468 ( .A1(n370), .A2(n355), .ZN(n365) );
  XNOR2_X1 U469 ( .A(n767), .B(n369), .ZN(n368) );
  XNOR2_X1 U470 ( .A(n761), .B(n371), .ZN(n370) );
  INV_X1 U471 ( .A(n760), .ZN(n371) );
  NOR2_X1 U472 ( .A1(n824), .A2(n823), .ZN(n664) );
  INV_X1 U473 ( .A(n660), .ZN(n375) );
  NAND2_X1 U474 ( .A1(n473), .A2(n393), .ZN(n815) );
  XNOR2_X1 U475 ( .A(n377), .B(n376), .ZN(n519) );
  XNOR2_X1 U476 ( .A(n379), .B(n378), .ZN(n377) );
  XNOR2_X1 U477 ( .A(n382), .B(KEYINPUT94), .ZN(n378) );
  XNOR2_X1 U478 ( .A(n381), .B(n383), .ZN(n379) );
  NAND2_X1 U479 ( .A1(n816), .A2(G234), .ZN(n380) );
  XNOR2_X2 U480 ( .A(G110), .B(KEYINPUT93), .ZN(n381) );
  XNOR2_X2 U481 ( .A(G128), .B(KEYINPUT23), .ZN(n382) );
  XNOR2_X2 U482 ( .A(G119), .B(KEYINPUT24), .ZN(n383) );
  NAND2_X1 U483 ( .A1(n388), .A2(n384), .ZN(n611) );
  NAND2_X1 U484 ( .A1(n356), .A2(n483), .ZN(n387) );
  BUF_X1 U485 ( .A(n732), .Z(n390) );
  AND2_X1 U486 ( .A1(n606), .A2(n485), .ZN(n484) );
  INV_X1 U487 ( .A(KEYINPUT79), .ZN(n478) );
  INV_X1 U488 ( .A(n649), .ZN(n467) );
  INV_X1 U489 ( .A(G900), .ZN(n469) );
  INV_X1 U490 ( .A(G224), .ZN(n502) );
  XNOR2_X1 U491 ( .A(n540), .B(n537), .ZN(n429) );
  NAND2_X1 U492 ( .A1(n770), .A2(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U493 ( .A(n463), .B(n462), .ZN(n628) );
  INV_X1 U494 ( .A(KEYINPUT110), .ZN(n462) );
  INV_X1 U495 ( .A(n414), .ZN(n410) );
  NAND2_X1 U496 ( .A1(n411), .A2(n416), .ZN(n409) );
  NAND2_X1 U497 ( .A1(n414), .A2(n412), .ZN(n407) );
  INV_X2 U498 ( .A(G953), .ZN(n816) );
  INV_X1 U499 ( .A(KEYINPUT81), .ZN(n483) );
  INV_X1 U500 ( .A(KEYINPUT109), .ZN(n471) );
  INV_X1 U501 ( .A(KEYINPUT76), .ZN(n612) );
  INV_X1 U502 ( .A(KEYINPUT44), .ZN(n493) );
  NOR2_X1 U503 ( .A1(n726), .A2(n815), .ZN(n730) );
  AND2_X1 U504 ( .A1(n544), .A2(n477), .ZN(n453) );
  INV_X1 U505 ( .A(G478), .ZN(n570) );
  AND2_X1 U506 ( .A1(n678), .A2(n392), .ZN(n499) );
  NOR2_X2 U507 ( .A1(n502), .A2(G953), .ZN(n501) );
  INV_X1 U508 ( .A(KEYINPUT108), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n430), .B(n426), .ZN(n744) );
  XNOR2_X1 U510 ( .A(n428), .B(n427), .ZN(n426) );
  XNOR2_X1 U511 ( .A(n578), .B(n538), .ZN(n427) );
  AND2_X1 U512 ( .A1(n489), .A2(n658), .ZN(n488) );
  INV_X1 U513 ( .A(KEYINPUT92), .ZN(n653) );
  INV_X1 U514 ( .A(G953), .ZN(n479) );
  XNOR2_X1 U515 ( .A(n569), .B(n568), .ZN(n793) );
  XNOR2_X1 U516 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U517 ( .A(n430), .B(n511), .ZN(n789) );
  XNOR2_X1 U518 ( .A(n749), .B(n748), .ZN(n796) );
  NAND2_X1 U519 ( .A1(n447), .A2(n391), .ZN(n446) );
  XNOR2_X1 U520 ( .A(n464), .B(n631), .ZN(n634) );
  NOR2_X1 U521 ( .A1(n638), .A2(n641), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n413), .A2(KEYINPUT35), .ZN(n405) );
  INV_X1 U523 ( .A(KEYINPUT111), .ZN(n459) );
  AND2_X1 U524 ( .A1(n617), .A2(n618), .ZN(n391) );
  AND2_X1 U525 ( .A1(n683), .A2(n677), .ZN(n392) );
  AND2_X1 U526 ( .A1(n751), .A2(n643), .ZN(n393) );
  AND2_X1 U527 ( .A1(n654), .A2(n630), .ZN(n395) );
  XOR2_X1 U528 ( .A(KEYINPUT6), .B(n667), .Z(n659) );
  AND2_X1 U529 ( .A1(n415), .A2(n654), .ZN(n396) );
  INV_X1 U530 ( .A(n770), .ZN(n617) );
  AND2_X1 U531 ( .A1(n476), .A2(n481), .ZN(n397) );
  AND2_X1 U532 ( .A1(n654), .A2(n412), .ZN(n398) );
  XNOR2_X1 U533 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n399) );
  OR2_X1 U534 ( .A1(n721), .A2(n431), .ZN(n401) );
  AND2_X1 U535 ( .A1(n607), .A2(n483), .ZN(n402) );
  INV_X1 U536 ( .A(KEYINPUT35), .ZN(n412) );
  INV_X1 U537 ( .A(KEYINPUT78), .ZN(n481) );
  XOR2_X1 U538 ( .A(n684), .B(KEYINPUT45), .Z(n403) );
  AND2_X1 U539 ( .A1(n725), .A2(n731), .ZN(n404) );
  NAND2_X1 U540 ( .A1(n406), .A2(n405), .ZN(n823) );
  NAND2_X1 U541 ( .A1(n417), .A2(n418), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n396), .A2(n416), .ZN(n413) );
  AND2_X1 U543 ( .A1(n674), .A2(KEYINPUT34), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n431), .A2(KEYINPUT34), .ZN(n415) );
  NOR2_X1 U545 ( .A1(n431), .A2(KEYINPUT34), .ZN(n417) );
  INV_X1 U546 ( .A(n674), .ZN(n418) );
  NAND2_X1 U547 ( .A1(n660), .A2(KEYINPUT106), .ZN(n419) );
  XNOR2_X2 U548 ( .A(n456), .B(n400), .ZN(n660) );
  INV_X1 U549 ( .A(n657), .ZN(n420) );
  NAND2_X1 U550 ( .A1(n437), .A2(n436), .ZN(n421) );
  NAND2_X1 U551 ( .A1(n437), .A2(n436), .ZN(n435) );
  XNOR2_X1 U552 ( .A(n472), .B(n471), .ZN(n470) );
  NAND2_X1 U553 ( .A1(n470), .A2(n469), .ZN(n468) );
  XNOR2_X2 U554 ( .A(n605), .B(n604), .ZN(n778) );
  OR2_X2 U555 ( .A1(n778), .A2(n608), .ZN(n606) );
  XNOR2_X1 U556 ( .A(n539), .B(n429), .ZN(n428) );
  BUF_X1 U557 ( .A(n812), .Z(n422) );
  NAND2_X1 U558 ( .A1(n439), .A2(n421), .ZN(n424) );
  NAND2_X1 U559 ( .A1(n439), .A2(n435), .ZN(n588) );
  BUF_X1 U560 ( .A(n600), .Z(n630) );
  INV_X1 U561 ( .A(n659), .ZN(n443) );
  XNOR2_X1 U562 ( .A(n425), .B(n445), .ZN(n444) );
  NAND2_X1 U563 ( .A1(n646), .A2(n690), .ZN(n425) );
  XNOR2_X1 U564 ( .A(n602), .B(n601), .ZN(n651) );
  NOR2_X1 U565 ( .A1(n660), .A2(n443), .ZN(n679) );
  XNOR2_X1 U566 ( .A(n432), .B(n577), .ZN(n581) );
  NOR2_X1 U567 ( .A1(n714), .A2(n431), .ZN(n715) );
  XNOR2_X2 U568 ( .A(n442), .B(n399), .ZN(n431) );
  XNOR2_X1 U569 ( .A(n433), .B(n576), .ZN(n432) );
  XNOR2_X1 U570 ( .A(n434), .B(n423), .ZN(n433) );
  XNOR2_X1 U571 ( .A(n503), .B(n501), .ZN(n434) );
  INV_X1 U572 ( .A(n441), .ZN(n436) );
  AND2_X2 U573 ( .A1(n438), .A2(KEYINPUT78), .ZN(n437) );
  NAND2_X1 U574 ( .A1(n452), .A2(n476), .ZN(n438) );
  AND2_X2 U575 ( .A1(n440), .A2(n451), .ZN(n439) );
  NAND2_X1 U576 ( .A1(n441), .A2(n481), .ZN(n440) );
  NAND2_X1 U577 ( .A1(n444), .A2(n443), .ZN(n442) );
  INV_X1 U578 ( .A(n637), .ZN(n447) );
  NAND2_X1 U579 ( .A1(n637), .A2(KEYINPUT40), .ZN(n450) );
  NAND2_X1 U580 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U581 ( .A1(n452), .A2(n397), .ZN(n451) );
  INV_X1 U582 ( .A(n672), .ZN(n452) );
  NAND2_X1 U583 ( .A1(n672), .A2(n478), .ZN(n454) );
  XNOR2_X1 U584 ( .A(n626), .B(KEYINPUT46), .ZN(n457) );
  NOR2_X1 U585 ( .A1(n457), .A2(n461), .ZN(n475) );
  XNOR2_X2 U586 ( .A(KEYINPUT32), .B(n663), .ZN(n825) );
  XNOR2_X1 U587 ( .A(n633), .B(n632), .ZN(n690) );
  XNOR2_X2 U588 ( .A(n616), .B(n615), .ZN(n637) );
  BUF_X2 U589 ( .A(n645), .Z(n646) );
  XNOR2_X2 U590 ( .A(n498), .B(n403), .ZN(n732) );
  XNOR2_X1 U591 ( .A(n455), .B(n635), .ZN(n473) );
  NAND2_X1 U592 ( .A1(n474), .A2(n475), .ZN(n455) );
  OR2_X2 U593 ( .A1(n531), .A2(n525), .ZN(n527) );
  NAND2_X1 U594 ( .A1(n593), .A2(n487), .ZN(n486) );
  XNOR2_X2 U595 ( .A(n589), .B(n459), .ZN(n593) );
  XNOR2_X1 U596 ( .A(n784), .B(KEYINPUT86), .ZN(n461) );
  NOR2_X1 U597 ( .A1(n659), .A2(n627), .ZN(n463) );
  NAND2_X1 U598 ( .A1(n466), .A2(n603), .ZN(n605) );
  NAND2_X1 U599 ( .A1(n689), .A2(n466), .ZN(n623) );
  XNOR2_X1 U600 ( .A(n613), .B(n612), .ZN(n474) );
  INV_X1 U601 ( .A(n625), .ZN(n752) );
  XNOR2_X2 U602 ( .A(n533), .B(KEYINPUT98), .ZN(n672) );
  NAND2_X1 U603 ( .A1(n394), .A2(n478), .ZN(n477) );
  NAND2_X1 U604 ( .A1(n732), .A2(n404), .ZN(n726) );
  AND2_X1 U605 ( .A1(n390), .A2(n479), .ZN(n807) );
  XNOR2_X2 U606 ( .A(G146), .B(G125), .ZN(n575) );
  XNOR2_X2 U607 ( .A(G104), .B(G110), .ZN(n798) );
  XNOR2_X2 U608 ( .A(G902), .B(KEYINPUT89), .ZN(n521) );
  XNOR2_X2 U609 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X2 U610 ( .A(n529), .B(n528), .ZN(n661) );
  NAND2_X1 U611 ( .A1(n356), .A2(n402), .ZN(n482) );
  AND2_X1 U612 ( .A1(n592), .A2(KEYINPUT81), .ZN(n487) );
  NAND2_X1 U613 ( .A1(n460), .A2(KEYINPUT106), .ZN(n489) );
  NAND2_X1 U614 ( .A1(n495), .A2(n491), .ZN(n500) );
  AND2_X1 U615 ( .A1(n665), .A2(n493), .ZN(n492) );
  INV_X1 U616 ( .A(n666), .ZN(n494) );
  NAND2_X1 U617 ( .A1(KEYINPUT74), .A2(KEYINPUT44), .ZN(n496) );
  NAND2_X1 U618 ( .A1(n666), .A2(KEYINPUT74), .ZN(n497) );
  XNOR2_X2 U619 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n503) );
  NAND2_X1 U620 ( .A1(n600), .A2(n708), .ZN(n602) );
  INV_X1 U621 ( .A(n826), .ZN(n624) );
  INV_X1 U622 ( .A(KEYINPUT74), .ZN(n665) );
  INV_X1 U623 ( .A(n594), .ZN(n692) );
  AND2_X1 U624 ( .A1(n655), .A2(n692), .ZN(n656) );
  INV_X1 U625 ( .A(KEYINPUT19), .ZN(n601) );
  INV_X1 U626 ( .A(KEYINPUT48), .ZN(n635) );
  XNOR2_X1 U627 ( .A(n571), .B(n570), .ZN(n572) );
  BUF_X1 U628 ( .A(n763), .Z(n765) );
  XNOR2_X1 U629 ( .A(n573), .B(n572), .ZN(n619) );
  XNOR2_X1 U630 ( .A(n670), .B(n653), .ZN(n674) );
  XNOR2_X1 U631 ( .A(n798), .B(KEYINPUT72), .ZN(n507) );
  XNOR2_X1 U632 ( .A(n539), .B(n507), .ZN(n577) );
  NAND2_X1 U633 ( .A1(n816), .A2(G227), .ZN(n508) );
  XNOR2_X1 U634 ( .A(n508), .B(G107), .ZN(n509) );
  XNOR2_X1 U635 ( .A(n509), .B(n517), .ZN(n510) );
  XNOR2_X1 U636 ( .A(n577), .B(n510), .ZN(n511) );
  NAND2_X1 U637 ( .A1(n789), .A2(n512), .ZN(n516) );
  XNOR2_X1 U638 ( .A(KEYINPUT71), .B(G469), .ZN(n514) );
  INV_X1 U639 ( .A(KEYINPUT70), .ZN(n513) );
  XNOR2_X1 U640 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X2 U641 ( .A(n516), .B(n515), .ZN(n633) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT10), .ZN(n551) );
  INV_X1 U643 ( .A(n517), .ZN(n518) );
  XNOR2_X1 U644 ( .A(n551), .B(n518), .ZN(n813) );
  XNOR2_X1 U645 ( .A(n519), .B(n813), .ZN(n754) );
  OR2_X2 U646 ( .A1(n754), .A2(G902), .ZN(n529) );
  XNOR2_X1 U647 ( .A(n521), .B(n520), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n582), .A2(G234), .ZN(n524) );
  XNOR2_X1 U649 ( .A(n522), .B(KEYINPUT96), .ZN(n523) );
  XNOR2_X1 U650 ( .A(n524), .B(n523), .ZN(n531) );
  INV_X1 U651 ( .A(G217), .ZN(n525) );
  XNOR2_X1 U652 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n526) );
  INV_X1 U653 ( .A(G221), .ZN(n530) );
  OR2_X1 U654 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U655 ( .A(n534), .B(KEYINPUT14), .ZN(n536) );
  NAND2_X1 U656 ( .A1(n536), .A2(G902), .ZN(n535) );
  XOR2_X1 U657 ( .A(KEYINPUT91), .B(n535), .Z(n647) );
  NAND2_X1 U658 ( .A1(G952), .A2(n536), .ZN(n719) );
  NOR2_X1 U659 ( .A1(n719), .A2(G953), .ZN(n649) );
  NAND2_X1 U660 ( .A1(G210), .A2(n547), .ZN(n540) );
  XNOR2_X2 U661 ( .A(n541), .B(G472), .ZN(n667) );
  NAND2_X1 U662 ( .A1(G214), .A2(n583), .ZN(n708) );
  INV_X1 U663 ( .A(n708), .ZN(n542) );
  NOR2_X1 U664 ( .A1(n667), .A2(n542), .ZN(n543) );
  XNOR2_X1 U665 ( .A(n543), .B(KEYINPUT30), .ZN(n544) );
  XOR2_X1 U666 ( .A(G104), .B(G140), .Z(n546) );
  XNOR2_X1 U667 ( .A(n546), .B(n545), .ZN(n549) );
  NAND2_X1 U668 ( .A1(G214), .A2(n547), .ZN(n548) );
  XNOR2_X1 U669 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U670 ( .A(n551), .B(n550), .Z(n558) );
  XOR2_X2 U671 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n553) );
  XNOR2_X1 U672 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U673 ( .A(n554), .B(KEYINPUT12), .Z(n556) );
  XNOR2_X1 U674 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U675 ( .A(n558), .B(n557), .ZN(n759) );
  NOR2_X1 U676 ( .A1(G902), .A2(n759), .ZN(n560) );
  XNOR2_X1 U677 ( .A(KEYINPUT103), .B(KEYINPUT13), .ZN(n559) );
  XNOR2_X1 U678 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U679 ( .A(n561), .B(G475), .ZN(n620) );
  XOR2_X1 U680 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n564) );
  NAND2_X1 U681 ( .A1(n562), .A2(G217), .ZN(n563) );
  XNOR2_X1 U682 ( .A(n564), .B(n563), .ZN(n569) );
  INV_X1 U683 ( .A(n565), .ZN(n567) );
  XNOR2_X1 U684 ( .A(G122), .B(n566), .ZN(n579) );
  XNOR2_X1 U685 ( .A(n567), .B(n579), .ZN(n568) );
  NOR2_X1 U686 ( .A1(G902), .A2(n793), .ZN(n573) );
  INV_X1 U687 ( .A(KEYINPUT104), .ZN(n571) );
  NOR2_X1 U688 ( .A1(n620), .A2(n619), .ZN(n654) );
  XNOR2_X1 U689 ( .A(n575), .B(KEYINPUT4), .ZN(n576) );
  XNOR2_X1 U690 ( .A(n580), .B(n579), .ZN(n799) );
  XNOR2_X1 U691 ( .A(n581), .B(n799), .ZN(n763) );
  INV_X1 U692 ( .A(n582), .ZN(n731) );
  INV_X1 U693 ( .A(n731), .ZN(n728) );
  NAND2_X1 U694 ( .A1(n763), .A2(n728), .ZN(n587) );
  INV_X1 U695 ( .A(n583), .ZN(n585) );
  NOR2_X1 U696 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X2 U697 ( .A(n587), .B(n586), .ZN(n600) );
  INV_X1 U698 ( .A(n619), .ZN(n590) );
  AND2_X1 U699 ( .A1(n620), .A2(n590), .ZN(n781) );
  OR2_X1 U700 ( .A1(n590), .A2(n620), .ZN(n770) );
  INV_X1 U701 ( .A(KEYINPUT47), .ZN(n608) );
  NOR2_X1 U702 ( .A1(n704), .A2(n608), .ZN(n591) );
  INV_X1 U703 ( .A(n591), .ZN(n592) );
  NOR2_X1 U704 ( .A1(n394), .A2(n594), .ZN(n595) );
  INV_X1 U705 ( .A(n661), .ZN(n657) );
  NAND2_X1 U706 ( .A1(n595), .A2(n657), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n667), .A2(n627), .ZN(n596) );
  XOR2_X1 U708 ( .A(KEYINPUT28), .B(n596), .Z(n599) );
  INV_X1 U709 ( .A(KEYINPUT112), .ZN(n597) );
  XNOR2_X1 U710 ( .A(n633), .B(n597), .ZN(n598) );
  INV_X1 U711 ( .A(n651), .ZN(n603) );
  INV_X1 U712 ( .A(KEYINPUT80), .ZN(n604) );
  INV_X1 U713 ( .A(KEYINPUT82), .ZN(n607) );
  AND2_X1 U714 ( .A1(n704), .A2(n608), .ZN(n609) );
  NAND2_X1 U715 ( .A1(n778), .A2(n609), .ZN(n610) );
  NAND2_X1 U716 ( .A1(n611), .A2(n610), .ZN(n613) );
  INV_X1 U717 ( .A(KEYINPUT38), .ZN(n614) );
  NAND2_X1 U718 ( .A1(n424), .A2(n709), .ZN(n616) );
  INV_X1 U719 ( .A(KEYINPUT39), .ZN(n615) );
  INV_X1 U720 ( .A(KEYINPUT40), .ZN(n618) );
  NAND2_X1 U721 ( .A1(n620), .A2(n619), .ZN(n711) );
  NAND2_X1 U722 ( .A1(n709), .A2(n708), .ZN(n705) );
  NOR2_X1 U723 ( .A1(n711), .A2(n705), .ZN(n621) );
  XOR2_X1 U724 ( .A(KEYINPUT41), .B(n621), .Z(n689) );
  XNOR2_X1 U725 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n622) );
  XNOR2_X1 U726 ( .A(n623), .B(n622), .ZN(n826) );
  XOR2_X1 U727 ( .A(KEYINPUT36), .B(KEYINPUT114), .Z(n631) );
  NOR2_X1 U728 ( .A1(n770), .A2(n628), .ZN(n629) );
  NAND2_X1 U729 ( .A1(n629), .A2(n708), .ZN(n638) );
  INV_X1 U730 ( .A(n630), .ZN(n641) );
  XNOR2_X1 U731 ( .A(KEYINPUT1), .B(KEYINPUT66), .ZN(n632) );
  INV_X1 U732 ( .A(n460), .ZN(n669) );
  OR2_X1 U733 ( .A1(n637), .A2(n636), .ZN(n751) );
  NOR2_X1 U734 ( .A1(n638), .A2(n460), .ZN(n640) );
  INV_X1 U735 ( .A(KEYINPUT43), .ZN(n639) );
  XNOR2_X1 U736 ( .A(n640), .B(n639), .ZN(n642) );
  AND2_X1 U737 ( .A1(n642), .A2(n641), .ZN(n786) );
  INV_X1 U738 ( .A(n786), .ZN(n643) );
  NAND2_X1 U739 ( .A1(n733), .A2(KEYINPUT2), .ZN(n644) );
  XNOR2_X1 U740 ( .A(n644), .B(KEYINPUT85), .ZN(n685) );
  XOR2_X1 U741 ( .A(G898), .B(KEYINPUT90), .Z(n806) );
  NAND2_X1 U742 ( .A1(G953), .A2(n806), .ZN(n802) );
  NOR2_X1 U743 ( .A1(n647), .A2(n802), .ZN(n648) );
  NOR2_X1 U744 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X2 U745 ( .A1(n651), .A2(n650), .ZN(n652) );
  INV_X1 U746 ( .A(n711), .ZN(n655) );
  AND2_X1 U747 ( .A1(n667), .A2(n657), .ZN(n658) );
  XNOR2_X1 U748 ( .A(n420), .B(KEYINPUT105), .ZN(n680) );
  INV_X1 U749 ( .A(n680), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n669), .A2(n693), .ZN(n662) );
  NAND2_X1 U751 ( .A1(n679), .A2(n662), .ZN(n663) );
  NAND2_X1 U752 ( .A1(n664), .A2(n825), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n666), .A2(KEYINPUT44), .ZN(n678) );
  INV_X1 U754 ( .A(n667), .ZN(n699) );
  NAND2_X1 U755 ( .A1(n699), .A2(n646), .ZN(n668) );
  NOR2_X1 U756 ( .A1(n669), .A2(n668), .ZN(n701) );
  NAND2_X1 U757 ( .A1(n670), .A2(n701), .ZN(n671) );
  OR2_X1 U758 ( .A1(n699), .A2(n672), .ZN(n673) );
  NOR2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n772) );
  XNOR2_X1 U760 ( .A(n675), .B(KEYINPUT99), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n676), .A2(n704), .ZN(n677) );
  XNOR2_X1 U762 ( .A(KEYINPUT87), .B(n679), .ZN(n682) );
  OR2_X1 U763 ( .A1(n460), .A2(n680), .ZN(n681) );
  INV_X1 U764 ( .A(n768), .ZN(n683) );
  INV_X1 U765 ( .A(KEYINPUT84), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n685), .A2(n390), .ZN(n740) );
  AND2_X1 U767 ( .A1(n733), .A2(n390), .ZN(n686) );
  INV_X1 U768 ( .A(n686), .ZN(n687) );
  INV_X1 U769 ( .A(KEYINPUT2), .ZN(n727) );
  NAND2_X1 U770 ( .A1(n687), .A2(n727), .ZN(n688) );
  INV_X1 U771 ( .A(n689), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n460), .A2(n646), .ZN(n691) );
  XOR2_X1 U773 ( .A(KEYINPUT50), .B(n691), .Z(n697) );
  NOR2_X1 U774 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U775 ( .A(KEYINPUT117), .B(n694), .Z(n695) );
  XNOR2_X1 U776 ( .A(KEYINPUT49), .B(n695), .ZN(n696) );
  NAND2_X1 U777 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U778 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U779 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U780 ( .A(KEYINPUT51), .B(n702), .Z(n703) );
  NOR2_X1 U781 ( .A1(n721), .A2(n703), .ZN(n716) );
  INV_X1 U782 ( .A(n704), .ZN(n706) );
  NOR2_X1 U783 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U784 ( .A(KEYINPUT118), .B(n707), .ZN(n713) );
  NOR2_X1 U785 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U786 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U788 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U789 ( .A(n717), .B(KEYINPUT52), .ZN(n718) );
  NAND2_X1 U790 ( .A1(n722), .A2(n401), .ZN(n723) );
  XNOR2_X1 U791 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n724) );
  XNOR2_X1 U792 ( .A(n358), .B(n724), .ZN(G75) );
  INV_X1 U793 ( .A(KEYINPUT83), .ZN(n725) );
  NOR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n730), .A2(n729), .ZN(n737) );
  NAND2_X1 U796 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U797 ( .A1(n735), .A2(KEYINPUT83), .ZN(n736) );
  NAND2_X1 U798 ( .A1(n737), .A2(n736), .ZN(n739) );
  INV_X1 U799 ( .A(KEYINPUT65), .ZN(n738) );
  XNOR2_X1 U800 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U801 ( .A1(n741), .A2(n740), .ZN(n743) );
  INV_X1 U802 ( .A(KEYINPUT64), .ZN(n742) );
  XNOR2_X2 U803 ( .A(n743), .B(n742), .ZN(n762) );
  NAND2_X1 U804 ( .A1(n762), .A2(G472), .ZN(n746) );
  XNOR2_X1 U805 ( .A(n744), .B(KEYINPUT62), .ZN(n745) );
  INV_X1 U806 ( .A(G952), .ZN(n747) );
  NAND2_X1 U807 ( .A1(n747), .A2(G953), .ZN(n749) );
  INV_X1 U808 ( .A(KEYINPUT88), .ZN(n748) );
  XNOR2_X1 U809 ( .A(n750), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U810 ( .A(n751), .B(G134), .ZN(G36) );
  XOR2_X1 U811 ( .A(G131), .B(n752), .Z(G33) );
  XNOR2_X1 U812 ( .A(G143), .B(KEYINPUT116), .ZN(n753) );
  XOR2_X1 U813 ( .A(n753), .B(n356), .Z(G45) );
  NAND2_X1 U814 ( .A1(n792), .A2(G217), .ZN(n756) );
  BUF_X1 U815 ( .A(n754), .Z(n755) );
  XNOR2_X1 U816 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U817 ( .A1(n757), .A2(n796), .ZN(G66) );
  NAND2_X1 U818 ( .A1(n762), .A2(G475), .ZN(n761) );
  XOR2_X1 U819 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n758) );
  NAND2_X1 U820 ( .A1(n762), .A2(G210), .ZN(n767) );
  XNOR2_X1 U821 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n764) );
  XNOR2_X1 U822 ( .A(G101), .B(n768), .ZN(n769) );
  XNOR2_X1 U823 ( .A(n769), .B(KEYINPUT115), .ZN(G3) );
  NAND2_X1 U824 ( .A1(n617), .A2(n772), .ZN(n771) );
  XNOR2_X1 U825 ( .A(G104), .B(n771), .ZN(G6) );
  XOR2_X1 U826 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n774) );
  NAND2_X1 U827 ( .A1(n772), .A2(n781), .ZN(n773) );
  XNOR2_X1 U828 ( .A(n774), .B(n773), .ZN(n775) );
  XNOR2_X1 U829 ( .A(G107), .B(n775), .ZN(G9) );
  XOR2_X1 U830 ( .A(G128), .B(KEYINPUT29), .Z(n777) );
  NAND2_X1 U831 ( .A1(n781), .A2(n778), .ZN(n776) );
  XNOR2_X1 U832 ( .A(n777), .B(n776), .ZN(G30) );
  NAND2_X1 U833 ( .A1(n778), .A2(n617), .ZN(n779) );
  XNOR2_X1 U834 ( .A(n779), .B(G146), .ZN(G48) );
  NAND2_X1 U835 ( .A1(n782), .A2(n617), .ZN(n780) );
  XNOR2_X1 U836 ( .A(n780), .B(G113), .ZN(G15) );
  NAND2_X1 U837 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U838 ( .A(n783), .B(G116), .ZN(G18) );
  XNOR2_X1 U839 ( .A(G125), .B(n784), .ZN(n785) );
  XNOR2_X1 U840 ( .A(n785), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U841 ( .A(G140), .B(n786), .Z(G42) );
  NAND2_X1 U842 ( .A1(n792), .A2(G469), .ZN(n791) );
  XOR2_X1 U843 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n787) );
  XNOR2_X1 U844 ( .A(n787), .B(KEYINPUT121), .ZN(n788) );
  XNOR2_X1 U845 ( .A(n789), .B(n788), .ZN(n790) );
  NAND2_X1 U846 ( .A1(n792), .A2(G478), .ZN(n795) );
  XNOR2_X1 U847 ( .A(n793), .B(KEYINPUT124), .ZN(n794) );
  XNOR2_X1 U848 ( .A(n795), .B(n794), .ZN(n797) );
  NOR2_X1 U849 ( .A1(n797), .A2(n796), .ZN(G63) );
  XNOR2_X1 U850 ( .A(G101), .B(n798), .ZN(n800) );
  XNOR2_X1 U851 ( .A(n800), .B(n799), .ZN(n801) );
  NAND2_X1 U852 ( .A1(n802), .A2(n801), .ZN(n810) );
  NAND2_X1 U853 ( .A1(G224), .A2(G953), .ZN(n803) );
  XNOR2_X1 U854 ( .A(n803), .B(KEYINPUT61), .ZN(n804) );
  XNOR2_X1 U855 ( .A(n804), .B(KEYINPUT125), .ZN(n805) );
  NOR2_X1 U856 ( .A1(n806), .A2(n805), .ZN(n808) );
  NOR2_X1 U857 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U858 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U859 ( .A(KEYINPUT126), .B(n811), .ZN(G69) );
  XNOR2_X1 U860 ( .A(n422), .B(KEYINPUT127), .ZN(n814) );
  XNOR2_X1 U861 ( .A(n814), .B(n813), .ZN(n818) );
  XNOR2_X1 U862 ( .A(n815), .B(n818), .ZN(n817) );
  NAND2_X1 U863 ( .A1(n817), .A2(n816), .ZN(n822) );
  XNOR2_X1 U864 ( .A(G227), .B(n818), .ZN(n819) );
  NAND2_X1 U865 ( .A1(n819), .A2(G900), .ZN(n820) );
  NAND2_X1 U866 ( .A1(n820), .A2(G953), .ZN(n821) );
  NAND2_X1 U867 ( .A1(n822), .A2(n821), .ZN(G72) );
  XOR2_X1 U868 ( .A(n823), .B(G122), .Z(G24) );
  XOR2_X1 U869 ( .A(n824), .B(G110), .Z(G12) );
  XNOR2_X1 U870 ( .A(G119), .B(n825), .ZN(G21) );
  XOR2_X1 U871 ( .A(G137), .B(n826), .Z(G39) );
endmodule

