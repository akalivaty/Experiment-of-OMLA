//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT99), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G78gat), .ZN(new_n204));
  INV_X1    g003(.A(G64gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G57gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n203), .B(new_n204), .C1(KEYINPUT99), .C2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT100), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n202), .A2(new_n210), .ZN(new_n211));
  OAI22_X1  g010(.A1(new_n207), .A2(new_n209), .B1(new_n204), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(G127gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n213), .B2(new_n212), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n217), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(G183gat), .B(G211gat), .Z(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n231), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT41), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT15), .ZN(new_n238));
  XNOR2_X1  g037(.A(G43gat), .B(G50gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT94), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n240), .B2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT14), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(G29gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G36gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT14), .B(G29gat), .Z(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(G36gat), .ZN(new_n247));
  OR3_X1    g046(.A1(new_n242), .A2(new_n247), .A3(KEYINPUT95), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT95), .B1(new_n242), .B2(new_n247), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n239), .A2(KEYINPUT15), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n248), .A2(new_n249), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G85gat), .A2(G92gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT7), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT103), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT8), .ZN(new_n256));
  AND2_X1   g055(.A1(G99gat), .A2(G106gat), .ZN(new_n257));
  OAI221_X1 g056(.A(new_n255), .B1(G85gat), .B2(G92gat), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(new_n253), .B2(KEYINPUT103), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(KEYINPUT103), .B2(new_n253), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(G99gat), .A2(G106gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n257), .A2(new_n262), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n258), .B2(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n252), .A2(KEYINPUT17), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT96), .B(KEYINPUT17), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n252), .B2(new_n268), .ZN(new_n269));
  OAI221_X1 g068(.A(new_n237), .B1(new_n252), .B2(new_n266), .C1(new_n267), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G190gat), .B(G218gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT104), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT105), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n236), .A2(KEYINPUT41), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT101), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT102), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n273), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n272), .A2(KEYINPUT105), .ZN(new_n282));
  XNOR2_X1  g081(.A(G134gat), .B(G162gat), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n278), .A2(new_n284), .A3(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n235), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G120gat), .B(G148gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G176gat), .B(G204gat), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n261), .A2(KEYINPUT106), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n212), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n266), .ZN(new_n297));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n263), .B(new_n265), .C1(new_n212), .C2(new_n295), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n294), .B1(new_n302), .B2(KEYINPUT107), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(KEYINPUT107), .B2(new_n302), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT10), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n266), .A2(new_n305), .A3(new_n212), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n297), .A2(new_n300), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n305), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n299), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n294), .B1(new_n309), .B2(new_n302), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT34), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  INV_X1    g119(.A(G127gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G134gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G113gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(G120gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(G120gat), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G120gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(G113gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n324), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT72), .B1(new_n326), .B2(new_n331), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(G113gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n328), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n323), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n321), .A2(KEYINPUT71), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G127gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n319), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n339), .A2(KEYINPUT73), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT73), .B1(new_n339), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n334), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  INV_X1    g153(.A(G176gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(KEYINPUT23), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT65), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(KEYINPUT67), .A3(new_n363), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT24), .ZN(new_n368));
  INV_X1    g167(.A(G183gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G183gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT25), .B1(new_n374), .B2(KEYINPUT23), .ZN(new_n375));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT24), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n373), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n366), .A2(new_n367), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT64), .B(G169gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n374), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n382), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n359), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n377), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n370), .A2(new_n372), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n368), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n380), .B1(new_n387), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n379), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n356), .A2(new_n393), .A3(new_n357), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n356), .A2(KEYINPUT69), .A3(new_n393), .A4(new_n357), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n385), .A2(KEYINPUT26), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n359), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n369), .A2(KEYINPUT27), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G183gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n400), .A2(new_n402), .A3(new_n371), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT27), .B(G183gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT28), .A3(new_n371), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT68), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT68), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n399), .A2(new_n408), .A3(new_n410), .A4(new_n376), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n338), .A2(new_n323), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n337), .B1(new_n336), .B2(new_n328), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n347), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n339), .A2(KEYINPUT73), .A3(new_n347), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(KEYINPUT75), .A3(new_n334), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n352), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n408), .A2(new_n410), .A3(new_n376), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n422), .A2(new_n399), .B1(new_n379), .B2(new_n391), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n351), .A3(new_n350), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G227gat), .ZN(new_n426));
  INV_X1    g225(.A(G233gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n318), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(KEYINPUT34), .B(new_n428), .C1(new_n421), .C2(new_n424), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n428), .A3(new_n424), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT32), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G71gat), .B(G99gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(KEYINPUT76), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT33), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(KEYINPUT32), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n432), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n432), .B1(new_n445), .B2(new_n441), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n317), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n441), .A2(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(new_n432), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n441), .A3(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(KEYINPUT91), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G211gat), .A2(G218gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT22), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(KEYINPUT78), .A3(new_n460), .ZN(new_n464));
  XNOR2_X1  g263(.A(G197gat), .B(G204gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G211gat), .ZN(new_n467));
  INV_X1    g266(.A(G218gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n466), .A2(new_n459), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT79), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n459), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n463), .A2(new_n473), .A3(new_n465), .A4(new_n464), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n470), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G226gat), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n427), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT80), .B1(new_n423), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT80), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n412), .A2(new_n482), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n423), .B2(KEYINPUT29), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n477), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n412), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n423), .A2(new_n480), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n488), .A2(new_n489), .A3(new_n476), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n458), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n485), .B(new_n477), .C1(new_n480), .C2(new_n423), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n481), .B2(new_n483), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n457), .C1(new_n493), .C2(new_n477), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(KEYINPUT30), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n486), .A2(new_n490), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n457), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT88), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n333), .B1(new_n417), .B2(new_n418), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506));
  AND2_X1   g305(.A1(G155gat), .A2(G162gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(G155gat), .A2(G162gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(G155gat), .A2(G162gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT81), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT2), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G141gat), .B(G148gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n509), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT82), .B1(new_n507), .B2(new_n512), .ZN(new_n516));
  AND2_X1   g315(.A1(G141gat), .A2(G148gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(G141gat), .A2(G148gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G155gat), .B(G162gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT82), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n510), .A2(new_n521), .A3(KEYINPUT2), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n516), .A2(new_n519), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT3), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT3), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n515), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n504), .B1(new_n505), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n527), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n515), .B2(new_n523), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n350), .A2(KEYINPUT83), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G225gat), .A2(G233gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n524), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n419), .A2(new_n334), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT4), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n333), .B(new_n524), .C1(new_n417), .C2(new_n418), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT4), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n534), .A2(new_n535), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(KEYINPUT84), .A2(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n535), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n536), .B1(new_n419), .B2(new_n334), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(new_n540), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT85), .B(new_n545), .C1(new_n546), .C2(new_n540), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(KEYINPUT5), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n537), .B(KEYINPUT4), .ZN(new_n552));
  INV_X1    g351(.A(new_n543), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n535), .A3(new_n534), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n544), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G1gat), .B(G29gat), .Z(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G85gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT6), .ZN(new_n562));
  INV_X1    g361(.A(new_n560), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n544), .A2(new_n551), .A3(new_n554), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AND4_X1   g364(.A1(new_n563), .A2(new_n544), .A3(new_n551), .A4(new_n554), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT87), .B1(new_n566), .B2(KEYINPUT6), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n564), .A2(new_n568), .A3(new_n562), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n565), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G50gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n527), .A2(new_n487), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n476), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G228gat), .A2(G233gat), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT29), .B1(new_n470), .B2(new_n474), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n524), .B1(new_n577), .B2(KEYINPUT3), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n472), .A2(new_n487), .A3(new_n475), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n536), .B1(new_n580), .B2(new_n526), .ZN(new_n581));
  OAI211_X1 g380(.A(G228gat), .B(G233gat), .C1(new_n581), .C2(new_n574), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n572), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G78gat), .B(G106gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G22gat), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n582), .A3(new_n572), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n583), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n454), .A2(new_n503), .A3(new_n570), .A4(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n591), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n597), .A2(new_n446), .A3(new_n447), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n598), .A3(new_n499), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n595), .A2(new_n596), .B1(new_n599), .B2(KEYINPUT35), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n566), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n568), .B1(new_n564), .B2(new_n562), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n593), .B1(new_n603), .B2(new_n565), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(KEYINPUT92), .A3(new_n503), .A4(new_n454), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n535), .B1(new_n552), .B2(new_n534), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n563), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n350), .A2(new_n524), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n535), .A3(new_n537), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT89), .ZN(new_n611));
  INV_X1    g410(.A(new_n534), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n541), .A2(new_n539), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n545), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n614), .A3(KEYINPUT39), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT40), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n616), .A2(new_n566), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(new_n615), .A3(KEYINPUT40), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n501), .A2(new_n502), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n597), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n621));
  AOI21_X1  g420(.A(new_n457), .B1(new_n496), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n622), .B1(new_n623), .B2(new_n496), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT38), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n493), .A2(new_n476), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n488), .A2(new_n489), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n623), .B1(new_n627), .B2(new_n476), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT38), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n622), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n494), .A3(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n619), .B(new_n620), .C1(new_n631), .C2(new_n570), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n446), .A2(new_n447), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT77), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n451), .A2(new_n452), .B1(new_n635), .B2(KEYINPUT36), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n570), .A2(new_n499), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n638), .B2(new_n597), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n600), .A2(new_n605), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n223), .B1(new_n252), .B2(new_n268), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n267), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G229gat), .A2(G233gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n252), .A2(new_n223), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(KEYINPUT18), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n643), .B(KEYINPUT13), .Z(new_n647));
  AND2_X1   g446(.A1(new_n252), .A2(new_n223), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n644), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n645), .B(new_n643), .C1(new_n267), .C2(new_n641), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G197gat), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT11), .B(G169gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT93), .B(KEYINPUT12), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT97), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n646), .A2(new_n652), .A3(new_n659), .A4(new_n649), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n653), .A2(KEYINPUT97), .A3(new_n660), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n316), .B1(new_n640), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n451), .A2(KEYINPUT91), .A3(new_n452), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT91), .B1(new_n451), .B2(new_n452), .ZN(new_n669));
  INV_X1    g468(.A(new_n502), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT88), .B1(new_n495), .B2(new_n498), .ZN(new_n671));
  OAI22_X1  g470(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n570), .A2(new_n594), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n596), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n599), .A2(KEYINPUT35), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n605), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n639), .A2(new_n632), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n666), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(KEYINPUT98), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n315), .B1(new_n667), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n570), .B(KEYINPUT108), .Z(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g483(.A(KEYINPUT109), .B(KEYINPUT16), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n222), .ZN(new_n686));
  AND4_X1   g485(.A1(new_n502), .A2(new_n681), .A3(new_n501), .A4(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n503), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n222), .B1(new_n681), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n687), .ZN(G1325gat));
  INV_X1    g490(.A(new_n681), .ZN(new_n692));
  INV_X1    g491(.A(new_n637), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n454), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n692), .B2(new_n696), .ZN(G1326gat));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n597), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n667), .A2(new_n680), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n234), .A2(new_n313), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n288), .ZN(new_n704));
  INV_X1    g503(.A(new_n682), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(G29gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n701), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n704), .A4(new_n706), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n640), .B2(new_n288), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n289), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n703), .A2(new_n666), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n712), .A2(new_n682), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G29gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n709), .A2(new_n710), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT110), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n709), .A2(new_n710), .A3(new_n719), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1328gat));
  AND2_X1   g520(.A1(new_n712), .A2(new_n713), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n688), .A3(new_n714), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G36gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n503), .A2(G36gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n701), .A2(new_n704), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n726), .A2(new_n727), .A3(KEYINPUT46), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(KEYINPUT46), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n724), .B1(KEYINPUT46), .B2(new_n726), .C1(new_n728), .C2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n637), .A3(new_n713), .A4(new_n714), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n695), .A2(G43gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n701), .A2(new_n704), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n731), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1330gat));
  NAND4_X1  g537(.A1(new_n712), .A2(new_n597), .A3(new_n713), .A4(new_n714), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n620), .A2(G50gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n701), .A2(new_n704), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g543(.A1(new_n290), .A2(new_n666), .A3(new_n313), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n640), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n682), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT113), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  XNOR2_X1  g548(.A(new_n503), .B(KEYINPUT114), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT49), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n205), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT115), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n746), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n205), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1333gat));
  INV_X1    g555(.A(new_n746), .ZN(new_n757));
  OAI21_X1  g556(.A(G71gat), .B1(new_n757), .B2(new_n693), .ZN(new_n758));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n746), .A2(new_n759), .A3(new_n454), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n597), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(G78gat), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n679), .A2(new_n234), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n314), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n722), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n705), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n288), .B1(new_n676), .B2(new_n677), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n766), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n314), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G85gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n682), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n778), .ZN(G1336gat));
  INV_X1    g578(.A(new_n750), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n769), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(G92gat), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n722), .A2(new_n688), .A3(new_n768), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n786), .A2(G92gat), .B1(new_n776), .B2(new_n782), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n769), .B2(new_n693), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n695), .A2(G99gat), .A3(new_n314), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT117), .Z(new_n791));
  AND4_X1   g590(.A1(KEYINPUT51), .A2(new_n678), .A3(new_n289), .A4(new_n766), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT51), .B1(new_n771), .B2(new_n766), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n789), .A2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n620), .A2(G106gat), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n313), .B(new_n797), .C1(new_n792), .C2(new_n793), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n712), .A2(new_n597), .A3(new_n713), .A4(new_n768), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(KEYINPUT118), .B(G106gat), .Z(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n799), .A2(new_n800), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n796), .B(new_n798), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n799), .A2(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n798), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(KEYINPUT53), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT119), .B(new_n796), .C1(new_n808), .C2(new_n798), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n293), .B1(new_n309), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n308), .A2(new_n299), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n308), .B2(new_n299), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n310), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n814), .B(KEYINPUT55), .C1(new_n815), .C2(new_n816), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n664), .A2(new_n819), .A3(new_n665), .A4(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n648), .A2(new_n644), .A3(new_n647), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT121), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n643), .B1(new_n642), .B2(new_n645), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n657), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n825), .A2(new_n663), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n313), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n289), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n819), .A2(new_n820), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n663), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n829), .A2(new_n288), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n235), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n290), .A2(new_n666), .A3(new_n314), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n705), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n598), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n780), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n679), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n833), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n695), .A2(new_n597), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n780), .A2(new_n682), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n666), .A2(new_n325), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(G1340gat));
  AOI21_X1  g643(.A(G120gat), .B1(new_n836), .B2(new_n313), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n314), .A2(new_n330), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(G1341gat));
  NAND4_X1  g646(.A1(new_n836), .A2(new_n340), .A3(new_n342), .A4(new_n234), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n340), .A2(new_n342), .ZN(new_n849));
  INV_X1    g648(.A(new_n842), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n235), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(G1342gat));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n319), .A3(new_n503), .A4(new_n289), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n850), .B2(new_n288), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n637), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n620), .B1(new_n832), .B2(new_n833), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n862), .B(new_n620), .C1(new_n832), .C2(new_n833), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n679), .A2(G141gat), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(G141gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n637), .A2(new_n620), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n834), .A2(new_n780), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n867), .B1(new_n869), .B2(new_n666), .ZN(new_n870));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n866), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n866), .B2(new_n870), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1344gat));
  OAI211_X1 g673(.A(new_n313), .B(new_n859), .C1(new_n861), .C2(new_n863), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n876));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(KEYINPUT59), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n875), .B2(new_n878), .ZN(new_n880));
  INV_X1    g679(.A(new_n863), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n289), .A2(new_n826), .A3(new_n820), .A4(new_n819), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n821), .A2(new_n827), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n289), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT125), .B1(new_n828), .B2(new_n831), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n235), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n620), .B1(new_n887), .B2(new_n833), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n881), .B1(new_n888), .B2(KEYINPUT57), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n841), .A2(new_n637), .A3(new_n314), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n877), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n879), .A2(new_n880), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n869), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n877), .A3(new_n313), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n864), .B2(new_n235), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n227), .A3(new_n234), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n864), .B2(new_n288), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n834), .A2(new_n868), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n688), .A2(new_n288), .A3(G162gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G1347gat));
  AOI21_X1  g702(.A(new_n682), .B1(new_n832), .B2(new_n833), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n904), .A2(new_n598), .A3(new_n750), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n381), .A3(new_n679), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n682), .A2(new_n503), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n838), .A2(new_n839), .A3(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n679), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT127), .B(new_n906), .C1(new_n911), .C2(new_n354), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n354), .B1(new_n910), .B2(new_n679), .ZN(new_n914));
  INV_X1    g713(.A(new_n906), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n905), .A2(new_n355), .A3(new_n313), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n910), .A2(new_n313), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n355), .ZN(G1349gat));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n406), .A3(new_n234), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n910), .A2(new_n234), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n369), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n369), .B1(new_n910), .B2(new_n234), .ZN(new_n925));
  INV_X1    g724(.A(new_n922), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n371), .A3(new_n289), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n910), .A2(new_n289), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(G190gat), .ZN(new_n932));
  AOI211_X1 g731(.A(KEYINPUT61), .B(new_n371), .C1(new_n910), .C2(new_n289), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(G1351gat));
  AND3_X1   g733(.A1(new_n904), .A2(new_n750), .A3(new_n868), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n679), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n907), .A2(new_n693), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n889), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n679), .A2(G197gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(G1352gat));
  INV_X1    g740(.A(G204gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n942), .A3(new_n313), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT62), .Z(new_n944));
  AND2_X1   g743(.A1(new_n939), .A2(new_n313), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n945), .B2(new_n942), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n935), .A2(new_n467), .A3(new_n234), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n889), .A2(new_n234), .A3(new_n938), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n468), .A3(new_n289), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n939), .A2(new_n289), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n468), .ZN(G1355gat));
endmodule


