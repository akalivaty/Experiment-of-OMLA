//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n568, new_n570, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR3_X1   g026(.A1(G221), .A2(G219), .A3(G218), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n437), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT67), .B(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G125), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n459), .A2(G137), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n464), .A2(new_n465), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n468), .B1(new_n474), .B2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n459), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT70), .Z(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n459), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n480), .A2(new_n485), .ZN(G162));
  NAND3_X1  g061(.A1(new_n466), .A2(new_n459), .A3(G138), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n466), .A2(new_n459), .A3(G138), .A4(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n494), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n466), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI211_X1 g083(.A(G50), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n510), .A2(new_n511), .B1(new_n507), .B2(new_n508), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n503), .A2(new_n519), .A3(G88), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n506), .B1(new_n516), .B2(new_n521), .ZN(G166));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n517), .B2(new_n518), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n511), .A2(new_n510), .ZN(new_n529));
  OAI21_X1  g104(.A(G89), .B1(new_n507), .B2(new_n508), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(G168));
  NAND3_X1  g108(.A1(new_n503), .A2(new_n519), .A3(G90), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n519), .A2(G52), .A3(G543), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(G64), .B1(new_n511), .B2(new_n510), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n505), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n519), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n512), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n543), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n524), .B(G53), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n529), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n501), .A2(new_n502), .B1(new_n517), .B2(new_n518), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n563), .A2(G651), .B1(new_n564), .B2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  AND2_X1   g142(.A1(new_n530), .A2(new_n531), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n525), .B(new_n527), .C1(new_n568), .C2(new_n529), .ZN(G286));
  INV_X1    g144(.A(new_n521), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT72), .B1(new_n520), .B2(new_n509), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(new_n505), .B2(new_n504), .ZN(G303));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n501), .A2(new_n573), .A3(new_n502), .ZN(new_n574));
  AOI22_X1  g149(.A1(G49), .A2(new_n524), .B1(new_n574), .B2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n564), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT75), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n529), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n564), .A2(G86), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  INV_X1    g160(.A(G48), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n543), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n524), .A2(KEYINPUT76), .A3(G48), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n503), .A2(G60), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n505), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n564), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND3_X1  g171(.A1(new_n564), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n512), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n529), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G299), .A2(new_n607), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n466), .A2(new_n469), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT77), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT78), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n478), .A2(G123), .B1(G135), .B2(new_n481), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n459), .C2(G111), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n628), .B1(new_n627), .B2(new_n629), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n626), .B(new_n633), .C1(new_n624), .C2(new_n623), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n644), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n652), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  OAI221_X1 g234(.A(new_n654), .B1(new_n653), .B2(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n654), .A2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT81), .B(G2096), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(G2100), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n674), .B(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT82), .Z(new_n681));
  OAI211_X1 g256(.A(new_n678), .B(new_n679), .C1(new_n681), .C2(new_n673), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G2090), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT99), .Z(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G21), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G168), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT97), .B(G1966), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n632), .A2(G29), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G19), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n547), .B2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(G1341), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n704), .B(new_n708), .C1(G1341), .C2(new_n707), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n481), .A2(G141), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n711), .A3(G105), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n494), .A2(G105), .A3(G2104), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(KEYINPUT95), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n494), .A2(KEYINPUT67), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2105), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n720), .A2(new_n466), .A3(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT26), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT96), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(G141), .A2(new_n481), .B1(new_n712), .B2(new_n714), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n728), .A2(new_n729), .A3(new_n721), .A4(new_n724), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(new_n693), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n693), .B2(G32), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n699), .A2(G4), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n614), .B2(new_n699), .ZN(new_n738));
  INV_X1    g313(.A(G1348), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n734), .A2(new_n735), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n709), .A2(new_n736), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G11), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT98), .B(G28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(new_n693), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n744), .A2(KEYINPUT30), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(G171), .A2(new_n699), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G5), .B2(new_n699), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(new_n701), .B2(new_n703), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n748), .B(new_n752), .C1(new_n751), .C2(new_n750), .ZN(new_n753));
  NOR2_X1   g328(.A1(G27), .A2(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G164), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n753), .B(new_n757), .C1(new_n696), .C2(G2090), .ZN(new_n758));
  AND2_X1   g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  NOR2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n693), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT94), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G160), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n693), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n481), .A2(G140), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n459), .A2(G116), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n478), .A2(KEYINPUT88), .A3(G128), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n720), .A2(new_n466), .A3(G128), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n771), .B1(new_n780), .B2(new_n693), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n765), .A2(new_n769), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n742), .A2(new_n758), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n693), .A2(G33), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT93), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n481), .A2(G139), .ZN(new_n788));
  AND2_X1   g363(.A1(G103), .A2(G2104), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n717), .A2(new_n719), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n717), .A2(new_n719), .A3(new_n789), .A4(KEYINPUT90), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n794));
  AND3_X1   g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n788), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n794), .ZN(new_n800));
  AOI21_X1  g375(.A(KEYINPUT90), .B1(new_n459), .B2(new_n789), .ZN(new_n801));
  INV_X1    g376(.A(new_n793), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n805), .A2(KEYINPUT91), .A3(new_n788), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G127), .ZN(new_n808));
  INV_X1    g383(.A(G115), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n472), .A2(new_n808), .B1(new_n809), .B2(new_n463), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI221_X1 g387(.A(KEYINPUT92), .B1(new_n809), .B2(new_n463), .C1(new_n472), .C2(new_n808), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n812), .A2(new_n720), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n787), .B1(new_n807), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g391(.A(KEYINPUT93), .B(new_n814), .C1(new_n799), .C2(new_n806), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n786), .B1(new_n818), .B2(new_n693), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n698), .B(new_n785), .C1(new_n819), .C2(G2072), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G2072), .B2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n481), .A2(G131), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT83), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT84), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n463), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .C1(G107), .C2(new_n459), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n478), .A2(G119), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT85), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n693), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(G25), .B2(new_n693), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT35), .B(G1991), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT86), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n832), .A2(new_n835), .ZN(new_n837));
  MUX2_X1   g412(.A(G24), .B(G290), .S(G16), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1986), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n699), .A2(G23), .ZN(new_n841));
  INV_X1    g416(.A(new_n577), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n699), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT33), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1976), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n699), .A2(G22), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G166), .B2(new_n699), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(G1971), .Z(new_n848));
  NOR2_X1   g423(.A1(G6), .A2(G16), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n587), .A2(new_n588), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n582), .A2(new_n583), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n849), .B1(new_n852), .B2(G16), .ZN(new_n853));
  XOR2_X1   g428(.A(KEYINPUT32), .B(G1981), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n845), .A2(new_n848), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(KEYINPUT34), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n840), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n859), .B(new_n860), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n821), .A2(new_n861), .ZN(G150));
  INV_X1    g437(.A(G150), .ZN(G311));
  NAND2_X1  g438(.A1(new_n614), .A2(G559), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT100), .B(G93), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n543), .A2(new_n866), .B1(new_n512), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n503), .A2(G67), .ZN(new_n869));
  NAND2_X1  g444(.A1(G80), .A2(G543), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n505), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n547), .A2(new_n872), .ZN(new_n873));
  OAI22_X1  g448(.A1(new_n542), .A2(new_n546), .B1(new_n868), .B2(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n865), .B(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n878));
  INV_X1    g453(.A(G860), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(KEYINPUT39), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n872), .A2(new_n879), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  OR3_X1    g459(.A1(new_n630), .A2(new_n631), .A3(G160), .ZN(new_n885));
  OAI21_X1  g460(.A(G160), .B1(new_n630), .B2(new_n631), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(G162), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(G162), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT103), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n887), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT101), .B1(new_n816), .B2(new_n817), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT91), .B1(new_n805), .B2(new_n788), .ZN(new_n896));
  INV_X1    g471(.A(new_n788), .ZN(new_n897));
  AOI211_X1 g472(.A(new_n798), .B(new_n897), .C1(new_n803), .C2(new_n804), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n815), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT93), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n807), .A2(new_n787), .A3(new_n815), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n780), .A2(new_n726), .A3(new_n730), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n776), .A2(new_n779), .ZN(new_n905));
  INV_X1    g480(.A(new_n775), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n726), .A2(new_n730), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n904), .A2(new_n907), .A3(new_n499), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n727), .B2(new_n731), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n780), .A2(new_n726), .A3(new_n730), .ZN(new_n911));
  AOI21_X1  g486(.A(G164), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n895), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n829), .B(new_n622), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n478), .A2(G130), .ZN(new_n916));
  OAI221_X1 g491(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n459), .C2(G118), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n481), .A2(G142), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n915), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n499), .B1(new_n904), .B2(new_n907), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(G164), .A3(new_n911), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n818), .A2(new_n902), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n914), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n914), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n894), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n894), .B(new_n930), .C1(new_n926), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n914), .A2(new_n925), .ZN(new_n933));
  INV_X1    g508(.A(new_n921), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n914), .A2(new_n921), .A3(new_n925), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n888), .A2(new_n889), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(KEYINPUT102), .A3(new_n936), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G37), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n932), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  NAND4_X1  g520(.A1(new_n560), .A2(new_n601), .A3(new_n565), .A4(new_n605), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n560), .A2(new_n565), .B1(new_n601), .B2(new_n605), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g525(.A1(G299), .A2(new_n606), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n946), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT105), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n875), .B(new_n617), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT41), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(new_n959), .A3(new_n946), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n957), .B1(new_n956), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(G290), .A2(new_n577), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n594), .A2(new_n595), .A3(new_n576), .A4(new_n575), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(G166), .A2(KEYINPUT107), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n506), .C1(new_n516), .C2(new_n521), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n852), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G303), .A2(new_n972), .ZN(new_n975));
  NAND2_X1  g550(.A1(G166), .A2(KEYINPUT107), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(G305), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n970), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n971), .A2(new_n973), .A3(new_n852), .ZN(new_n979));
  AOI21_X1  g554(.A(G305), .B1(new_n975), .B2(new_n976), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G47), .ZN(new_n982));
  INV_X1    g557(.A(G85), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n543), .A2(new_n982), .B1(new_n512), .B2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n577), .A2(new_n593), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n594), .A2(new_n595), .B1(new_n575), .B2(new_n576), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT108), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n968), .A2(new_n969), .A3(new_n967), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n978), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT42), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n966), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n965), .A2(KEYINPUT109), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n966), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(G868), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G868), .B2(new_n872), .ZN(G295));
  OAI21_X1  g571(.A(new_n995), .B1(G868), .B2(new_n872), .ZN(G331));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n536), .B2(new_n539), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n537), .A2(new_n538), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G651), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n1001), .A3(new_n535), .A4(new_n534), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1002), .A3(G286), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G168), .A2(G171), .A3(new_n1001), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n875), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1003), .A2(new_n873), .A3(new_n1004), .A4(new_n874), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n876), .A2(KEYINPUT111), .A3(new_n1004), .A4(new_n1003), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n949), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n987), .B1(new_n979), .B2(new_n980), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n989), .A2(new_n974), .A3(new_n977), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n961), .B2(new_n963), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1018), .A2(new_n943), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n958), .A2(new_n960), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1009), .A2(new_n1010), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n950), .A2(new_n954), .A3(new_n1008), .A4(new_n1006), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n990), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1019), .A2(KEYINPUT43), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT41), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n959), .B1(new_n951), .B2(new_n946), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1029), .A2(new_n962), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n952), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n990), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT43), .B1(new_n1019), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT43), .ZN(new_n1035));
  AND4_X1   g610(.A1(new_n1035), .A2(new_n1024), .A3(new_n1018), .A4(new_n943), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n943), .A3(new_n1018), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT43), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(KEYINPUT112), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1040), .A3(KEYINPUT43), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1034), .B1(new_n1042), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g618(.A1(G160), .A2(G40), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n499), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1049), .B(KEYINPUT113), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n909), .A2(G2067), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n780), .A2(new_n782), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1054), .B(KEYINPUT114), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT115), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1050), .A2(new_n732), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1049), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1059), .A2(G1996), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(G1996), .B2(new_n732), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n830), .A2(new_n835), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT125), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1057), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1050), .B1(new_n1065), .B2(new_n1053), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1060), .B(KEYINPUT46), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1058), .A3(new_n1056), .ZN(new_n1068));
  XOR2_X1   g643(.A(new_n1068), .B(KEYINPUT47), .Z(new_n1069));
  XNOR2_X1  g644(.A(new_n829), .B(new_n834), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1051), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(G290), .A2(G1986), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1049), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1073), .B(KEYINPUT48), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n1062), .A2(new_n1057), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1066), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  AND2_X1   g652(.A1(G160), .A2(G40), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1046), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT45), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1080), .A3(new_n756), .A4(new_n1048), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT53), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1078), .A2(new_n1083), .A3(KEYINPUT122), .A4(new_n1084), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n751), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(G301), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1077), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1082), .A2(new_n1089), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G171), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1090), .A3(KEYINPUT54), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  INV_X1    g672(.A(G8), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1078), .A2(new_n1080), .A3(new_n1048), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n702), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1084), .A2(G40), .A3(G160), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n764), .A3(new_n1083), .ZN(new_n1104));
  AOI21_X1  g679(.A(G286), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1104), .A3(G286), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1104), .A3(G168), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n1109), .B2(G8), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1976), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(G288), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1079), .A2(G40), .A3(G160), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n842), .A2(G1976), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1113), .A2(G8), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(G8), .A3(new_n1115), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT52), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n850), .A2(new_n851), .A3(G1981), .ZN(new_n1120));
  INV_X1    g695(.A(G1981), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n584), .B2(new_n589), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(G1981), .B1(new_n850), .B2(new_n851), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n584), .A2(new_n1121), .A3(new_n589), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(KEYINPUT49), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1123), .A2(G8), .A3(new_n1114), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1116), .A2(new_n1118), .A3(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1048), .A2(G40), .A3(G160), .ZN(new_n1129));
  AOI21_X1  g704(.A(G1971), .B1(new_n1129), .B2(new_n1080), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT116), .B(G2090), .Z(new_n1131));
  AND4_X1   g706(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .A4(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(G8), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G166), .A2(new_n1098), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT55), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1128), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(G8), .B(new_n1135), .C1(new_n1130), .C2(new_n1132), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1093), .A2(new_n1096), .A3(new_n1111), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1114), .A2(KEYINPUT121), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1079), .A2(G160), .A3(new_n1142), .A4(G40), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT58), .B(G1341), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1144), .A2(new_n1145), .B1(G1996), .B2(new_n1101), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n547), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1146), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g729(.A(G299), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT119), .B(G1956), .Z(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1103), .B2(new_n1083), .ZN(new_n1160));
  XNOR2_X1  g735(.A(KEYINPUT56), .B(G2072), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1078), .A2(new_n1080), .A3(new_n1048), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1158), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1129), .A2(new_n1080), .A3(new_n1161), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1085), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1164), .B(new_n1157), .C1(new_n1165), .C2(new_n1159), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1152), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1151), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1087), .A2(new_n739), .A3(new_n1088), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1144), .A2(new_n782), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT60), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1171), .A2(new_n1172), .A3(new_n1175), .A4(KEYINPUT60), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n614), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1174), .A2(new_n1180), .A3(new_n614), .A4(new_n1176), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1167), .A2(new_n1168), .A3(new_n1152), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1170), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n606), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1163), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1166), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1140), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(G288), .A2(G1976), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1120), .B1(new_n1127), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT117), .ZN(new_n1192));
  OAI211_X1 g767(.A(G8), .B(new_n1114), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n1193), .A2(new_n1194), .B1(new_n1138), .B2(new_n1128), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1098), .B(G286), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1128), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1138), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT63), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1137), .A2(KEYINPUT63), .A3(new_n1138), .A4(new_n1197), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1195), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT118), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1206), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1107), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1099), .B1(new_n1208), .B2(new_n1105), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1110), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT62), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1207), .A2(new_n1139), .A3(new_n1211), .A4(new_n1092), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1212), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1189), .A2(new_n1205), .A3(new_n1213), .ZN(new_n1214));
  AND2_X1   g789(.A1(G290), .A2(G1986), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1049), .B1(new_n1072), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g791(.A1(new_n1057), .A2(new_n1062), .A3(new_n1216), .A4(new_n1071), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1076), .B1(new_n1214), .B2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n666), .A2(new_n669), .A3(G319), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1221), .A2(KEYINPUT126), .ZN(new_n1222));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n1223));
  NAND4_X1  g797(.A1(new_n666), .A2(new_n669), .A3(new_n1223), .A4(G319), .ZN(new_n1224));
  AOI21_X1  g798(.A(G401), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n1225), .B1(new_n690), .B2(new_n691), .ZN(new_n1226));
  AOI21_X1  g800(.A(new_n1226), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1227));
  AND3_X1   g801(.A1(new_n944), .A2(new_n1220), .A3(new_n1227), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1220), .B1(new_n944), .B2(new_n1227), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1228), .A2(new_n1229), .ZN(G308));
  NAND2_X1  g804(.A1(new_n944), .A2(new_n1227), .ZN(new_n1231));
  NAND2_X1  g805(.A1(new_n1231), .A2(KEYINPUT127), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n944), .A2(new_n1227), .A3(new_n1220), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1233), .ZN(G225));
endmodule


