//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT93), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT93), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n202), .A2(new_n206), .A3(new_n203), .ZN(new_n207));
  AND2_X1   g006(.A1(G57gat), .A2(G64gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G57gat), .A2(G64gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT92), .B1(G71gat), .B2(G78gat), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n213), .B1(new_n211), .B2(new_n214), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(G127gat), .ZN(new_n220));
  XOR2_X1   g019(.A(G15gat), .B(G22gat), .Z(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G8gat), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n214), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n212), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n231), .B1(new_n235), .B2(KEYINPUT21), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n220), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  XNOR2_X1  g037(.A(G155gat), .B(G183gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n237), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G231gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(G211gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n241), .B(new_n244), .Z(new_n245));
  INV_X1    g044(.A(KEYINPUT97), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT14), .ZN(new_n247));
  INV_X1    g046(.A(G29gat), .ZN(new_n248));
  INV_X1    g047(.A(G36gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(KEYINPUT88), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT88), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G29gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n255), .A3(G36gat), .ZN(new_n256));
  INV_X1    g055(.A(G43gat), .ZN(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260));
  NAND2_X1  g059(.A1(G43gat), .A2(G50gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n252), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n261), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n252), .B2(new_n256), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT15), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n252), .A2(new_n256), .A3(new_n262), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT15), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT17), .ZN(new_n271));
  NAND2_X1  g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT7), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(G85gat), .A3(G92gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G99gat), .A2(G106gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G85gat), .ZN(new_n281));
  INV_X1    g080(.A(G92gat), .ZN(new_n282));
  AOI22_X1  g081(.A1(KEYINPUT8), .A2(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n276), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n280), .B1(new_n276), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT94), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n276), .A2(new_n283), .ZN(new_n287));
  INV_X1    g086(.A(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n276), .A2(new_n280), .A3(new_n283), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n270), .A2(new_n271), .A3(new_n286), .A4(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT88), .B(G29gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(G36gat), .B1(new_n250), .B2(new_n251), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT15), .B1(new_n295), .B2(new_n262), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n267), .B1(new_n295), .B2(new_n264), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(KEYINPUT15), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n286), .A2(new_n292), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(KEYINPUT17), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G190gat), .B(G218gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n303), .B(KEYINPUT95), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n293), .A2(new_n300), .A3(new_n304), .A4(new_n301), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT96), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n246), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT96), .B(KEYINPUT97), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n306), .A2(KEYINPUT96), .A3(new_n307), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G134gat), .ZN(new_n315));
  INV_X1    g114(.A(G162gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n318), .B1(new_n310), .B2(new_n311), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n245), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324));
  OR3_X1    g123(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n325), .A2(new_n326), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT25), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT24), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT66), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT64), .B(G190gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OR3_X1    g138(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(G169gat), .ZN(new_n342));
  INV_X1    g141(.A(G176gat), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n340), .B(new_n341), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n335), .A3(new_n334), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n330), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n333), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n338), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT65), .B1(new_n348), .B2(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT65), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n338), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n331), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n328), .B1(new_n353), .B2(new_n327), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n324), .B1(new_n355), .B2(KEYINPUT29), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n335), .B(KEYINPUT66), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT28), .B1(new_n357), .B2(new_n348), .ZN(new_n358));
  INV_X1    g157(.A(new_n346), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n332), .B2(new_n329), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n353), .A2(new_n327), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(G226gat), .A3(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT22), .ZN(new_n366));
  XOR2_X1   g165(.A(KEYINPUT72), .B(G211gat), .Z(new_n367));
  INV_X1    g166(.A(G218gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n374), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n365), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n378), .A3(new_n364), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(KEYINPUT85), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n356), .A2(new_n383), .A3(new_n364), .A4(new_n378), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(KEYINPUT37), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT86), .ZN(new_n386));
  XOR2_X1   g185(.A(G8gat), .B(G36gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G64gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(new_n282), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n380), .A2(new_n381), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT37), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n382), .A2(new_n395), .A3(KEYINPUT37), .A4(new_n384), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n386), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT38), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n394), .B(KEYINPUT38), .C1(new_n393), .C2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G141gat), .B(G148gat), .Z(new_n402));
  INV_X1    g201(.A(G155gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT2), .B1(new_n403), .B2(new_n316), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G155gat), .B(G162gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT3), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT68), .B(G113gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(G120gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G127gat), .B(G134gat), .ZN(new_n411));
  INV_X1    g210(.A(G113gat), .ZN(new_n412));
  INV_X1    g211(.A(G120gat), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT1), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT69), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g218(.A(new_n411), .B(KEYINPUT67), .Z(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n412), .B2(new_n413), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n417), .A2(new_n418), .B1(new_n421), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n407), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n407), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT74), .B(KEYINPUT4), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT5), .ZN(new_n433));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n408), .B2(new_n423), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n436), .B(new_n434), .C1(new_n437), .C2(new_n429), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n428), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n426), .ZN(new_n440));
  INV_X1    g239(.A(new_n434), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n438), .A2(KEYINPUT5), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n449), .B(KEYINPUT80), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  INV_X1    g256(.A(new_n449), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n444), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n458), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n456), .A2(new_n460), .B1(KEYINPUT6), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n392), .A2(new_n390), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n401), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n426), .A3(new_n434), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT39), .B(new_n466), .C1(new_n432), .C2(new_n434), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT81), .B(KEYINPUT39), .Z(new_n468));
  NAND4_X1  g267(.A1(new_n427), .A2(new_n441), .A3(new_n431), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(KEYINPUT82), .A3(new_n450), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT82), .B1(new_n469), .B2(new_n450), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT84), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n472), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n470), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT40), .A4(new_n467), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(new_n474), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n391), .B2(new_n389), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n392), .A2(new_n482), .A3(new_n390), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n454), .B2(new_n455), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G78gat), .B(G106gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT31), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(new_n258), .ZN(new_n491));
  INV_X1    g290(.A(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT3), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT29), .B1(new_n407), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n379), .A2(new_n495), .A3(KEYINPUT77), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT77), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n378), .B2(new_n494), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n376), .A2(new_n371), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n375), .A2(KEYINPUT76), .A3(new_n377), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT3), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n496), .B(new_n498), .C1(new_n503), .C2(new_n407), .ZN(new_n504));
  AND2_X1   g303(.A1(G228gat), .A2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n378), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n407), .B1(new_n513), .B2(new_n493), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n378), .A2(new_n494), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n514), .A2(new_n506), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n492), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  AOI211_X1 g317(.A(G22gat), .B(new_n516), .C1(new_n508), .C2(new_n510), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n491), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n510), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n509), .B1(new_n504), .B2(new_n506), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G22gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n511), .A2(new_n492), .A3(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n520), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n465), .A2(new_n488), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n460), .A2(new_n461), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n462), .A2(new_n459), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n532), .A2(new_n533), .B1(new_n485), .B2(new_n484), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n355), .A2(new_n537), .A3(new_n425), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n360), .A2(new_n425), .A3(new_n362), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT70), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n363), .A2(new_n423), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(G227gat), .A2(G233gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT33), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(KEYINPUT32), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G43gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G71gat), .ZN(new_n548));
  INV_X1    g347(.A(G99gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT32), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n542), .B2(new_n543), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(KEYINPUT33), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n555), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT71), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n556), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT34), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n551), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n542), .A2(new_n543), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT36), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n566), .B1(new_n560), .B2(new_n565), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n559), .A2(KEYINPUT34), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n564), .B1(new_n563), .B2(new_n551), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n572), .A2(new_n573), .B1(new_n543), .B2(new_n542), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT36), .B1(new_n574), .B2(new_n567), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n531), .B(new_n536), .C1(new_n571), .C2(new_n575), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n568), .A2(new_n570), .A3(new_n529), .ZN(new_n577));
  INV_X1    g376(.A(new_n486), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n463), .A2(KEYINPUT35), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n530), .A2(new_n574), .A3(new_n567), .A4(new_n534), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT35), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n323), .B1(new_n576), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT90), .B1(new_n228), .B2(new_n230), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n270), .B1(new_n585), .B2(KEYINPUT17), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT90), .B1(new_n298), .B2(new_n271), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n231), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT18), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n266), .A2(new_n271), .A3(new_n269), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT90), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n231), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n223), .A2(new_n226), .A3(new_n229), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n229), .B1(new_n223), .B2(new_n226), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n596), .A2(new_n271), .B1(new_n266), .B2(new_n269), .ZN(new_n597));
  OAI211_X1 g396(.A(KEYINPUT18), .B(new_n589), .C1(new_n593), .C2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n594), .A2(new_n595), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n270), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n589), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n600), .A2(new_n601), .A3(new_n607), .A4(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n589), .B1(new_n593), .B2(new_n597), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT18), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(new_n612), .A3(new_n607), .A4(new_n598), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT91), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n612), .ZN(new_n619));
  INV_X1    g418(.A(new_n607), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n613), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  INV_X1    g421(.A(G233gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n287), .A2(KEYINPUT98), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n215), .B2(new_n216), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n284), .A2(new_n285), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n628), .B(new_n626), .C1(new_n215), .C2(new_n216), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT10), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n299), .A2(new_n235), .A3(KEYINPUT10), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n625), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n624), .A3(new_n631), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT99), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(new_n343), .ZN(new_n640));
  INV_X1    g439(.A(G204gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n621), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n584), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n532), .A2(new_n533), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT100), .B(G1gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1324gat));
  NAND2_X1  g452(.A1(new_n225), .A2(new_n229), .ZN(new_n654));
  NAND2_X1  g453(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n578), .A2(new_n648), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n229), .B1(new_n648), .B2(new_n578), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  NOR2_X1   g458(.A1(new_n568), .A2(new_n570), .ZN(new_n660));
  AOI21_X1  g459(.A(G15gat), .B1(new_n648), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n571), .B2(new_n575), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n574), .A2(KEYINPUT36), .A3(new_n567), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(KEYINPUT101), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(G15gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n661), .B1(new_n648), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n529), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT102), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n648), .A2(new_n673), .A3(new_n529), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT43), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G22gat), .ZN(G1327gat));
  AOI21_X1  g476(.A(new_n322), .B1(new_n576), .B2(new_n583), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n245), .A2(new_n646), .A3(new_n621), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n294), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n650), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n685), .B(new_n322), .C1(new_n576), .C2(new_n583), .ZN(new_n686));
  INV_X1    g485(.A(new_n322), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n531), .A2(new_n536), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n666), .B2(new_n663), .ZN(new_n689));
  INV_X1    g488(.A(new_n583), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n686), .B1(new_n691), .B2(new_n685), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n679), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n294), .B1(new_n693), .B2(new_n649), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n684), .A2(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n249), .A3(new_n578), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT46), .Z(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n693), .B2(new_n486), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1329gat));
  OAI21_X1  g500(.A(G43gat), .B1(new_n693), .B2(new_n667), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n257), .A3(new_n660), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n702), .B(new_n703), .C1(KEYINPUT105), .C2(KEYINPUT47), .ZN(new_n704));
  NAND2_X1  g503(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1330gat));
  NAND3_X1  g505(.A1(new_n692), .A2(new_n529), .A3(new_n679), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n530), .A2(G50gat), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n707), .A2(G50gat), .B1(new_n680), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT48), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n709), .A2(KEYINPUT106), .A3(KEYINPUT48), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n709), .A2(new_n714), .A3(KEYINPUT48), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n709), .B2(KEYINPUT48), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n712), .A2(new_n713), .B1(new_n715), .B2(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n646), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n399), .A2(new_n400), .B1(new_n392), .B2(new_n390), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(new_n463), .B1(new_n481), .B2(new_n487), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n535), .B1(new_n720), .B2(new_n530), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n571), .A2(new_n575), .A3(new_n662), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT101), .B1(new_n664), .B2(new_n665), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n718), .B1(new_n724), .B2(new_n583), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n619), .A2(new_n620), .ZN(new_n726));
  INV_X1    g525(.A(new_n618), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n617), .A2(KEYINPUT91), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n323), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n650), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n486), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  AND2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT108), .ZN(G1333gat));
  NOR3_X1   g539(.A1(new_n731), .A2(new_n568), .A3(new_n570), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n663), .A2(G71gat), .A3(new_n666), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n741), .A2(G71gat), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n732), .A2(new_n529), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g545(.A1(new_n678), .A2(KEYINPUT44), .ZN(new_n747));
  INV_X1    g546(.A(new_n245), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n621), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n646), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n322), .B1(new_n724), .B2(new_n583), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n747), .B(new_n752), .C1(new_n753), .C2(KEYINPUT44), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n649), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n687), .B(new_n750), .C1(new_n689), .C2(new_n690), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n756), .A2(new_n757), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n761), .A2(new_n763), .A3(KEYINPUT111), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT111), .B1(new_n761), .B2(new_n763), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n281), .B(new_n646), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n755), .B1(new_n766), .B2(new_n649), .ZN(G1336gat));
  OAI21_X1  g566(.A(KEYINPUT112), .B1(new_n754), .B2(new_n486), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n692), .A2(new_n769), .A3(new_n578), .A4(new_n752), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n770), .A3(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n486), .A2(G92gat), .A3(new_n718), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n761), .A2(new_n763), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT113), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n771), .A2(new_n777), .A3(new_n772), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G92gat), .B1(new_n754), .B2(new_n486), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n753), .B2(new_n750), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n762), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n784), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n660), .A2(new_n549), .A3(new_n646), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT114), .Z(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n764), .B2(new_n765), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n754), .B2(new_n667), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  NOR3_X1   g589(.A1(new_n530), .A2(G106gat), .A3(new_n718), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n761), .A2(new_n763), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g592(.A(G106gat), .B1(new_n754), .B2(new_n530), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n762), .B2(new_n781), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT116), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(KEYINPUT115), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(KEYINPUT116), .ZN(new_n800));
  AND4_X1   g599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n795), .B1(new_n801), .B2(new_n793), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT10), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n628), .B1(new_n235), .B2(new_n626), .ZN(new_n804));
  INV_X1    g603(.A(new_n631), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(new_n624), .A3(new_n633), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n635), .A3(KEYINPUT54), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n807), .A2(new_n635), .A3(KEYINPUT117), .A4(KEYINPUT54), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n625), .C1(new_n632), .C2(new_n634), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n643), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT118), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(new_n817), .A3(new_n643), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n812), .A2(new_n819), .A3(KEYINPUT55), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n645), .A3(new_n729), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n606), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n588), .A2(new_n589), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n609), .A2(new_n611), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n646), .B(new_n829), .C1(new_n727), .C2(new_n728), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n687), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n613), .B2(new_n618), .ZN(new_n832));
  AOI22_X1  g631(.A1(new_n810), .A2(new_n811), .B1(new_n816), .B2(new_n818), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(KEYINPUT55), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n823), .A2(new_n645), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n322), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT119), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n823), .A2(new_n645), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n687), .A2(new_n839), .A3(new_n832), .A4(new_n822), .ZN(new_n840));
  INV_X1    g639(.A(new_n830), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(new_n812), .B2(new_n819), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n621), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(new_n839), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n838), .B(new_n840), .C1(new_n844), .C2(new_n687), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n748), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n730), .A2(new_n718), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n577), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n649), .A2(new_n578), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n729), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G113gat), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n409), .B2(new_n853), .ZN(G1340gat));
  NOR2_X1   g654(.A1(new_n851), .A2(new_n718), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(new_n413), .ZN(G1341gat));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n245), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g658(.A1(new_n851), .A2(new_n322), .ZN(new_n860));
  NOR2_X1   g659(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n861));
  AND2_X1   g660(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n860), .B2(new_n861), .ZN(G1343gat));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n323), .A2(new_n646), .A3(new_n729), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n824), .A2(new_n830), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n836), .B1(new_n867), .B2(new_n322), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n245), .B1(new_n868), .B2(new_n838), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n866), .B1(new_n869), .B2(new_n837), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT120), .B(new_n865), .C1(new_n870), .C2(new_n530), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n530), .B1(new_n846), .B2(new_n847), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n847), .B1(new_n245), .B2(new_n868), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .A3(new_n529), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n667), .A2(new_n850), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n621), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  INV_X1    g681(.A(new_n873), .ZN(new_n883));
  NOR4_X1   g682(.A1(new_n878), .A2(new_n883), .A3(G141gat), .A4(new_n621), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n887), .A3(new_n879), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n877), .B2(new_n879), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n729), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(G141gat), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n882), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n880), .A2(KEYINPUT121), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n621), .B1(new_n895), .B2(new_n888), .ZN(new_n896));
  INV_X1    g695(.A(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT122), .B1(new_n898), .B2(KEYINPUT58), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n886), .B1(new_n894), .B2(new_n899), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n878), .A2(new_n883), .ZN(new_n901));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n646), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n718), .B1(new_n895), .B2(new_n888), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(KEYINPUT59), .A3(new_n902), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n875), .A2(new_n529), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n865), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n646), .ZN(new_n910));
  OAI21_X1  g709(.A(G148gat), .B1(new_n910), .B2(new_n878), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT59), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n905), .B2(new_n912), .ZN(G1345gat));
  AOI21_X1  g712(.A(G155gat), .B1(new_n901), .B2(new_n245), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n888), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n245), .A2(G155gat), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT123), .Z(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(G1346gat));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n316), .A3(new_n687), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n322), .B1(new_n895), .B2(new_n888), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n316), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n577), .A2(new_n578), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT125), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n870), .A2(new_n650), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n342), .A3(new_n729), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n650), .A2(new_n486), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n849), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G169gat), .B1(new_n929), .B2(new_n621), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n929), .B2(new_n718), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n870), .A2(new_n650), .A3(new_n718), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n343), .A3(new_n924), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1349gat));
  NAND3_X1  g734(.A1(new_n926), .A2(new_n337), .A3(new_n245), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n929), .B2(new_n748), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT126), .ZN(new_n939));
  XOR2_X1   g738(.A(new_n939), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n929), .B2(new_n322), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT61), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n338), .A3(new_n687), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1351gat));
  AOI211_X1 g743(.A(new_n486), .B(new_n530), .C1(new_n663), .C2(new_n666), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n945), .A2(new_n925), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n729), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n667), .A2(new_n928), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n907), .B2(new_n908), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(new_n729), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n951), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n945), .A3(new_n641), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT62), .Z(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n910), .B2(new_n949), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n946), .A2(new_n367), .A3(new_n245), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n950), .A2(new_n245), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n946), .B2(new_n687), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n322), .A2(new_n368), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n950), .B2(new_n964), .ZN(G1355gat));
endmodule


