

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760;

  INV_X2 U372 ( .A(G953), .ZN(n737) );
  XNOR2_X1 U373 ( .A(n609), .B(KEYINPUT33), .ZN(n661) );
  INV_X2 U374 ( .A(n630), .ZN(n729) );
  XNOR2_X2 U375 ( .A(n459), .B(n458), .ZN(n630) );
  INV_X2 U376 ( .A(G143), .ZN(n473) );
  NOR2_X2 U377 ( .A1(n370), .A2(n667), .ZN(n673) );
  XNOR2_X2 U378 ( .A(n433), .B(n372), .ZN(n667) );
  XNOR2_X2 U379 ( .A(n489), .B(KEYINPUT35), .ZN(n758) );
  XOR2_X2 U380 ( .A(G131), .B(KEYINPUT66), .Z(n553) );
  XNOR2_X2 U381 ( .A(n412), .B(n472), .ZN(n507) );
  AND2_X1 U382 ( .A1(n394), .A2(n389), .ZN(n388) );
  XNOR2_X1 U383 ( .A(n492), .B(KEYINPUT96), .ZN(n637) );
  AND2_X1 U384 ( .A1(n597), .A2(n353), .ZN(n602) );
  AND2_X1 U385 ( .A1(n359), .A2(n474), .ZN(n349) );
  XNOR2_X1 U386 ( .A(n682), .B(n562), .ZN(n608) );
  NOR2_X1 U387 ( .A1(n575), .A2(n581), .ZN(n669) );
  NAND2_X1 U388 ( .A1(n401), .A2(n397), .ZN(n446) );
  XNOR2_X1 U389 ( .A(n558), .B(n557), .ZN(n581) );
  OR2_X1 U390 ( .A1(n517), .A2(n481), .ZN(n480) );
  XNOR2_X1 U391 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U392 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U393 ( .A(n555), .B(n430), .ZN(n714) );
  XNOR2_X1 U394 ( .A(n386), .B(n508), .ZN(n385) );
  XNOR2_X1 U395 ( .A(n418), .B(G125), .ZN(n531) );
  XNOR2_X1 U396 ( .A(n487), .B(KEYINPUT3), .ZN(n503) );
  XNOR2_X1 U397 ( .A(KEYINPUT87), .B(G110), .ZN(n735) );
  NOR2_X1 U398 ( .A1(G953), .A2(G237), .ZN(n551) );
  XNOR2_X1 U399 ( .A(G101), .B(G119), .ZN(n487) );
  XNOR2_X1 U400 ( .A(n387), .B(n384), .ZN(n465) );
  XNOR2_X1 U401 ( .A(n385), .B(n506), .ZN(n384) );
  XNOR2_X1 U402 ( .A(n423), .B(n571), .ZN(n760) );
  BUF_X1 U403 ( .A(n706), .Z(n348) );
  XNOR2_X1 U404 ( .A(n465), .B(n734), .ZN(n706) );
  NOR2_X1 U405 ( .A1(n585), .A2(n467), .ZN(n394) );
  AND2_X1 U406 ( .A1(n757), .A2(n577), .ZN(n390) );
  NAND2_X1 U407 ( .A1(n434), .A2(n457), .ZN(n411) );
  NOR2_X1 U408 ( .A1(n456), .A2(n625), .ZN(n408) );
  NAND2_X1 U409 ( .A1(n482), .A2(n399), .ZN(n481) );
  XNOR2_X1 U410 ( .A(n743), .B(n418), .ZN(n405) );
  OR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n519) );
  NAND2_X1 U412 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U413 ( .A1(n518), .A2(G902), .ZN(n484) );
  INV_X1 U414 ( .A(KEYINPUT30), .ZN(n478) );
  NAND2_X1 U415 ( .A1(n400), .A2(n399), .ZN(n398) );
  XNOR2_X1 U416 ( .A(n501), .B(n498), .ZN(n416) );
  AND2_X1 U417 ( .A1(n551), .A2(G210), .ZN(n501) );
  XNOR2_X1 U418 ( .A(n352), .B(G116), .ZN(n417) );
  XOR2_X1 U419 ( .A(G137), .B(KEYINPUT5), .Z(n499) );
  NOR2_X1 U420 ( .A1(n659), .A2(n594), .ZN(n595) );
  XNOR2_X1 U421 ( .A(n426), .B(G140), .ZN(n536) );
  INV_X1 U422 ( .A(G137), .ZN(n426) );
  XNOR2_X1 U423 ( .A(n537), .B(n538), .ZN(n404) );
  XNOR2_X1 U424 ( .A(n382), .B(n466), .ZN(n381) );
  INV_X1 U425 ( .A(KEYINPUT45), .ZN(n458) );
  INV_X1 U426 ( .A(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n605) );
  INV_X1 U428 ( .A(KEYINPUT22), .ZN(n368) );
  NOR2_X1 U429 ( .A1(n620), .A2(n462), .ZN(n369) );
  NAND2_X1 U430 ( .A1(n669), .A2(n351), .ZN(n462) );
  XNOR2_X1 U431 ( .A(n561), .B(KEYINPUT6), .ZN(n562) );
  INV_X1 U432 ( .A(KEYINPUT100), .ZN(n561) );
  XNOR2_X1 U433 ( .A(G128), .B(G119), .ZN(n532) );
  XNOR2_X1 U434 ( .A(n536), .B(n450), .ZN(n449) );
  XNOR2_X1 U435 ( .A(n451), .B(n535), .ZN(n450) );
  INV_X1 U436 ( .A(KEYINPUT24), .ZN(n535) );
  XNOR2_X1 U437 ( .A(KEYINPUT78), .B(KEYINPUT23), .ZN(n451) );
  INV_X1 U438 ( .A(KEYINPUT10), .ZN(n452) );
  XNOR2_X1 U439 ( .A(n380), .B(n378), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n379), .B(KEYINPUT12), .ZN(n378) );
  NAND2_X1 U441 ( .A1(n551), .A2(G214), .ZN(n380) );
  INV_X1 U442 ( .A(KEYINPUT97), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n374) );
  XNOR2_X1 U444 ( .A(KEYINPUT11), .B(G122), .ZN(n376) );
  XNOR2_X1 U445 ( .A(G143), .B(G140), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n507), .B(n523), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n371), .B(KEYINPUT41), .ZN(n690) );
  XNOR2_X1 U448 ( .A(n588), .B(n431), .ZN(n566) );
  INV_X1 U449 ( .A(KEYINPUT107), .ZN(n431) );
  NAND2_X1 U450 ( .A1(n560), .A2(n589), .ZN(n455) );
  BUF_X1 U451 ( .A(n677), .Z(n424) );
  XNOR2_X1 U452 ( .A(n455), .B(KEYINPUT19), .ZN(n597) );
  NOR2_X1 U453 ( .A1(n605), .A2(n616), .ZN(n603) );
  XNOR2_X1 U454 ( .A(n427), .B(G478), .ZN(n580) );
  NOR2_X1 U455 ( .A1(n720), .A2(G902), .ZN(n427) );
  NOR2_X1 U456 ( .A1(n714), .A2(G902), .ZN(n557) );
  XNOR2_X1 U457 ( .A(n471), .B(n364), .ZN(n470) );
  XNOR2_X1 U458 ( .A(n582), .B(n583), .ZN(n367) );
  XOR2_X1 U459 ( .A(G107), .B(G104), .Z(n521) );
  XNOR2_X1 U460 ( .A(n536), .B(n425), .ZN(n744) );
  INV_X1 U461 ( .A(KEYINPUT90), .ZN(n425) );
  XOR2_X1 U462 ( .A(KEYINPUT17), .B(KEYINPUT76), .Z(n508) );
  XNOR2_X1 U463 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U464 ( .A(KEYINPUT18), .ZN(n504) );
  INV_X1 U465 ( .A(KEYINPUT4), .ZN(n472) );
  XNOR2_X1 U466 ( .A(n735), .B(KEYINPUT68), .ZN(n523) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n511) );
  XNOR2_X1 U468 ( .A(n510), .B(n509), .ZN(n592) );
  AND2_X1 U469 ( .A1(n476), .A2(n475), .ZN(n474) );
  OR2_X1 U470 ( .A1(n589), .A2(n478), .ZN(n475) );
  NAND2_X1 U471 ( .A1(n477), .A2(n361), .ZN(n476) );
  NOR2_X1 U472 ( .A1(n676), .A2(n563), .ZN(n396) );
  NAND2_X1 U473 ( .A1(G469), .A2(G902), .ZN(n402) );
  NAND2_X1 U474 ( .A1(n596), .A2(n351), .ZN(n676) );
  XNOR2_X1 U475 ( .A(n405), .B(n502), .ZN(n517) );
  XNOR2_X1 U476 ( .A(n419), .B(n500), .ZN(n502) );
  XNOR2_X1 U477 ( .A(n416), .B(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n631), .B(n436), .ZN(n742) );
  INV_X1 U479 ( .A(KEYINPUT79), .ZN(n436) );
  AND2_X1 U480 ( .A1(n381), .A2(n595), .ZN(n631) );
  XNOR2_X1 U481 ( .A(n464), .B(n463), .ZN(n734) );
  XNOR2_X1 U482 ( .A(n552), .B(n486), .ZN(n463) );
  XNOR2_X1 U483 ( .A(n503), .B(n546), .ZN(n464) );
  INV_X1 U484 ( .A(KEYINPUT16), .ZN(n486) );
  XNOR2_X1 U485 ( .A(G134), .B(KEYINPUT98), .ZN(n429) );
  XOR2_X1 U486 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n548) );
  XNOR2_X1 U487 ( .A(n488), .B(G122), .ZN(n546) );
  XNOR2_X1 U488 ( .A(G116), .B(G107), .ZN(n488) );
  XNOR2_X1 U489 ( .A(G902), .B(KEYINPUT15), .ZN(n628) );
  NOR2_X2 U490 ( .A1(n630), .A2(n626), .ZN(n627) );
  XNOR2_X1 U491 ( .A(n422), .B(KEYINPUT80), .ZN(n626) );
  BUF_X1 U492 ( .A(n592), .Z(n433) );
  XNOR2_X1 U493 ( .A(n448), .B(n453), .ZN(n726) );
  XNOR2_X1 U494 ( .A(n454), .B(n534), .ZN(n453) );
  XNOR2_X1 U495 ( .A(n556), .B(n449), .ZN(n448) );
  XNOR2_X1 U496 ( .A(n554), .B(n373), .ZN(n555) );
  XNOR2_X1 U497 ( .A(n377), .B(n374), .ZN(n373) );
  XNOR2_X1 U498 ( .A(n576), .B(n428), .ZN(n757) );
  XNOR2_X1 U499 ( .A(KEYINPUT42), .B(KEYINPUT106), .ZN(n428) );
  NOR2_X1 U500 ( .A1(n586), .A2(n651), .ZN(n423) );
  XNOR2_X1 U501 ( .A(n567), .B(n432), .ZN(n568) );
  XNOR2_X1 U502 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n432) );
  INV_X1 U503 ( .A(KEYINPUT34), .ZN(n420) );
  XNOR2_X1 U504 ( .A(n607), .B(KEYINPUT32), .ZN(n383) );
  XNOR2_X1 U505 ( .A(n579), .B(KEYINPUT77), .ZN(n648) );
  NAND2_X1 U506 ( .A1(n414), .A2(n360), .ZN(n641) );
  XNOR2_X1 U507 ( .A(n603), .B(KEYINPUT102), .ZN(n414) );
  INV_X1 U508 ( .A(n679), .ZN(n413) );
  NOR2_X1 U509 ( .A1(n616), .A2(n615), .ZN(n635) );
  NAND2_X1 U510 ( .A1(n470), .A2(n469), .ZN(n468) );
  NAND2_X1 U511 ( .A1(n438), .A2(n469), .ZN(n437) );
  XNOR2_X1 U512 ( .A(n439), .B(n363), .ZN(n438) );
  NAND2_X1 U513 ( .A1(n415), .A2(n361), .ZN(n350) );
  XNOR2_X1 U514 ( .A(n573), .B(KEYINPUT28), .ZN(n574) );
  XOR2_X1 U515 ( .A(KEYINPUT21), .B(n542), .Z(n351) );
  XOR2_X1 U516 ( .A(G113), .B(KEYINPUT95), .Z(n352) );
  OR2_X1 U517 ( .A1(n600), .A2(n599), .ZN(n353) );
  AND2_X1 U518 ( .A1(n575), .A2(n581), .ZN(n354) );
  AND2_X1 U519 ( .A1(n396), .A2(n446), .ZN(n355) );
  NAND2_X1 U520 ( .A1(n395), .A2(n446), .ZN(n356) );
  AND2_X1 U521 ( .A1(n446), .A2(n574), .ZN(n357) );
  AND2_X1 U522 ( .A1(n480), .A2(KEYINPUT30), .ZN(n358) );
  AND2_X1 U523 ( .A1(n350), .A2(n479), .ZN(n359) );
  INV_X1 U524 ( .A(G902), .ZN(n399) );
  INV_X2 U525 ( .A(G146), .ZN(n418) );
  AND2_X1 U526 ( .A1(n618), .A2(n413), .ZN(n360) );
  AND2_X1 U527 ( .A1(n589), .A2(n478), .ZN(n361) );
  AND2_X1 U528 ( .A1(n595), .A2(KEYINPUT2), .ZN(n362) );
  INV_X1 U529 ( .A(n574), .ZN(n447) );
  XOR2_X1 U530 ( .A(n348), .B(n495), .Z(n363) );
  XOR2_X1 U531 ( .A(n517), .B(KEYINPUT62), .Z(n364) );
  XNOR2_X1 U532 ( .A(n531), .B(n452), .ZN(n556) );
  INV_X1 U533 ( .A(n556), .ZN(n430) );
  XNOR2_X1 U534 ( .A(n507), .B(n497), .ZN(n743) );
  NOR2_X1 U535 ( .A1(G952), .A2(n737), .ZN(n728) );
  INV_X1 U536 ( .A(n728), .ZN(n469) );
  XNOR2_X1 U537 ( .A(KEYINPUT81), .B(KEYINPUT56), .ZN(n365) );
  XOR2_X1 U538 ( .A(n634), .B(KEYINPUT86), .Z(n366) );
  NAND2_X1 U539 ( .A1(n367), .A2(n584), .ZN(n467) );
  NAND2_X1 U540 ( .A1(n391), .A2(n388), .ZN(n382) );
  NAND2_X1 U541 ( .A1(n485), .A2(n484), .ZN(n415) );
  NAND2_X1 U542 ( .A1(n597), .A2(n578), .ZN(n579) );
  NAND2_X1 U543 ( .A1(n381), .A2(n362), .ZN(n422) );
  INV_X1 U544 ( .A(n669), .ZN(n370) );
  NAND2_X1 U545 ( .A1(n673), .A2(n589), .ZN(n371) );
  INV_X1 U546 ( .A(KEYINPUT38), .ZN(n372) );
  NAND2_X1 U547 ( .A1(n383), .A2(n641), .ZN(n612) );
  XNOR2_X1 U548 ( .A(n383), .B(G119), .ZN(n759) );
  NOR2_X2 U549 ( .A1(n605), .A2(n608), .ZN(n614) );
  XNOR2_X2 U550 ( .A(n602), .B(n601), .ZN(n620) );
  INV_X1 U551 ( .A(n531), .ZN(n386) );
  XNOR2_X2 U552 ( .A(n473), .B(G128), .ZN(n412) );
  NAND2_X1 U553 ( .A1(n760), .A2(n390), .ZN(n389) );
  NOR2_X1 U554 ( .A1(n393), .A2(n392), .ZN(n391) );
  NOR2_X1 U555 ( .A1(n757), .A2(n577), .ZN(n392) );
  NOR2_X1 U556 ( .A1(n760), .A2(n577), .ZN(n393) );
  INV_X1 U557 ( .A(n676), .ZN(n395) );
  OR2_X1 U558 ( .A1(n707), .A2(n398), .ZN(n397) );
  INV_X1 U559 ( .A(G469), .ZN(n400) );
  AND2_X1 U560 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U561 ( .A1(n707), .A2(G469), .ZN(n403) );
  NAND2_X1 U562 ( .A1(n404), .A2(G221), .ZN(n454) );
  NAND2_X1 U563 ( .A1(n404), .A2(G217), .ZN(n547) );
  XNOR2_X1 U564 ( .A(n526), .B(n405), .ZN(n707) );
  NAND2_X1 U565 ( .A1(n406), .A2(G475), .ZN(n716) );
  NAND2_X1 U566 ( .A1(n406), .A2(G478), .ZN(n722) );
  NAND2_X1 U567 ( .A1(n406), .A2(G210), .ZN(n439) );
  NAND2_X1 U568 ( .A1(n406), .A2(G472), .ZN(n471) );
  NAND2_X1 U569 ( .A1(n406), .A2(G469), .ZN(n710) );
  NAND2_X1 U570 ( .A1(n406), .A2(G217), .ZN(n725) );
  AND2_X4 U571 ( .A1(n491), .A2(n662), .ZN(n406) );
  AND2_X1 U572 ( .A1(n446), .A2(n447), .ZN(n444) );
  XNOR2_X1 U573 ( .A(n446), .B(n407), .ZN(n677) );
  NAND2_X1 U574 ( .A1(n408), .A2(n613), .ZN(n410) );
  NAND2_X1 U575 ( .A1(n410), .A2(n409), .ZN(n461) );
  NAND2_X1 U576 ( .A1(n411), .A2(n613), .ZN(n409) );
  XNOR2_X1 U577 ( .A(n412), .B(n429), .ZN(n545) );
  NAND2_X1 U578 ( .A1(n661), .A2(n435), .ZN(n421) );
  INV_X1 U579 ( .A(n415), .ZN(n483) );
  XNOR2_X1 U580 ( .A(n421), .B(n420), .ZN(n490) );
  XNOR2_X1 U581 ( .A(n611), .B(KEYINPUT69), .ZN(n460) );
  XNOR2_X1 U582 ( .A(n539), .B(n540), .ZN(n596) );
  NAND2_X1 U583 ( .A1(n349), .A2(n355), .ZN(n543) );
  NAND2_X1 U584 ( .A1(n648), .A2(n665), .ZN(n582) );
  NAND2_X1 U585 ( .A1(n565), .A2(n608), .ZN(n588) );
  AND2_X2 U586 ( .A1(n663), .A2(n629), .ZN(n491) );
  NAND2_X1 U587 ( .A1(n625), .A2(KEYINPUT83), .ZN(n434) );
  INV_X1 U588 ( .A(n661), .ZN(n675) );
  INV_X1 U589 ( .A(n620), .ZN(n435) );
  XNOR2_X1 U590 ( .A(n437), .B(n365), .ZN(G51) );
  NAND2_X1 U591 ( .A1(n442), .A2(n440), .ZN(n578) );
  NAND2_X1 U592 ( .A1(n444), .A2(n441), .ZN(n440) );
  NOR2_X1 U593 ( .A1(n572), .A2(n618), .ZN(n441) );
  NAND2_X1 U594 ( .A1(n357), .A2(n443), .ZN(n442) );
  NAND2_X1 U595 ( .A1(n445), .A2(n682), .ZN(n443) );
  INV_X1 U596 ( .A(n572), .ZN(n445) );
  NOR2_X1 U597 ( .A1(n566), .A2(n455), .ZN(n567) );
  OR2_X1 U598 ( .A1(n635), .A2(KEYINPUT83), .ZN(n456) );
  NAND2_X1 U599 ( .A1(n635), .A2(KEYINPUT83), .ZN(n457) );
  NAND2_X1 U600 ( .A1(n461), .A2(n460), .ZN(n459) );
  NAND2_X2 U601 ( .A1(n483), .A2(n480), .ZN(n682) );
  INV_X1 U602 ( .A(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U603 ( .A(n468), .B(n366), .ZN(G57) );
  INV_X1 U604 ( .A(n480), .ZN(n477) );
  NAND2_X1 U605 ( .A1(n358), .A2(n483), .ZN(n479) );
  INV_X1 U606 ( .A(n518), .ZN(n482) );
  NAND2_X1 U607 ( .A1(n517), .A2(n518), .ZN(n485) );
  NAND2_X1 U608 ( .A1(n490), .A2(n354), .ZN(n489) );
  XNOR2_X2 U609 ( .A(n627), .B(KEYINPUT73), .ZN(n662) );
  NAND2_X1 U610 ( .A1(n637), .A2(n653), .ZN(n622) );
  NAND2_X1 U611 ( .A1(n493), .A2(n618), .ZN(n492) );
  XNOR2_X1 U612 ( .A(n617), .B(n494), .ZN(n493) );
  INV_X1 U613 ( .A(KEYINPUT93), .ZN(n494) );
  XNOR2_X1 U614 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U615 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U616 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n495) );
  INV_X1 U617 ( .A(n660), .ZN(n594) );
  XNOR2_X1 U618 ( .A(n503), .B(n499), .ZN(n500) );
  XNOR2_X1 U619 ( .A(n553), .B(n496), .ZN(n497) );
  INV_X1 U620 ( .A(KEYINPUT104), .ZN(n573) );
  INV_X1 U621 ( .A(KEYINPUT63), .ZN(n634) );
  XOR2_X1 U622 ( .A(G134), .B(KEYINPUT67), .Z(n496) );
  XNOR2_X1 U623 ( .A(KEYINPUT72), .B(KEYINPUT94), .ZN(n498) );
  XOR2_X1 U624 ( .A(G113), .B(G104), .Z(n552) );
  NAND2_X1 U625 ( .A1(G224), .A2(n737), .ZN(n505) );
  NAND2_X1 U626 ( .A1(n706), .A2(n628), .ZN(n510) );
  NAND2_X1 U627 ( .A1(G210), .A2(n519), .ZN(n509) );
  XNOR2_X1 U628 ( .A(n511), .B(KEYINPUT88), .ZN(n512) );
  XNOR2_X1 U629 ( .A(KEYINPUT14), .B(n512), .ZN(n514) );
  NAND2_X1 U630 ( .A1(n514), .A2(G952), .ZN(n513) );
  XOR2_X1 U631 ( .A(KEYINPUT89), .B(n513), .Z(n697) );
  NOR2_X1 U632 ( .A1(G953), .A2(n697), .ZN(n600) );
  AND2_X1 U633 ( .A1(n514), .A2(G953), .ZN(n515) );
  NAND2_X1 U634 ( .A1(G902), .A2(n515), .ZN(n598) );
  NOR2_X1 U635 ( .A1(G900), .A2(n598), .ZN(n516) );
  NOR2_X1 U636 ( .A1(n600), .A2(n516), .ZN(n563) );
  XNOR2_X1 U637 ( .A(G472), .B(KEYINPUT70), .ZN(n518) );
  NAND2_X1 U638 ( .A1(G214), .A2(n519), .ZN(n589) );
  NAND2_X1 U639 ( .A1(G227), .A2(n737), .ZN(n520) );
  XNOR2_X1 U640 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U641 ( .A(n522), .B(n744), .Z(n525) );
  XNOR2_X1 U642 ( .A(G101), .B(n523), .ZN(n524) );
  XNOR2_X1 U643 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U644 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n529) );
  NAND2_X1 U645 ( .A1(G234), .A2(n628), .ZN(n527) );
  XNOR2_X1 U646 ( .A(KEYINPUT20), .B(n527), .ZN(n541) );
  NAND2_X1 U647 ( .A1(G217), .A2(n541), .ZN(n528) );
  XNOR2_X1 U648 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U649 ( .A(KEYINPUT92), .B(n530), .ZN(n540) );
  XOR2_X1 U650 ( .A(KEYINPUT91), .B(G110), .Z(n533) );
  XNOR2_X1 U651 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n737), .A2(G234), .ZN(n538) );
  XNOR2_X1 U653 ( .A(KEYINPUT8), .B(KEYINPUT65), .ZN(n537) );
  NOR2_X1 U654 ( .A1(G902), .A2(n726), .ZN(n539) );
  NAND2_X1 U655 ( .A1(n541), .A2(G221), .ZN(n542) );
  XNOR2_X1 U656 ( .A(n543), .B(KEYINPUT74), .ZN(n569) );
  OR2_X1 U657 ( .A1(n433), .A2(n569), .ZN(n544) );
  XNOR2_X1 U658 ( .A(KEYINPUT103), .B(n544), .ZN(n559) );
  XNOR2_X1 U659 ( .A(n546), .B(n545), .ZN(n550) );
  XNOR2_X1 U660 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U661 ( .A(n550), .B(n549), .ZN(n720) );
  INV_X1 U662 ( .A(n580), .ZN(n575) );
  XNOR2_X1 U663 ( .A(KEYINPUT13), .B(G475), .ZN(n558) );
  XNOR2_X1 U664 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U665 ( .A1(n559), .A2(n354), .ZN(n647) );
  INV_X1 U666 ( .A(n592), .ZN(n560) );
  INV_X1 U667 ( .A(n589), .ZN(n671) );
  NAND2_X1 U668 ( .A1(n581), .A2(n580), .ZN(n651) );
  NOR2_X1 U669 ( .A1(n596), .A2(n563), .ZN(n564) );
  NAND2_X1 U670 ( .A1(n564), .A2(n351), .ZN(n572) );
  NOR2_X1 U671 ( .A1(n651), .A2(n572), .ZN(n565) );
  INV_X1 U672 ( .A(n424), .ZN(n616) );
  NAND2_X1 U673 ( .A1(n568), .A2(n616), .ZN(n657) );
  NAND2_X1 U674 ( .A1(n647), .A2(n657), .ZN(n585) );
  NOR2_X1 U675 ( .A1(n569), .A2(n667), .ZN(n570) );
  XNOR2_X1 U676 ( .A(n570), .B(KEYINPUT39), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n571) );
  INV_X1 U678 ( .A(n682), .ZN(n618) );
  NAND2_X1 U679 ( .A1(n578), .A2(n690), .ZN(n576) );
  XOR2_X1 U680 ( .A(KEYINPUT46), .B(KEYINPUT82), .Z(n577) );
  NOR2_X1 U681 ( .A1(KEYINPUT71), .A2(KEYINPUT47), .ZN(n583) );
  NOR2_X1 U682 ( .A1(n581), .A2(n580), .ZN(n642) );
  INV_X1 U683 ( .A(n642), .ZN(n654) );
  XOR2_X1 U684 ( .A(KEYINPUT99), .B(n654), .Z(n587) );
  NAND2_X1 U685 ( .A1(n587), .A2(n651), .ZN(n665) );
  NAND2_X1 U686 ( .A1(KEYINPUT71), .A2(KEYINPUT47), .ZN(n584) );
  NOR2_X1 U687 ( .A1(n587), .A2(n586), .ZN(n659) );
  NOR2_X1 U688 ( .A1(n616), .A2(n588), .ZN(n590) );
  NAND2_X1 U689 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U690 ( .A(n591), .B(KEYINPUT43), .ZN(n593) );
  NAND2_X1 U691 ( .A1(n593), .A2(n433), .ZN(n660) );
  BUF_X1 U692 ( .A(n596), .Z(n679) );
  NOR2_X1 U693 ( .A1(G898), .A2(n598), .ZN(n599) );
  XNOR2_X1 U694 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n601) );
  NOR2_X1 U695 ( .A1(n679), .A2(n424), .ZN(n604) );
  XOR2_X1 U696 ( .A(KEYINPUT101), .B(n604), .Z(n606) );
  NAND2_X1 U697 ( .A1(n606), .A2(n614), .ZN(n607) );
  NOR2_X1 U698 ( .A1(n677), .A2(n676), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n619), .A2(n608), .ZN(n609) );
  OR2_X2 U700 ( .A1(n758), .A2(KEYINPUT44), .ZN(n610) );
  NOR2_X2 U701 ( .A1(n612), .A2(n610), .ZN(n611) );
  NAND2_X1 U702 ( .A1(n612), .A2(KEYINPUT44), .ZN(n613) );
  NAND2_X1 U703 ( .A1(n679), .A2(n614), .ZN(n615) );
  NAND2_X1 U704 ( .A1(KEYINPUT44), .A2(n758), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n620), .A2(n356), .ZN(n617) );
  NAND2_X1 U706 ( .A1(n619), .A2(n682), .ZN(n687) );
  NOR2_X1 U707 ( .A1(n687), .A2(n620), .ZN(n621) );
  XNOR2_X1 U708 ( .A(n621), .B(KEYINPUT31), .ZN(n653) );
  NAND2_X1 U709 ( .A1(n622), .A2(n665), .ZN(n623) );
  INV_X1 U710 ( .A(n628), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n729), .A2(n742), .ZN(n633) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n663) );
  XOR2_X1 U714 ( .A(G101), .B(n635), .Z(G3) );
  NOR2_X1 U715 ( .A1(n637), .A2(n651), .ZN(n636) );
  XOR2_X1 U716 ( .A(G104), .B(n636), .Z(G6) );
  NOR2_X1 U717 ( .A1(n637), .A2(n654), .ZN(n639) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U720 ( .A(G107), .B(n640), .ZN(G9) );
  XNOR2_X1 U721 ( .A(n641), .B(G110), .ZN(G12) );
  XOR2_X1 U722 ( .A(KEYINPUT29), .B(KEYINPUT109), .Z(n644) );
  NAND2_X1 U723 ( .A1(n648), .A2(n642), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n644), .B(n643), .ZN(n646) );
  XOR2_X1 U725 ( .A(G128), .B(KEYINPUT108), .Z(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(G30) );
  XNOR2_X1 U727 ( .A(G143), .B(n647), .ZN(G45) );
  INV_X1 U728 ( .A(n651), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U730 ( .A(G146), .B(n650), .ZN(G48) );
  NOR2_X1 U731 ( .A1(n651), .A2(n653), .ZN(n652) );
  XOR2_X1 U732 ( .A(G113), .B(n652), .Z(G15) );
  NOR2_X1 U733 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U734 ( .A(G116), .B(n655), .Z(G18) );
  XOR2_X1 U735 ( .A(KEYINPUT110), .B(KEYINPUT37), .Z(n656) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(G125), .B(n658), .ZN(G27) );
  XOR2_X1 U738 ( .A(G134), .B(n659), .Z(G36) );
  XNOR2_X1 U739 ( .A(G140), .B(n660), .ZN(G42) );
  XNOR2_X1 U740 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n705) );
  NAND2_X1 U741 ( .A1(n661), .A2(n690), .ZN(n702) );
  NAND2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n737), .A2(n664), .ZN(n700) );
  INV_X1 U744 ( .A(n665), .ZN(n666) );
  NOR2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U747 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U749 ( .A1(n675), .A2(n674), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n424), .A2(n676), .ZN(n678) );
  XNOR2_X1 U751 ( .A(KEYINPUT50), .B(n678), .ZN(n685) );
  NOR2_X1 U752 ( .A1(n679), .A2(n351), .ZN(n681) );
  XNOR2_X1 U753 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n680) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(n683) );
  NOR2_X1 U755 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U758 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U760 ( .A(KEYINPUT112), .B(n691), .Z(n692) );
  NOR2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U762 ( .A(n694), .B(KEYINPUT113), .Z(n695) );
  XNOR2_X1 U763 ( .A(KEYINPUT52), .B(n695), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(KEYINPUT114), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U768 ( .A(n703), .B(KEYINPUT53), .ZN(n704) );
  XNOR2_X1 U769 ( .A(n705), .B(n704), .ZN(G75) );
  XNOR2_X1 U770 ( .A(KEYINPUT58), .B(KEYINPUT117), .ZN(n709) );
  XNOR2_X1 U771 ( .A(n707), .B(KEYINPUT57), .ZN(n708) );
  XNOR2_X1 U772 ( .A(n709), .B(n708), .ZN(n711) );
  XNOR2_X1 U773 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U774 ( .A1(n728), .A2(n712), .ZN(G54) );
  XOR2_X1 U775 ( .A(KEYINPUT59), .B(KEYINPUT64), .Z(n713) );
  NOR2_X2 U776 ( .A1(n717), .A2(n728), .ZN(n718) );
  XNOR2_X1 U777 ( .A(n718), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U778 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n719) );
  NOR2_X2 U779 ( .A1(n723), .A2(n728), .ZN(n724) );
  XNOR2_X1 U780 ( .A(n724), .B(KEYINPUT120), .ZN(G63) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U783 ( .A1(n737), .A2(n729), .ZN(n733) );
  NAND2_X1 U784 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U785 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n731), .A2(G898), .ZN(n732) );
  NAND2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n741) );
  XNOR2_X1 U788 ( .A(n734), .B(KEYINPUT121), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n735), .B(n736), .ZN(n739) );
  NOR2_X1 U790 ( .A1(G898), .A2(n737), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n741), .B(n740), .ZN(G69) );
  XNOR2_X1 U793 ( .A(n742), .B(KEYINPUT124), .ZN(n748) );
  XOR2_X1 U794 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n746) );
  XOR2_X1 U795 ( .A(n744), .B(n430), .Z(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n743), .B(n747), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n748), .B(n751), .ZN(n749) );
  NOR2_X1 U799 ( .A1(G953), .A2(n749), .ZN(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(KEYINPUT125), .ZN(n755) );
  XNOR2_X1 U801 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U803 ( .A1(G953), .A2(n753), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U805 ( .A(G137), .B(KEYINPUT127), .Z(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(G39) );
  XOR2_X1 U807 ( .A(n758), .B(G122), .Z(G24) );
  XNOR2_X1 U808 ( .A(n759), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U809 ( .A(n760), .B(G131), .ZN(G33) );
endmodule

