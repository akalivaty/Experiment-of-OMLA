//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n592, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT67), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n465), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n464), .A2(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT66), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n470), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n469), .A2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n466), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n485), .A2(G126), .ZN(new_n495));
  AND2_X1   g070(.A1(KEYINPUT68), .A2(G114), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT68), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT69), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT69), .A2(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n513), .A2(G543), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n511), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT69), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT69), .A2(G651), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n519), .A2(new_n520), .A3(new_n514), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n515), .B1(new_n503), .B2(new_n504), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n513), .A2(new_n526), .A3(KEYINPUT70), .A4(new_n515), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n517), .B1(G88), .B2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n533), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n526), .A2(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n516), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n528), .B2(G89), .ZN(G168));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(new_n524), .B2(new_n525), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT71), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n544), .B(new_n541), .C1(new_n505), .C2(new_n539), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n510), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT72), .A4(new_n510), .ZN(new_n549));
  INV_X1    g124(.A(new_n516), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n523), .A2(G90), .A3(new_n527), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(new_n524), .B2(new_n525), .ZN(new_n556));
  AND2_X1   g131(.A1(G68), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n510), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n513), .A2(G43), .A3(G543), .A4(new_n515), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n523), .A2(G81), .A3(new_n527), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n523), .A2(G91), .A3(new_n527), .ZN(new_n571));
  AND2_X1   g146(.A1(G53), .A2(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n513), .A2(new_n515), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n526), .A2(G65), .ZN(new_n577));
  AND2_X1   g152(.A1(G78), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n571), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n573), .A2(new_n574), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n515), .A4(new_n572), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(KEYINPUT9), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n570), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n571), .A2(new_n576), .A3(new_n579), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n581), .A2(KEYINPUT9), .A3(new_n582), .ZN(new_n586));
  NOR3_X1   g161(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT75), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(G299));
  NAND2_X1  g163(.A1(new_n523), .A2(new_n527), .ZN(new_n589));
  INV_X1    g164(.A(G89), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n535), .B1(new_n536), .B2(new_n516), .C1(new_n589), .C2(new_n590), .ZN(G286));
  INV_X1    g166(.A(G88), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n511), .B1(new_n512), .B2(new_n516), .C1(new_n589), .C2(new_n592), .ZN(G303));
  NAND2_X1  g168(.A1(new_n528), .A2(G87), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n526), .A2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n550), .A2(G49), .B1(new_n595), .B2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n510), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G48), .B2(new_n550), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n528), .A2(G86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(new_n528), .A2(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n505), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n550), .A2(G47), .B1(new_n607), .B2(new_n510), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n604), .A2(KEYINPUT76), .A3(new_n608), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT77), .B(KEYINPUT10), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n589), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n589), .B2(new_n615), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n505), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n550), .A2(G54), .B1(new_n621), .B2(G651), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n614), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n614), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n464), .A2(new_n474), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n470), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n485), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n465), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n642), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT78), .B(KEYINPUT14), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT80), .Z(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT81), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n670), .B2(new_n671), .ZN(new_n675));
  INV_X1    g250(.A(new_n671), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n676), .A2(new_n672), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n673), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G6), .A2(G16), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n601), .A2(new_n602), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(G16), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT32), .ZN(new_n703));
  INV_X1    g278(.A(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1971), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n706), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT33), .B(G1976), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n709), .B2(new_n710), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n705), .A2(new_n711), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  MUX2_X1   g294(.A(G24), .B(G290), .S(G16), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT85), .B(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G29), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G25), .ZN(new_n724));
  AOI22_X1  g299(.A1(G119), .A2(new_n485), .B1(new_n470), .B2(G131), .ZN(new_n725));
  OR2_X1    g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n727), .A2(KEYINPUT82), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(KEYINPUT82), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT83), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n724), .B1(new_n731), .B2(new_n723), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT84), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n732), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n722), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n719), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n705), .A2(new_n711), .A3(new_n718), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT34), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT87), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT87), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n741), .A3(KEYINPUT34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n737), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT88), .B(KEYINPUT36), .Z(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(G299), .A2(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n706), .A2(G20), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT23), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G1956), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n723), .A2(G35), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G162), .B2(new_n723), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n756), .B(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT25), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n464), .A2(G127), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n465), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n764), .B(new_n767), .C1(G139), .C2(new_n470), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n723), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n723), .B2(G33), .ZN(new_n770));
  INV_X1    g345(.A(G2072), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT30), .B(G28), .ZN(new_n773));
  OR2_X1    g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  NAND2_X1  g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n723), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n772), .B(new_n776), .C1(new_n723), .C2(new_n647), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n706), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n706), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(G1966), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n781), .A2(KEYINPUT93), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT26), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G129), .B2(new_n485), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(new_n723), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n723), .A2(G32), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OR3_X1    g367(.A1(new_n790), .A2(new_n791), .A3(new_n784), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n792), .B(new_n793), .C1(new_n770), .C2(new_n771), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n777), .A2(new_n782), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(KEYINPUT93), .B2(new_n781), .ZN(new_n796));
  NOR2_X1   g371(.A1(G27), .A2(G29), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G164), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  INV_X1    g374(.A(G2084), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n723), .B1(KEYINPUT24), .B2(G34), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(KEYINPUT24), .B2(G34), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n482), .B2(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n799), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G171), .A2(new_n706), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G5), .B2(new_n706), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n759), .A2(new_n754), .B1(G1966), .B2(new_n779), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n804), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n803), .A2(new_n800), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n807), .B2(new_n806), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n796), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n760), .A2(new_n761), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n624), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G4), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1348), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n470), .A2(G140), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n485), .A2(G128), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n465), .A2(G116), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n723), .A2(G26), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT28), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT90), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2067), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n817), .A2(new_n818), .ZN(new_n831));
  NOR2_X1   g406(.A1(G16), .A2(G19), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n563), .B2(G16), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT89), .B(G1341), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n819), .A2(new_n830), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT91), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n762), .A2(new_n814), .A3(new_n815), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n746), .A2(new_n747), .A3(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  NAND2_X1  g415(.A1(new_n624), .A2(G559), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT38), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n524), .B2(new_n525), .ZN(new_n844));
  AND2_X1   g419(.A1(G80), .A2(G543), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n510), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(KEYINPUT97), .A2(G55), .ZN(new_n847));
  NOR2_X1   g422(.A1(KEYINPUT97), .A2(G55), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n513), .A2(new_n849), .A3(G543), .A4(new_n515), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n523), .A2(G93), .A3(new_n527), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n561), .A2(new_n560), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n561), .A2(new_n560), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n842), .B(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n857), .A2(new_n858), .A3(G860), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(new_n852), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n859), .A2(new_n862), .ZN(G145));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n470), .A2(G142), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT98), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n485), .A2(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n465), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT99), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n638), .ZN(new_n872));
  INV_X1    g447(.A(new_n731), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n871), .A2(new_n638), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n638), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n731), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(KEYINPUT100), .A3(new_n877), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n500), .B(new_n824), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n789), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(new_n768), .Z(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n482), .B(new_n647), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n489), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n881), .A2(new_n884), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n885), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n864), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n894), .A2(KEYINPUT40), .A3(new_n890), .A4(new_n889), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n893), .A2(new_n895), .ZN(G395));
  NAND2_X1  g471(.A1(new_n860), .A2(new_n627), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n584), .B2(new_n587), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n580), .A2(new_n570), .A3(new_n583), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT75), .B1(new_n585), .B2(new_n586), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n624), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(G299), .A2(new_n900), .A3(new_n623), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n633), .B(new_n855), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n912), .B2(new_n907), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n714), .A2(G303), .ZN(new_n914));
  NAND2_X1  g489(.A1(G288), .A2(G166), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n612), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT76), .B1(new_n604), .B2(new_n608), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n917), .A2(new_n701), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G305), .B1(new_n611), .B2(new_n612), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n701), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n611), .A2(G305), .A3(new_n612), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n915), .A4(new_n914), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n925), .A2(KEYINPUT102), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n913), .B(new_n932), .Z(new_n933));
  OAI21_X1  g508(.A(new_n897), .B1(new_n933), .B2(new_n627), .ZN(G331));
  XNOR2_X1  g509(.A(G331), .B(KEYINPUT103), .ZN(G295));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g511(.A1(G301), .A2(G286), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n552), .A2(new_n551), .ZN(new_n938));
  NAND4_X1  g513(.A1(G168), .A2(new_n938), .A3(new_n549), .A4(new_n548), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n855), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n853), .ZN(new_n941));
  INV_X1    g516(.A(new_n854), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n937), .A2(new_n939), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n936), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n936), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n949), .A2(new_n910), .A3(new_n911), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n946), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n855), .A2(new_n937), .A3(new_n939), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n903), .A2(new_n904), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n953), .A2(new_n925), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n890), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT106), .B1(new_n949), .B2(new_n905), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n951), .A2(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n910), .A2(new_n911), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n906), .A2(new_n964), .A3(new_n948), .A4(new_n944), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n926), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n950), .A2(new_n953), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n926), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n959), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n959), .A2(new_n974), .A3(new_n969), .A4(new_n971), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n968), .A2(new_n973), .A3(KEYINPUT44), .A4(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n950), .A2(new_n957), .A3(new_n954), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n957), .B1(new_n950), .B2(new_n954), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n953), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT41), .B1(new_n903), .B2(new_n904), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(new_n949), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n890), .B1(new_n984), .B2(new_n925), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT43), .B1(new_n966), .B2(new_n926), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n959), .A2(new_n987), .A3(new_n890), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT107), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n992), .B(KEYINPUT44), .C1(new_n986), .C2(new_n988), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n976), .B1(new_n991), .B2(new_n993), .ZN(G397));
  XOR2_X1   g569(.A(KEYINPUT109), .B(G40), .Z(new_n995));
  NAND4_X1  g570(.A1(new_n473), .A2(new_n481), .A3(new_n475), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n500), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2067), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n824), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT110), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(new_n789), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1000), .A2(G1996), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1004), .A2(new_n1006), .B1(new_n789), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1000), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n873), .A2(new_n734), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n873), .A2(new_n734), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT125), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n500), .A2(new_n998), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n996), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  OAI21_X1  g594(.A(G1981), .B1(new_n600), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n701), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1020), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G305), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G305), .B(new_n1020), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT112), .B1(new_n1027), .B2(KEYINPUT49), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1021), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1026), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1034), .A2(new_n999), .A3(new_n996), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n500), .A2(new_n1037), .A3(new_n998), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n997), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n1035), .A2(G1971), .B1(new_n1039), .B2(G2090), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT55), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1043), .A3(G8), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1018), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1045), .B(new_n1047), .C1(new_n1046), .C2(G288), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G288), .A2(new_n1046), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n1018), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1032), .A2(new_n1044), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1036), .A2(new_n1053), .A3(new_n997), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1037), .B1(new_n500), .B2(new_n998), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT113), .B1(new_n1055), .B2(new_n996), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1056), .A3(new_n1038), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1057), .A2(G2090), .B1(G1971), .B2(new_n1035), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1043), .B1(new_n1058), .B2(G8), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1016), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(G8), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1042), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1027), .A2(KEYINPUT112), .A3(KEYINPUT49), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1066), .B2(new_n1026), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1067), .A3(KEYINPUT125), .A4(new_n1044), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1060), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1034), .A2(new_n999), .ZN(new_n1070));
  INV_X1    g645(.A(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n481), .A2(KEYINPUT53), .A3(G40), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n476), .B2(KEYINPUT123), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1070), .B(new_n1073), .C1(KEYINPUT123), .C2(new_n476), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT45), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1017), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n997), .A3(new_n1033), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1078), .B2(G2078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1039), .A2(new_n807), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1074), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1035), .A2(KEYINPUT53), .A3(new_n1071), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1082), .B(KEYINPUT54), .C1(G171), .C2(new_n1084), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT114), .B(G2084), .Z(new_n1086));
  NAND4_X1  g661(.A1(new_n1036), .A2(new_n997), .A3(new_n1038), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1035), .B2(G1966), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(G286), .ZN(new_n1089));
  OAI211_X1 g664(.A(G168), .B(new_n1087), .C1(new_n1035), .C2(G1966), .ZN(new_n1090));
  INV_X1    g665(.A(G8), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT121), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1090), .A2(KEYINPUT51), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1085), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1084), .A2(G171), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1074), .A2(new_n1079), .A3(G301), .A4(new_n1080), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT124), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1096), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(KEYINPUT124), .A3(new_n1100), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1069), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1057), .A2(new_n752), .B1(new_n1035), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n585), .A2(new_n586), .B1(KEYINPUT116), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT117), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n996), .A2(new_n1017), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1039), .A2(new_n818), .B1(new_n1001), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n623), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1111), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1112), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT119), .B(new_n1121), .C1(new_n1122), .C2(new_n1112), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1111), .A2(KEYINPUT61), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1077), .A2(new_n997), .A3(new_n1005), .A4(new_n1033), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1117), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  AOI22_X1  g708(.A1(new_n1130), .A2(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1035), .A2(KEYINPUT118), .A3(new_n1005), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n562), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT59), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1118), .A2(new_n623), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT60), .B1(new_n1138), .B2(new_n1119), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1118), .A2(new_n1140), .A3(new_n624), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1128), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1115), .A4(new_n1113), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1127), .A2(new_n1129), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1104), .B1(new_n1120), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1088), .A2(G8), .A3(G168), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1052), .A2(new_n1059), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT115), .B1(new_n1150), .B2(KEYINPUT63), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1067), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1044), .A2(KEYINPUT63), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1043), .B1(new_n1040), .B2(G8), .ZN(new_n1154));
  OR4_X1    g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1149), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT115), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1062), .A2(new_n1067), .A3(new_n1044), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1156), .B(new_n1157), .C1(new_n1158), .C2(new_n1149), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1095), .A2(KEYINPUT62), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1097), .B1(new_n1095), .B2(KEYINPUT62), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1069), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1032), .A2(new_n1046), .A3(new_n714), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(G1981), .B2(G305), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1044), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1165), .A2(new_n1045), .B1(new_n1166), .B2(new_n1067), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1160), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1015), .B1(new_n1148), .B2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(G290), .A2(new_n1000), .A3(G1986), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1013), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1008), .A2(KEYINPUT126), .A3(new_n1012), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n824), .A2(G2067), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1000), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1007), .B(KEYINPUT46), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1179), .A2(new_n1004), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT47), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1175), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1169), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g758(.A1(new_n894), .A2(new_n890), .A3(new_n889), .ZN(new_n1185));
  NOR4_X1   g759(.A1(G401), .A2(G229), .A3(new_n460), .A4(G227), .ZN(new_n1186));
  NAND3_X1  g760(.A1(new_n1185), .A2(new_n989), .A3(new_n1186), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


