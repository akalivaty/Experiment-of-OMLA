//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n202), .B2(new_n203), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(G50gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT89), .B(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n207), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n215), .B2(KEYINPUT90), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(KEYINPUT90), .B2(new_n215), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n210), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT91), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT91), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n211), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n205), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT92), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT92), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(new_n225), .A3(new_n205), .A4(new_n222), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n213), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G15gat), .B(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(G1gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(G1gat), .B2(new_n230), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n227), .A2(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G229gat), .A2(G233gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n237), .B1(new_n229), .B2(new_n235), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n239), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n227), .A2(new_n235), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n237), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n239), .B(KEYINPUT13), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n242), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT11), .B(G169gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G197gat), .ZN(new_n251));
  XOR2_X1   g050(.A(G113gat), .B(G141gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n242), .A2(new_n244), .A3(new_n248), .A4(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  INV_X1    g059(.A(G85gat), .ZN(new_n261));
  INV_X1    g060(.A(G92gat), .ZN(new_n262));
  AOI22_X1  g061(.A1(KEYINPUT8), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT97), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G85gat), .A2(G92gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT7), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G99gat), .B(G106gat), .Z(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n269), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n271), .A3(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G64gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(G57gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(G57gat), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(KEYINPUT94), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(KEYINPUT94), .B2(new_n276), .ZN(new_n278));
  XOR2_X1   g077(.A(G71gat), .B(G78gat), .Z(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT93), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n276), .B2(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n279), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n273), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n270), .A2(new_n285), .A3(new_n283), .A4(new_n272), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT99), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT99), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(new_n288), .A3(new_n293), .A4(new_n289), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G230gat), .A2(G233gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G120gat), .B(G148gat), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(G204gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(new_n274), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(new_n262), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(KEYINPUT22), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n328), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT66), .B1(new_n333), .B2(G183gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT65), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G190gat), .ZN(new_n336));
  INV_X1    g135(.A(G190gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT65), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT27), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(G183gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT66), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n332), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(KEYINPUT65), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n335), .A2(G190gat), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(new_n346), .B1(new_n341), .B2(KEYINPUT66), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT66), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n333), .A2(G183gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n340), .A2(KEYINPUT27), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n351), .A3(KEYINPUT67), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n344), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n349), .A2(new_n350), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n345), .A2(new_n346), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT28), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n331), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n327), .B(KEYINPUT23), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n324), .B(KEYINPUT64), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n340), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n330), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n362), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n365), .B(new_n366), .C1(G183gat), .C2(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n359), .A2(new_n324), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n361), .A2(new_n368), .B1(new_n370), .B2(new_n362), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n323), .B1(new_n358), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n357), .ZN(new_n374));
  INV_X1    g173(.A(new_n331), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n368), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n362), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n373), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n321), .B(new_n372), .C1(new_n380), .C2(new_n323), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n358), .A2(new_n371), .ZN(new_n382));
  OAI211_X1 g181(.A(KEYINPUT72), .B(new_n322), .C1(new_n382), .C2(new_n373), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n320), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n322), .B1(new_n382), .B2(KEYINPUT29), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n319), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT30), .B(new_n312), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n384), .A2(new_n386), .A3(new_n312), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(KEYINPUT73), .ZN(new_n389));
  AND2_X1   g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G141gat), .B(G148gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(G155gat), .B2(G162gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G141gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G148gat), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G155gat), .B(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT2), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT3), .ZN(new_n407));
  INV_X1    g206(.A(G134gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(G127gat), .ZN(new_n409));
  INV_X1    g208(.A(G127gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(G134gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G113gat), .B(G120gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(KEYINPUT1), .ZN(new_n414));
  INV_X1    g213(.A(G120gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G113gat), .ZN(new_n416));
  INV_X1    g215(.A(G113gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G120gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n424));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n405), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G225gat), .A2(G233gat), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n414), .A2(new_n396), .A3(new_n422), .A4(new_n405), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT68), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n419), .A2(new_n421), .B1(new_n409), .B2(new_n411), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n422), .A3(KEYINPUT68), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n396), .A2(new_n405), .A3(KEYINPUT75), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT75), .B1(new_n396), .B2(new_n405), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n435), .B(new_n436), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n426), .B(new_n431), .C1(new_n439), .C2(new_n430), .ZN(new_n440));
  INV_X1    g239(.A(new_n429), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n422), .A2(new_n414), .B1(new_n396), .B2(new_n405), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n428), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT76), .B1(new_n443), .B2(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n406), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n427), .B1(new_n445), .B2(new_n429), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT76), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n440), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G57gat), .B(G85gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n429), .A2(KEYINPUT4), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT78), .B(new_n456), .C1(new_n439), .C2(KEYINPUT4), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n435), .A2(new_n436), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n406), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n396), .A2(new_n405), .A3(KEYINPUT75), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n459), .A3(new_n430), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n457), .A2(new_n426), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n455), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n455), .B1(new_n450), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT80), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n450), .A2(new_n466), .ZN(new_n474));
  INV_X1    g273(.A(new_n455), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n469), .A4(new_n467), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n473), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n376), .A2(new_n379), .ZN(new_n481));
  INV_X1    g280(.A(new_n373), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n323), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n372), .A2(new_n321), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n383), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n386), .B1(new_n485), .B2(new_n319), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n480), .B1(new_n486), .B2(new_n311), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n319), .ZN(new_n488));
  INV_X1    g287(.A(new_n386), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT73), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT30), .A4(new_n312), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n389), .A2(new_n479), .A3(new_n487), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR4_X1   g294(.A1(new_n486), .A2(KEYINPUT73), .A3(new_n480), .A4(new_n311), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT30), .B1(new_n490), .B2(new_n312), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(KEYINPUT81), .A3(new_n479), .A4(new_n389), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n382), .A2(new_n458), .ZN(new_n500));
  INV_X1    g299(.A(new_n458), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n358), .B2(new_n371), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G227gat), .ZN(new_n504));
  INV_X1    g303(.A(G233gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT33), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(KEYINPUT32), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G43gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G71gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G99gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n506), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n500), .B2(new_n502), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n512), .A2(new_n508), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT69), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522));
  NOR4_X1   g321(.A1(new_n516), .A2(new_n522), .A3(new_n517), .A4(new_n519), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n514), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n503), .A2(new_n506), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT34), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(G22gat), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n406), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(new_n407), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT83), .B(new_n406), .C1(new_n532), .C2(KEYINPUT3), .ZN(new_n536));
  NAND2_X1  g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n425), .A2(new_n482), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n319), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n535), .A2(new_n536), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n424), .B1(new_n319), .B2(new_n373), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(new_n462), .A3(new_n461), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n540), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n537), .B(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G50gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT84), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n547), .A2(new_n549), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n531), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g352(.A1(new_n547), .A2(new_n549), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(new_n530), .A3(new_n550), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n526), .B(new_n514), .C1(new_n521), .C2(new_n523), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n528), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n495), .A2(new_n499), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT35), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n455), .B(KEYINPUT86), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(new_n450), .B2(new_n466), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n470), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n473), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT35), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n556), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n528), .A2(KEYINPUT70), .A3(new_n557), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n524), .A2(new_n527), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT85), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n492), .A2(new_n487), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n311), .B1(new_n488), .B2(new_n489), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n488), .A2(new_n489), .A3(new_n311), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT30), .A2(new_n574), .B1(new_n575), .B2(new_n491), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n572), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n389), .A2(KEYINPUT85), .A3(new_n487), .A4(new_n492), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n495), .A2(new_n499), .ZN(new_n582));
  INV_X1    g381(.A(new_n556), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n457), .A2(new_n426), .A3(new_n464), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n428), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n586), .A2(KEYINPUT39), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n445), .A2(new_n427), .A3(new_n429), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT39), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT87), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n561), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n594), .A2(new_n595), .A3(new_n562), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n578), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT88), .B(KEYINPUT37), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n384), .B2(new_n386), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n385), .A2(new_n319), .A3(new_n372), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT37), .B(new_n601), .C1(new_n485), .C2(new_n319), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n599), .A2(new_n600), .A3(new_n311), .A4(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n574), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n603), .A2(new_n604), .A3(new_n565), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n311), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT38), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n583), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n597), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n528), .B2(new_n557), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n568), .A2(new_n570), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n584), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  AOI211_X1 g414(.A(new_n259), .B(new_n308), .C1(new_n581), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n619));
  XOR2_X1   g418(.A(G134gat), .B(G162gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT41), .ZN(new_n623));
  INV_X1    g422(.A(G232gat), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n623), .A2(new_n624), .A3(new_n505), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n227), .A2(new_n273), .ZN(new_n626));
  AOI211_X1 g425(.A(new_n625), .B(new_n626), .C1(new_n229), .C2(new_n273), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n618), .A2(KEYINPUT98), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n629), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n625), .B1(new_n229), .B2(new_n273), .ZN(new_n632));
  INV_X1    g431(.A(new_n626), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n628), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n622), .B1(new_n630), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n629), .B1(new_n627), .B2(new_n628), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n635), .A3(new_n631), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n621), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT21), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n235), .B1(new_n286), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G183gat), .ZN(new_n644));
  XOR2_X1   g443(.A(G127gat), .B(G155gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT95), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT96), .B(G211gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n646), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n286), .A2(new_n642), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n651), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n641), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n616), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n479), .B(KEYINPUT100), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  INV_X1    g461(.A(new_n579), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n665), .A2(new_n667), .B1(KEYINPUT101), .B2(KEYINPUT42), .ZN(new_n668));
  OR2_X1    g467(.A1(KEYINPUT101), .A2(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n658), .A2(KEYINPUT42), .A3(new_n663), .A4(new_n667), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n670), .B(new_n671), .C1(new_n234), .C2(new_n665), .ZN(G1325gat));
  AOI21_X1  g471(.A(G15gat), .B1(new_n658), .B2(new_n613), .ZN(new_n673));
  INV_X1    g472(.A(new_n614), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n658), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n673), .B1(new_n675), .B2(G15gat), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n583), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  AOI21_X1  g478(.A(new_n641), .B1(new_n581), .B2(new_n615), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n259), .A2(new_n655), .A3(new_n308), .ZN(new_n681));
  AND2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n202), .A3(new_n660), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n681), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G29gat), .B1(new_n687), .B2(new_n659), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n682), .A2(new_n203), .A3(new_n663), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  OAI21_X1  g490(.A(G36gat), .B1(new_n687), .B2(new_n579), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1329gat));
  OAI21_X1  g492(.A(G43gat), .B1(new_n687), .B2(new_n614), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n682), .A2(new_n207), .A3(new_n613), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT47), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n696), .B(new_n698), .ZN(G1330gat));
  AND2_X1   g498(.A1(new_n682), .A2(new_n583), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n583), .A2(new_n214), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n700), .A2(new_n214), .B1(new_n687), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g502(.A(new_n308), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n656), .A2(new_n258), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT104), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n581), .A2(new_n615), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n659), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT105), .B(G57gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n579), .ZN(new_n712));
  NOR2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  AND2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n712), .B2(new_n713), .ZN(G1333gat));
  OAI21_X1  g515(.A(G71gat), .B1(new_n708), .B2(new_n614), .ZN(new_n717));
  INV_X1    g516(.A(new_n708), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n613), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n719), .B2(G71gat), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n583), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n258), .A2(new_n655), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n685), .A2(new_n308), .A3(new_n686), .A4(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n659), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT106), .Z(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n724), .B1(new_n680), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  AOI211_X1 g529(.A(KEYINPUT107), .B(new_n641), .C1(new_n581), .C2(new_n615), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n308), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n660), .A2(new_n261), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n727), .A2(new_n261), .B1(new_n737), .B2(new_n738), .ZN(G1336gat));
  NOR2_X1   g538(.A1(new_n579), .A2(G92gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n704), .B(new_n741), .C1(new_n733), .C2(new_n734), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n579), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n262), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT52), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n737), .B2(new_n741), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(new_n744), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n725), .B2(new_n614), .ZN(new_n749));
  INV_X1    g548(.A(G99gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n735), .A2(new_n750), .A3(new_n308), .A4(new_n736), .ZN(new_n751));
  INV_X1    g550(.A(new_n613), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT109), .B(new_n749), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1338gat));
  NOR3_X1   g556(.A1(new_n704), .A2(G106gat), .A3(new_n556), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n735), .A2(new_n736), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  OAI21_X1  g559(.A(G106gat), .B1(new_n725), .B2(new_n556), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n724), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n637), .A2(new_n640), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n584), .A2(new_n610), .A3(new_n614), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n559), .A2(KEYINPUT35), .B1(new_n571), .B2(new_n579), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n767), .B2(KEYINPUT107), .ZN(new_n768));
  INV_X1    g567(.A(new_n731), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT51), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n758), .B1(new_n770), .B2(new_n732), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n773), .B(new_n758), .C1(new_n770), .C2(new_n732), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n761), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(KEYINPUT53), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n762), .B1(new_n777), .B2(new_n778), .ZN(G1339gat));
  NOR3_X1   g578(.A1(new_n656), .A2(new_n258), .A3(new_n308), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n295), .A2(new_n781), .A3(new_n296), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n305), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n291), .A2(new_n299), .A3(new_n292), .A4(new_n294), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n297), .A2(KEYINPUT54), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(KEYINPUT55), .A3(new_n785), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n306), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n243), .A2(new_n239), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n246), .A2(new_n247), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n253), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n257), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n764), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n257), .A2(new_n308), .A3(new_n794), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n797), .B1(new_n791), .B2(new_n258), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n798), .B2(new_n764), .ZN(new_n799));
  INV_X1    g598(.A(new_n655), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n780), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n558), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n660), .A2(new_n579), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n417), .A3(new_n258), .ZN(new_n805));
  INV_X1    g604(.A(new_n780), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n257), .A2(new_n794), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n641), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n797), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n259), .B2(new_n807), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n809), .B1(new_n811), .B2(new_n641), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n806), .B1(new_n812), .B2(new_n655), .ZN(new_n813));
  INV_X1    g612(.A(new_n803), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n752), .A2(new_n583), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n816), .A2(new_n258), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n805), .B1(new_n817), .B2(new_n417), .ZN(G1340gat));
  NAND3_X1  g617(.A1(new_n804), .A2(new_n415), .A3(new_n308), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n816), .A2(new_n308), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n415), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n804), .B2(new_n655), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n800), .A2(new_n410), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n816), .B2(new_n823), .ZN(G1342gat));
  AOI21_X1  g623(.A(new_n408), .B1(new_n816), .B2(new_n764), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n813), .A2(new_n764), .A3(new_n558), .A4(new_n814), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT113), .B1(new_n826), .B2(G134gat), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n804), .A2(new_n828), .A3(new_n408), .A4(new_n764), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n825), .B1(new_n830), .B2(KEYINPUT56), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n827), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n827), .A2(new_n829), .A3(KEYINPUT114), .A4(new_n832), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n831), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n831), .A2(new_n835), .A3(KEYINPUT115), .A4(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1343gat));
  NAND2_X1  g640(.A1(new_n783), .A2(new_n785), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n788), .A3(new_n306), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n256), .A2(new_n257), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n789), .A2(KEYINPUT116), .A3(new_n844), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n797), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n796), .B1(new_n849), .B2(new_n764), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n780), .B1(new_n850), .B2(new_n800), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT57), .B1(new_n851), .B2(new_n556), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n813), .A2(new_n853), .A3(new_n583), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n674), .A2(new_n803), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n854), .A3(new_n258), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G141gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n258), .A2(new_n397), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT117), .ZN(new_n859));
  AND4_X1   g658(.A1(new_n583), .A2(new_n813), .A3(new_n855), .A4(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(KEYINPUT118), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n857), .B2(new_n861), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT118), .B(new_n860), .C1(new_n856), .C2(G141gat), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n866), .A2(new_n870), .ZN(G1344gat));
  NOR2_X1   g670(.A1(new_n801), .A2(new_n556), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n872), .A2(new_n855), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n399), .A3(new_n308), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n846), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n258), .A2(new_n876), .A3(new_n848), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n764), .B1(new_n877), .B2(new_n810), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n800), .B1(new_n878), .B2(new_n809), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n806), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n583), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n801), .A2(new_n853), .A3(new_n556), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT119), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n308), .A3(new_n855), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n875), .B1(new_n888), .B2(G148gat), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n852), .A2(new_n855), .ZN(new_n890));
  INV_X1    g689(.A(new_n854), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n399), .C1(new_n892), .C2(new_n308), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n874), .B1(new_n889), .B2(new_n893), .ZN(G1345gat));
  AOI21_X1  g693(.A(G155gat), .B1(new_n873), .B2(new_n655), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n890), .A2(new_n891), .A3(new_n800), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g696(.A(G162gat), .B1(new_n873), .B2(new_n764), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n892), .A2(G162gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n764), .ZN(G1347gat));
  NOR2_X1   g699(.A1(new_n660), .A2(new_n579), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n801), .A2(new_n802), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n904), .A3(new_n258), .ZN(new_n905));
  XOR2_X1   g704(.A(new_n905), .B(KEYINPUT120), .Z(new_n906));
  NOR2_X1   g705(.A1(new_n801), .A2(new_n902), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n815), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT121), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n907), .A2(new_n910), .A3(new_n815), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n259), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n906), .A2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n903), .B2(new_n308), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n704), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(G176gat), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n903), .A2(new_n655), .A3(new_n355), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n912), .A2(new_n800), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n340), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT60), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT60), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n922), .B(new_n918), .C1(new_n919), .C2(new_n340), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n764), .A3(new_n356), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n764), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n928), .B2(G190gat), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT61), .B(new_n337), .C1(new_n927), .C2(new_n764), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n902), .A2(new_n674), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n887), .A2(new_n258), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT123), .B(G197gat), .Z(new_n935));
  INV_X1    g734(.A(new_n932), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n883), .B2(new_n886), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n258), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n934), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n614), .A2(new_n663), .A3(new_n583), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT122), .ZN(new_n943));
  NOR4_X1   g742(.A1(new_n801), .A2(new_n660), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n935), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n258), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n940), .A2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n887), .A2(new_n308), .A3(new_n932), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n937), .A2(new_n950), .A3(new_n308), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n949), .A2(G204gat), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n944), .A2(new_n304), .A3(new_n308), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT62), .Z(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n314), .A3(new_n655), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n887), .A2(new_n655), .A3(new_n932), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n957), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT63), .B1(new_n957), .B2(G211gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n315), .B1(new_n937), .B2(new_n764), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n315), .A3(new_n764), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n641), .B(new_n936), .C1(new_n883), .C2(new_n886), .ZN(new_n966));
  OAI211_X1 g765(.A(KEYINPUT126), .B(new_n963), .C1(new_n966), .C2(new_n315), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1355gat));
endmodule


