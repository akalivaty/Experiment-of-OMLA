//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G104), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n187), .A2(G107), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT4), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(new_n191), .A3(new_n193), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT75), .A2(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(new_n198), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n202), .B(new_n203), .C1(new_n205), .C2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n212), .A2(new_n202), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(new_n214), .A3(new_n202), .A4(new_n203), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n190), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n187), .A2(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  AND4_X1   g039(.A1(new_n225), .A2(new_n210), .A3(new_n211), .A4(G128), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n194), .B(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n201), .A2(new_n217), .B1(new_n218), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n231), .A2(new_n234), .A3(new_n237), .A4(new_n232), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n194), .A2(new_n221), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT76), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n194), .A2(new_n221), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n222), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n210), .A2(KEYINPUT65), .A3(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G128), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n226), .B1(new_n248), .B2(new_n212), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n244), .A2(new_n250), .A3(KEYINPUT10), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n228), .A2(new_n239), .A3(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G140), .ZN(new_n253));
  INV_X1    g067(.A(G227), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(G953), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n253), .B(new_n255), .Z(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT81), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n241), .A3(new_n243), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n227), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n236), .A2(new_n238), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(KEYINPUT12), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n260), .A2(KEYINPUT77), .A3(KEYINPUT12), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n239), .B1(new_n260), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(KEYINPUT78), .A3(new_n227), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n252), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n244), .A2(new_n250), .A3(KEYINPUT10), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n226), .B1(new_n212), .B2(new_n223), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n218), .B1(new_n275), .B2(new_n240), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n196), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n277), .B1(new_n198), .B2(new_n195), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n278), .B2(new_n216), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n261), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT80), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n201), .A2(new_n217), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n251), .A3(new_n276), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n261), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n273), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n286), .A2(KEYINPUT82), .A3(new_n256), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT82), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n281), .B(new_n239), .C1(new_n228), .C2(new_n251), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT80), .B1(new_n284), .B2(new_n261), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n252), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n256), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n272), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G469), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n252), .B1(new_n266), .B2(new_n270), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT79), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT79), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n300), .B(new_n252), .C1(new_n266), .C2(new_n270), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n292), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n256), .B(new_n252), .C1(new_n289), .C2(new_n290), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(G469), .A3(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n295), .A2(new_n296), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT9), .B(G234), .Z(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n296), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(G221), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT74), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n314), .B2(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n313), .A3(KEYINPUT72), .A4(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT71), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G140), .ZN(new_n322));
  AND4_X1   g136(.A1(KEYINPUT71), .A2(new_n314), .A3(new_n322), .A4(KEYINPUT16), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n318), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n206), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n314), .A2(new_n322), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n316), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n319), .A2(KEYINPUT71), .A3(KEYINPUT16), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(G146), .A3(new_n318), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G214), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT86), .A3(G143), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT86), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n204), .ZN(new_n337));
  NOR2_X1   g151(.A1(G237), .A2(G953), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT86), .A2(G143), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n337), .A2(G214), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT17), .A3(G131), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n325), .A2(new_n331), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT88), .B1(new_n341), .B2(new_n237), .ZN(new_n348));
  AOI21_X1  g162(.A(G131), .B1(new_n335), .B2(new_n340), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n342), .A2(KEYINPUT88), .A3(G131), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n325), .A2(new_n331), .A3(new_n343), .A4(KEYINPUT89), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n187), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n342), .A2(KEYINPUT18), .A3(G131), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n327), .A2(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n319), .A2(new_n206), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT87), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT18), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n341), .B1(new_n361), .B2(new_n237), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n319), .A2(KEYINPUT87), .A3(new_n206), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n357), .A2(new_n360), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n354), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n356), .B1(new_n354), .B2(new_n364), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n296), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT91), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n296), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT90), .B(G475), .Z(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n354), .A2(new_n356), .A3(new_n364), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n350), .A2(new_n351), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n319), .B(KEYINPUT19), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n206), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n331), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n364), .ZN(new_n379));
  INV_X1    g193(.A(new_n356), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n373), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G475), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n296), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT20), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT20), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(new_n386), .A3(new_n383), .A4(new_n296), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n372), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G128), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(G143), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(KEYINPUT13), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT92), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n392), .A2(KEYINPUT13), .ZN(new_n395));
  OAI21_X1  g209(.A(G134), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n391), .A3(new_n230), .ZN(new_n398));
  XNOR2_X1  g212(.A(G116), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n190), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n399), .ZN(new_n402));
  INV_X1    g216(.A(G116), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n403), .B2(G122), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(G107), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n399), .B1(KEYINPUT14), .B2(new_n190), .ZN(new_n406));
  INV_X1    g220(.A(new_n398), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n230), .B1(new_n397), .B2(new_n391), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n308), .A2(G217), .A3(new_n333), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT93), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n410), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n413), .A2(new_n296), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n413), .B2(new_n296), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n389), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n307), .A2(new_n311), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT67), .A3(G116), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT67), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(new_n403), .B2(G119), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n403), .A2(G119), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(KEYINPUT2), .A2(G113), .ZN(new_n429));
  NOR2_X1   g243(.A1(KEYINPUT2), .A2(G113), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(KEYINPUT66), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n428), .B2(KEYINPUT66), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n261), .A2(new_n213), .A3(new_n209), .A4(new_n215), .ZN(new_n437));
  INV_X1    g251(.A(new_n232), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n230), .A2(G137), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n205), .A2(new_n207), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n390), .B1(new_n222), .B2(new_n245), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n247), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n238), .B(new_n440), .C1(new_n443), .C2(new_n226), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n437), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n436), .B1(new_n437), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT28), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT70), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n440), .A2(new_n238), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n216), .A2(new_n239), .B1(new_n249), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n435), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n433), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n450), .B1(new_n455), .B2(new_n445), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n445), .A2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n459), .B2(KEYINPUT70), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n338), .A2(G210), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G101), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT29), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n296), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n437), .A2(new_n444), .A3(KEYINPUT30), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(new_n454), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(new_n445), .ZN(new_n472));
  INV_X1    g286(.A(new_n465), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n465), .B1(new_n456), .B2(new_n458), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT29), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G472), .B1(new_n467), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT32), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n465), .B1(new_n448), .B2(new_n457), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n445), .A3(new_n465), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT31), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n471), .A2(KEYINPUT31), .A3(new_n445), .A4(new_n465), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT69), .Z(new_n486));
  OAI21_X1  g300(.A(new_n478), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(new_n483), .ZN(new_n488));
  INV_X1    g302(.A(new_n479), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n486), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT32), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n477), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT22), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(G137), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n423), .A2(G128), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(KEYINPUT23), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(KEYINPUT23), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n499), .B(new_n500), .C1(G119), .C2(new_n390), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G110), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  XNOR2_X1  g317(.A(G119), .B(G128), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n324), .A2(new_n206), .ZN(new_n506));
  AOI21_X1  g320(.A(G146), .B1(new_n330), .B2(new_n318), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n502), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT73), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n501), .A2(G110), .B1(new_n504), .B2(new_n503), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n331), .A3(new_n359), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n497), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n511), .A3(new_n496), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n296), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G217), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n521), .B1(G234), .B2(new_n296), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n514), .A2(new_n515), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n493), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n321), .B1(new_n443), .B2(new_n226), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n321), .B2(new_n216), .ZN(new_n529));
  INV_X1    g343(.A(G224), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(G953), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n529), .B(new_n531), .Z(new_n532));
  OR2_X1    g346(.A1(new_n428), .A2(new_n432), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n427), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(G113), .B(new_n535), .C1(new_n428), .C2(new_n534), .ZN(new_n536));
  INV_X1    g350(.A(new_n243), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n242), .B1(new_n194), .B2(new_n221), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n533), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n436), .B2(new_n278), .ZN(new_n540));
  XOR2_X1   g354(.A(G110), .B(G122), .Z(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n539), .B(new_n543), .C1(new_n436), .C2(new_n278), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n546), .A3(new_n541), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n532), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n536), .A2(new_n533), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n240), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT83), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT83), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n552), .A3(new_n240), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n539), .A3(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n541), .B(KEYINPUT8), .Z(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n557));
  OAI221_X1 g371(.A(new_n528), .B1(new_n557), .B2(new_n531), .C1(new_n321), .C2(new_n216), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n529), .B(KEYINPUT7), .C1(new_n530), .C2(G953), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n544), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n548), .A2(new_n560), .A3(new_n296), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT84), .Z(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT85), .ZN(new_n565));
  INV_X1    g379(.A(new_n563), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n548), .A2(new_n560), .A3(new_n296), .A4(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n567), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G214), .B1(G237), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(G234), .A2(G237), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(G952), .A3(new_n333), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT21), .B(G898), .Z(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(G902), .A3(G953), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n570), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n422), .A2(new_n527), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G101), .ZN(G3));
  NAND2_X1  g395(.A1(new_n523), .A2(new_n526), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G472), .B1(new_n484), .B2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n490), .A2(new_n491), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n307), .A2(new_n583), .A3(new_n311), .A4(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n413), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n414), .B1(new_n588), .B2(G902), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT94), .B1(new_n410), .B2(new_n412), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(new_n413), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n296), .A2(G478), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n572), .B1(new_n564), .B2(new_n567), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n389), .A3(new_n577), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n587), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT34), .B(G104), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  INV_X1    g414(.A(new_n389), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(new_n577), .A3(new_n420), .A4(new_n596), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n587), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NOR2_X1   g419(.A1(new_n512), .A2(new_n513), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n497), .A2(KEYINPUT36), .ZN(new_n607));
  OR2_X1    g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n608), .A2(new_n525), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n523), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n522), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n518), .B2(new_n519), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT95), .B1(new_n615), .B2(new_n610), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n422), .A2(new_n579), .A3(new_n586), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT37), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G110), .ZN(G12));
  INV_X1    g435(.A(new_n311), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT82), .B1(new_n286), .B2(new_n256), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n291), .A2(new_n288), .A3(new_n292), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n272), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n305), .B1(new_n626), .B2(new_n295), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n622), .B1(new_n627), .B2(new_n304), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n613), .A2(new_n493), .A3(new_n616), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n576), .A2(G900), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n574), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n389), .A2(new_n419), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n628), .A2(new_n596), .A3(new_n629), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  XNOR2_X1  g449(.A(new_n631), .B(KEYINPUT97), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT39), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n628), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n570), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n472), .A2(new_n473), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n455), .A2(new_n473), .A3(new_n445), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n296), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n492), .A2(new_n487), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n492), .A2(new_n487), .A3(new_n645), .A4(KEYINPUT96), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n419), .B1(new_n372), .B2(new_n388), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n641), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n618), .A2(new_n572), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n628), .A2(new_n654), .A3(new_n637), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n639), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT98), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G143), .ZN(G45));
  NAND3_X1  g472(.A1(new_n595), .A2(new_n389), .A3(new_n631), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n628), .A2(new_n596), .A3(new_n629), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  AOI22_X1  g477(.A1(new_n623), .A2(new_n624), .B1(new_n271), .B2(new_n258), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(G902), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n294), .A2(KEYINPUT99), .A3(new_n296), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(G469), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n297), .A2(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n310), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT100), .A4(G469), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n527), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n597), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT41), .B(G113), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G15));
  NOR2_X1   g489(.A1(new_n672), .A2(new_n602), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n403), .ZN(G18));
  NAND4_X1  g491(.A1(new_n669), .A2(new_n670), .A3(new_n596), .A4(new_n671), .ZN(new_n678));
  INV_X1    g492(.A(new_n629), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n421), .A2(new_n577), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n423), .ZN(G21));
  AND3_X1   g496(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n460), .A2(new_n473), .ZN(new_n684));
  INV_X1    g498(.A(new_n488), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n491), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n584), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n583), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n389), .A2(new_n420), .A3(new_n596), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT101), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n651), .A2(new_n691), .A3(new_n596), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n688), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n683), .A2(KEYINPUT102), .A3(new_n693), .A4(new_n577), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n695));
  INV_X1    g509(.A(new_n688), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n691), .A2(new_n389), .A3(new_n420), .A4(new_n596), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n691), .B1(new_n651), .B2(new_n596), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n669), .A2(new_n577), .A3(new_n670), .A4(new_n671), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n694), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  INV_X1    g517(.A(new_n678), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n687), .A2(new_n613), .A3(new_n616), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n659), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NAND2_X1  g522(.A1(new_n304), .A2(KEYINPUT103), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n302), .A2(new_n710), .A3(G469), .A4(new_n303), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n709), .A2(new_n297), .A3(new_n306), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n572), .B(new_n310), .C1(new_n568), .C2(new_n569), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n527), .B(new_n660), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n712), .A2(new_n714), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(KEYINPUT104), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n527), .A4(new_n660), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G131), .ZN(G33));
  OAI211_X1 g540(.A(new_n527), .B(new_n633), .C1(new_n715), .C2(new_n716), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  NAND2_X1  g542(.A1(new_n302), .A2(new_n303), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT46), .A3(new_n306), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(G469), .C1(new_n730), .C2(G902), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n731), .A2(KEYINPUT105), .A3(KEYINPUT46), .A4(new_n306), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n736), .A3(new_n297), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n586), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n601), .A2(new_n595), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(KEYINPUT43), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(new_n740), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n739), .B(new_n618), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n738), .A2(new_n670), .A3(new_n637), .A4(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n570), .A2(new_n571), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n746), .B2(new_n747), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n233), .ZN(G39));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n738), .A2(new_n755), .A3(new_n670), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n755), .B1(new_n738), .B2(new_n670), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n659), .A2(new_n750), .A3(new_n583), .A4(new_n493), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  INV_X1    g576(.A(new_n641), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n740), .A2(new_n582), .A3(new_n572), .A4(new_n622), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(KEYINPUT108), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n650), .B(new_n765), .C1(KEYINPUT108), .C2(new_n764), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n669), .A2(new_n671), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT109), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n767), .B(new_n769), .Z(new_n770));
  OAI211_X1 g584(.A(new_n766), .B(new_n770), .C1(KEYINPUT109), .C2(new_n768), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n743), .A2(new_n745), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n574), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n696), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n767), .A2(new_n311), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n751), .B(new_n775), .C1(new_n758), .C2(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n767), .A2(new_n310), .A3(new_n750), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n773), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n618), .A3(new_n687), .ZN(new_n780));
  INV_X1    g594(.A(new_n574), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n650), .A2(new_n582), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OR3_X1    g597(.A1(new_n783), .A2(new_n389), .A3(new_n595), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n780), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n767), .A2(new_n571), .A3(new_n310), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n775), .B(new_n763), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n786), .B(new_n792), .C1(new_n793), .C2(KEYINPUT51), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n792), .A2(new_n777), .A3(new_n780), .A4(new_n784), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n795), .B(new_n796), .C1(KEYINPUT112), .C2(new_n785), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(G952), .B2(new_n333), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n775), .B2(new_n704), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n595), .A2(new_n389), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n779), .A2(new_n527), .ZN(new_n802));
  OAI221_X1 g616(.A(new_n800), .B1(new_n801), .B2(new_n783), .C1(new_n802), .C2(KEYINPUT48), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(KEYINPUT48), .B2(new_n802), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n794), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n672), .B1(new_n597), .B2(new_n602), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n681), .ZN(new_n807));
  INV_X1    g621(.A(new_n587), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n801), .B1(new_n419), .B2(new_n389), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n579), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n619), .A3(new_n580), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n706), .B1(new_n715), .B2(new_n716), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n750), .A2(new_n420), .A3(new_n389), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n628), .A3(new_n631), .A4(new_n629), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n807), .A2(new_n702), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n725), .A2(new_n727), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n632), .A2(new_n310), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n697), .B2(new_n698), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n615), .A2(new_n610), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n712), .A2(new_n650), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n712), .A2(new_n650), .A3(new_n823), .ZN(new_n826));
  INV_X1    g640(.A(new_n821), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n690), .B2(new_n692), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n828), .A3(KEYINPUT110), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n706), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n634), .B(new_n661), .C1(new_n678), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n832), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n825), .A2(new_n829), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n707), .A2(new_n634), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n840), .A2(new_n834), .A3(new_n836), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n819), .A2(new_n838), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n727), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n719), .B2(new_n724), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n813), .A2(new_n815), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n811), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n845), .A2(new_n702), .A3(new_n847), .A4(new_n807), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n837), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT53), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n843), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n819), .A2(new_n838), .A3(KEYINPUT53), .A4(new_n842), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n839), .B1(new_n848), .B2(new_n849), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(KEYINPUT113), .A2(G953), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n805), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n771), .B1(new_n858), .B2(new_n859), .ZN(G75));
  NOR2_X1   g674(.A1(new_n333), .A2(G952), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n545), .A2(new_n547), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(new_n532), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT55), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NOR4_X1   g679(.A1(new_n848), .A2(new_n849), .A3(new_n839), .A4(new_n841), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n819), .B2(new_n838), .ZN(new_n867));
  OAI21_X1  g681(.A(G902), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n865), .B1(new_n868), .B2(new_n566), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n869), .B2(KEYINPUT114), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n872), .B(new_n865), .C1(new_n868), .C2(new_n566), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n861), .B(new_n870), .C1(new_n874), .C2(new_n864), .ZN(G51));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n305), .B(KEYINPUT57), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n866), .B2(new_n867), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n879), .B2(new_n855), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n664), .B(KEYINPUT115), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n876), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n881), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(KEYINPUT116), .A3(new_n886), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n731), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT117), .B1(new_n868), .B2(new_n731), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n882), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n861), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(G54));
  INV_X1    g706(.A(new_n868), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  INV_X1    g708(.A(new_n382), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n861), .ZN(G60));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n414), .A2(new_n296), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n593), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n879), .B2(new_n855), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n899), .B1(new_n906), .B2(new_n861), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n856), .A2(new_n902), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n593), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n904), .B1(new_n883), .B2(new_n884), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(KEYINPUT119), .A3(new_n891), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n907), .A2(new_n911), .A3(new_n914), .A4(new_n909), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n852), .B2(new_n854), .ZN(new_n921));
  OAI211_X1 g735(.A(KEYINPUT61), .B(new_n891), .C1(new_n921), .C2(new_n524), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n608), .A2(new_n609), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n923), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n891), .B1(new_n921), .B2(new_n524), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n926), .A2(new_n934), .ZN(G66));
  AOI21_X1  g749(.A(new_n333), .B1(new_n575), .B2(G224), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n807), .A2(new_n702), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n812), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n938), .B2(new_n333), .ZN(new_n939));
  INV_X1    g753(.A(G898), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n862), .B1(new_n940), .B2(G953), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  AOI21_X1  g756(.A(new_n753), .B1(new_n758), .B2(new_n760), .ZN(new_n943));
  INV_X1    g757(.A(new_n638), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n527), .A3(new_n751), .A4(new_n809), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n832), .B(KEYINPUT124), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n657), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT62), .B1(new_n657), .B2(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n943), .B(new_n945), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n657), .A2(new_n946), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n657), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n955), .A2(new_n956), .A3(new_n943), .A4(new_n945), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n469), .A2(new_n470), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(new_n375), .Z(new_n959));
  NAND3_X1  g773(.A1(new_n950), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n697), .A2(new_n698), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n527), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n738), .A2(new_n670), .A3(new_n637), .A4(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n845), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n946), .B1(new_n749), .B2(new_n752), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n761), .B(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n959), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n960), .A2(new_n972), .A3(new_n333), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n971), .A2(G900), .A3(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(G900), .ZN(new_n976));
  OAI221_X1 g790(.A(G953), .B1(new_n254), .B2(new_n976), .C1(new_n959), .C2(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n973), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n642), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n843), .A2(new_n474), .A3(new_n850), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n970), .A2(new_n938), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n984), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n891), .B(new_n986), .C1(new_n988), .C2(new_n474), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n950), .A2(new_n957), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n983), .B1(new_n990), .B2(new_n938), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n642), .B2(new_n991), .ZN(G57));
endmodule


