

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U556 ( .A(n747), .B(n706), .ZN(n735) );
  NAND2_X1 U557 ( .A1(n735), .A2(G2072), .ZN(n707) );
  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n706) );
  XNOR2_X1 U559 ( .A(n757), .B(KEYINPUT32), .ZN(n766) );
  INV_X1 U560 ( .A(G2105), .ZN(n533) );
  XNOR2_X1 U561 ( .A(n537), .B(KEYINPUT97), .ZN(G164) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X2 U563 ( .A(KEYINPUT17), .B(n525), .Z(n885) );
  NAND2_X1 U564 ( .A1(G138), .A2(n885), .ZN(n528) );
  NAND2_X1 U565 ( .A1(n533), .A2(G2104), .ZN(n526) );
  XNOR2_X2 U566 ( .A(n526), .B(KEYINPUT65), .ZN(n884) );
  NAND2_X1 U567 ( .A1(G102), .A2(n884), .ZN(n527) );
  NAND2_X1 U568 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n529), .B(KEYINPUT96), .ZN(n532) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U571 ( .A1(G114), .A2(n881), .ZN(n530) );
  XNOR2_X1 U572 ( .A(KEYINPUT95), .B(n530), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n532), .A2(n531), .ZN(n536) );
  NOR2_X1 U574 ( .A1(G2104), .A2(n533), .ZN(n880) );
  NAND2_X1 U575 ( .A1(n880), .A2(G126), .ZN(n534) );
  XNOR2_X1 U576 ( .A(n534), .B(KEYINPUT94), .ZN(n535) );
  NAND2_X1 U577 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U578 ( .A1(G137), .A2(n885), .ZN(n539) );
  NAND2_X1 U579 ( .A1(G113), .A2(n881), .ZN(n538) );
  NAND2_X1 U580 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U581 ( .A(KEYINPUT66), .B(n540), .Z(n542) );
  NAND2_X1 U582 ( .A1(n880), .A2(G125), .ZN(n541) );
  NAND2_X1 U583 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U584 ( .A1(G101), .A2(n884), .ZN(n543) );
  XNOR2_X1 U585 ( .A(KEYINPUT23), .B(n543), .ZN(n544) );
  NOR2_X1 U586 ( .A1(n545), .A2(n544), .ZN(G160) );
  INV_X1 U587 ( .A(G96), .ZN(G221) );
  XOR2_X1 U588 ( .A(G2443), .B(G2446), .Z(n547) );
  XNOR2_X1 U589 ( .A(G2427), .B(G2451), .ZN(n546) );
  XNOR2_X1 U590 ( .A(n547), .B(n546), .ZN(n553) );
  XOR2_X1 U591 ( .A(G2430), .B(G2454), .Z(n549) );
  XNOR2_X1 U592 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U593 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U594 ( .A(G2435), .B(G2438), .Z(n550) );
  XNOR2_X1 U595 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U596 ( .A(n553), .B(n552), .Z(n554) );
  AND2_X1 U597 ( .A1(G14), .A2(n554), .ZN(G401) );
  INV_X1 U598 ( .A(G651), .ZN(n560) );
  NOR2_X1 U599 ( .A1(G543), .A2(n560), .ZN(n555) );
  XOR2_X1 U600 ( .A(KEYINPUT1), .B(n555), .Z(n674) );
  NAND2_X1 U601 ( .A1(n674), .A2(G64), .ZN(n558) );
  XOR2_X1 U602 ( .A(G543), .B(KEYINPUT0), .Z(n660) );
  NOR2_X1 U603 ( .A1(G651), .A2(n660), .ZN(n556) );
  XNOR2_X1 U604 ( .A(KEYINPUT64), .B(n556), .ZN(n675) );
  NAND2_X1 U605 ( .A1(G52), .A2(n675), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n558), .A2(n557), .ZN(n565) );
  NOR2_X1 U607 ( .A1(G651), .A2(G543), .ZN(n671) );
  NAND2_X1 U608 ( .A1(n671), .A2(G90), .ZN(n559) );
  XNOR2_X1 U609 ( .A(n559), .B(KEYINPUT70), .ZN(n562) );
  NOR2_X1 U610 ( .A1(n660), .A2(n560), .ZN(n672) );
  NAND2_X1 U611 ( .A1(G77), .A2(n672), .ZN(n561) );
  NAND2_X1 U612 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U614 ( .A1(n565), .A2(n564), .ZN(G171) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U616 ( .A1(G123), .A2(n880), .ZN(n566) );
  XNOR2_X1 U617 ( .A(n566), .B(KEYINPUT18), .ZN(n573) );
  NAND2_X1 U618 ( .A1(G99), .A2(n884), .ZN(n568) );
  NAND2_X1 U619 ( .A1(G135), .A2(n885), .ZN(n567) );
  NAND2_X1 U620 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U621 ( .A1(G111), .A2(n881), .ZN(n569) );
  XNOR2_X1 U622 ( .A(KEYINPUT81), .B(n569), .ZN(n570) );
  NOR2_X1 U623 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U624 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U625 ( .A(KEYINPUT82), .B(n574), .ZN(n930) );
  XNOR2_X1 U626 ( .A(n930), .B(G2096), .ZN(n575) );
  OR2_X1 U627 ( .A1(G2100), .A2(n575), .ZN(G156) );
  INV_X1 U628 ( .A(G860), .ZN(n641) );
  NAND2_X1 U629 ( .A1(n671), .A2(G81), .ZN(n576) );
  XNOR2_X1 U630 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U631 ( .A1(G68), .A2(n672), .ZN(n577) );
  NAND2_X1 U632 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U633 ( .A(n579), .B(KEYINPUT13), .ZN(n581) );
  NAND2_X1 U634 ( .A1(G43), .A2(n675), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U636 ( .A1(n674), .A2(G56), .ZN(n582) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n582), .Z(n583) );
  NOR2_X1 U638 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U639 ( .A(KEYINPUT74), .B(n585), .Z(n983) );
  OR2_X1 U640 ( .A1(n641), .A2(n983), .ZN(G153) );
  INV_X1 U641 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U642 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U643 ( .A1(G120), .A2(G69), .ZN(n586) );
  NOR2_X1 U644 ( .A1(G237), .A2(n586), .ZN(n587) );
  XNOR2_X1 U645 ( .A(KEYINPUT92), .B(n587), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n588), .A2(G108), .ZN(n895) );
  NAND2_X1 U647 ( .A1(G567), .A2(n895), .ZN(n589) );
  XNOR2_X1 U648 ( .A(n589), .B(KEYINPUT93), .ZN(n596) );
  NAND2_X1 U649 ( .A1(G132), .A2(G82), .ZN(n590) );
  XNOR2_X1 U650 ( .A(n590), .B(KEYINPUT90), .ZN(n591) );
  XNOR2_X1 U651 ( .A(n591), .B(KEYINPUT22), .ZN(n592) );
  NOR2_X1 U652 ( .A1(G218), .A2(n592), .ZN(n593) );
  XNOR2_X1 U653 ( .A(n593), .B(KEYINPUT91), .ZN(n594) );
  OR2_X1 U654 ( .A1(G221), .A2(n594), .ZN(n896) );
  AND2_X1 U655 ( .A1(G2106), .A2(n896), .ZN(n595) );
  NOR2_X1 U656 ( .A1(n596), .A2(n595), .ZN(G319) );
  NAND2_X1 U657 ( .A1(G75), .A2(n672), .ZN(n598) );
  NAND2_X1 U658 ( .A1(G88), .A2(n671), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U660 ( .A(KEYINPUT85), .B(n599), .ZN(n603) );
  NAND2_X1 U661 ( .A1(n675), .A2(G50), .ZN(n601) );
  NAND2_X1 U662 ( .A1(n674), .A2(G62), .ZN(n600) );
  AND2_X1 U663 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n603), .A2(n602), .ZN(G303) );
  NAND2_X1 U665 ( .A1(G78), .A2(n672), .ZN(n605) );
  NAND2_X1 U666 ( .A1(G91), .A2(n671), .ZN(n604) );
  NAND2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U668 ( .A1(G53), .A2(n675), .ZN(n606) );
  XNOR2_X1 U669 ( .A(KEYINPUT71), .B(n606), .ZN(n607) );
  NOR2_X1 U670 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U671 ( .A1(n674), .A2(G65), .ZN(n609) );
  NAND2_X1 U672 ( .A1(n610), .A2(n609), .ZN(G299) );
  NAND2_X1 U673 ( .A1(n672), .A2(G76), .ZN(n611) );
  XNOR2_X1 U674 ( .A(KEYINPUT78), .B(n611), .ZN(n615) );
  XOR2_X1 U675 ( .A(KEYINPUT77), .B(KEYINPUT4), .Z(n613) );
  NAND2_X1 U676 ( .A1(G89), .A2(n671), .ZN(n612) );
  XNOR2_X1 U677 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U678 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U679 ( .A(n616), .B(KEYINPUT5), .ZN(n622) );
  NAND2_X1 U680 ( .A1(G51), .A2(n675), .ZN(n617) );
  XOR2_X1 U681 ( .A(KEYINPUT79), .B(n617), .Z(n619) );
  NAND2_X1 U682 ( .A1(n674), .A2(G63), .ZN(n618) );
  NAND2_X1 U683 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U684 ( .A(KEYINPUT6), .B(n620), .Z(n621) );
  NAND2_X1 U685 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U686 ( .A(n623), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U687 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U688 ( .A1(G7), .A2(G661), .ZN(n624) );
  XNOR2_X1 U689 ( .A(n624), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U690 ( .A(G223), .B(KEYINPUT72), .Z(n842) );
  NAND2_X1 U691 ( .A1(n842), .A2(G567), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n625), .B(KEYINPUT73), .ZN(n626) );
  XNOR2_X1 U693 ( .A(KEYINPUT11), .B(n626), .ZN(G234) );
  INV_X1 U694 ( .A(G171), .ZN(G301) );
  NAND2_X1 U695 ( .A1(G868), .A2(G301), .ZN(n637) );
  NAND2_X1 U696 ( .A1(n672), .A2(G79), .ZN(n628) );
  NAND2_X1 U697 ( .A1(G54), .A2(n675), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT76), .B(n629), .ZN(n634) );
  NAND2_X1 U700 ( .A1(G66), .A2(n674), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G92), .A2(n671), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT75), .B(n632), .Z(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT15), .B(n635), .Z(n988) );
  INV_X1 U706 ( .A(n988), .ZN(n724) );
  INV_X1 U707 ( .A(G868), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n724), .A2(n638), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(G284) );
  NOR2_X1 U710 ( .A1(G286), .A2(n638), .ZN(n640) );
  NOR2_X1 U711 ( .A1(G868), .A2(G299), .ZN(n639) );
  NOR2_X1 U712 ( .A1(n640), .A2(n639), .ZN(G297) );
  NAND2_X1 U713 ( .A1(G559), .A2(n641), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT80), .B(n642), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n643), .A2(n988), .ZN(n644) );
  XNOR2_X1 U716 ( .A(KEYINPUT16), .B(n644), .ZN(G148) );
  NOR2_X1 U717 ( .A1(n983), .A2(G868), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n988), .A2(G868), .ZN(n645) );
  NOR2_X1 U719 ( .A1(G559), .A2(n645), .ZN(n646) );
  NOR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(G282) );
  NAND2_X1 U721 ( .A1(n674), .A2(G67), .ZN(n649) );
  NAND2_X1 U722 ( .A1(G55), .A2(n675), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n654) );
  NAND2_X1 U724 ( .A1(G80), .A2(n672), .ZN(n651) );
  NAND2_X1 U725 ( .A1(G93), .A2(n671), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U727 ( .A(KEYINPUT83), .B(n652), .Z(n653) );
  NOR2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n688) );
  NAND2_X1 U729 ( .A1(n988), .A2(G559), .ZN(n695) );
  XNOR2_X1 U730 ( .A(n983), .B(n695), .ZN(n655) );
  NOR2_X1 U731 ( .A1(G860), .A2(n655), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n688), .B(n656), .ZN(G145) );
  NAND2_X1 U733 ( .A1(G651), .A2(G74), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G49), .A2(n675), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U736 ( .A1(n674), .A2(n659), .ZN(n662) );
  NAND2_X1 U737 ( .A1(n660), .A2(G87), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G288) );
  NAND2_X1 U739 ( .A1(n675), .A2(G48), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n663), .B(KEYINPUT84), .ZN(n670) );
  NAND2_X1 U741 ( .A1(G61), .A2(n674), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G86), .A2(n671), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U744 ( .A1(n672), .A2(G73), .ZN(n666) );
  XOR2_X1 U745 ( .A(KEYINPUT2), .B(n666), .Z(n667) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(G305) );
  NAND2_X1 U748 ( .A1(n671), .A2(G85), .ZN(n682) );
  NAND2_X1 U749 ( .A1(n672), .A2(G72), .ZN(n673) );
  XNOR2_X1 U750 ( .A(KEYINPUT67), .B(n673), .ZN(n680) );
  NAND2_X1 U751 ( .A1(n674), .A2(G60), .ZN(n677) );
  NAND2_X1 U752 ( .A1(G47), .A2(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U754 ( .A(KEYINPUT68), .B(n678), .ZN(n679) );
  NOR2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U756 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U757 ( .A(KEYINPUT69), .B(n683), .Z(G290) );
  NOR2_X1 U758 ( .A1(G868), .A2(n688), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n684), .B(KEYINPUT89), .ZN(n698) );
  XOR2_X1 U760 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n686) );
  XNOR2_X1 U761 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n685) );
  XNOR2_X1 U762 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U763 ( .A(n688), .B(n687), .Z(n689) );
  XNOR2_X1 U764 ( .A(G288), .B(n689), .ZN(n692) );
  XNOR2_X1 U765 ( .A(n983), .B(G299), .ZN(n690) );
  XNOR2_X1 U766 ( .A(n690), .B(G305), .ZN(n691) );
  XNOR2_X1 U767 ( .A(n692), .B(n691), .ZN(n694) );
  XOR2_X1 U768 ( .A(G290), .B(G303), .Z(n693) );
  XNOR2_X1 U769 ( .A(n694), .B(n693), .ZN(n846) );
  XNOR2_X1 U770 ( .A(n846), .B(n695), .ZN(n696) );
  NAND2_X1 U771 ( .A1(G868), .A2(n696), .ZN(n697) );
  NAND2_X1 U772 ( .A1(n698), .A2(n697), .ZN(G295) );
  NAND2_X1 U773 ( .A1(G2078), .A2(G2084), .ZN(n699) );
  XOR2_X1 U774 ( .A(KEYINPUT20), .B(n699), .Z(n700) );
  NAND2_X1 U775 ( .A1(G2090), .A2(n700), .ZN(n701) );
  XNOR2_X1 U776 ( .A(KEYINPUT21), .B(n701), .ZN(n702) );
  NAND2_X1 U777 ( .A1(n702), .A2(G2072), .ZN(G158) );
  INV_X1 U778 ( .A(G319), .ZN(n704) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n703) );
  NOR2_X1 U780 ( .A1(n704), .A2(n703), .ZN(n845) );
  NAND2_X1 U781 ( .A1(n845), .A2(G36), .ZN(G176) );
  NOR2_X1 U782 ( .A1(G164), .A2(G1384), .ZN(n789) );
  NAND2_X1 U783 ( .A1(G160), .A2(G40), .ZN(n790) );
  INV_X1 U784 ( .A(n790), .ZN(n705) );
  NAND2_X2 U785 ( .A1(n789), .A2(n705), .ZN(n747) );
  XOR2_X1 U786 ( .A(n707), .B(KEYINPUT27), .Z(n710) );
  INV_X1 U787 ( .A(n735), .ZN(n708) );
  NAND2_X1 U788 ( .A1(n708), .A2(G1956), .ZN(n709) );
  NAND2_X1 U789 ( .A1(n710), .A2(n709), .ZN(n729) );
  NOR2_X1 U790 ( .A1(G299), .A2(n729), .ZN(n711) );
  XNOR2_X1 U791 ( .A(n711), .B(KEYINPUT107), .ZN(n728) );
  XNOR2_X1 U792 ( .A(G1996), .B(KEYINPUT103), .ZN(n955) );
  NOR2_X1 U793 ( .A1(n747), .A2(n955), .ZN(n712) );
  XNOR2_X1 U794 ( .A(n712), .B(KEYINPUT26), .ZN(n713) );
  NOR2_X1 U795 ( .A1(n983), .A2(n713), .ZN(n715) );
  NAND2_X1 U796 ( .A1(G1341), .A2(n747), .ZN(n714) );
  NAND2_X1 U797 ( .A1(n715), .A2(n714), .ZN(n723) );
  NOR2_X1 U798 ( .A1(n724), .A2(n723), .ZN(n716) );
  XOR2_X1 U799 ( .A(n716), .B(KEYINPUT104), .Z(n722) );
  NAND2_X1 U800 ( .A1(G1348), .A2(n747), .ZN(n717) );
  XOR2_X1 U801 ( .A(KEYINPUT105), .B(n717), .Z(n719) );
  NAND2_X1 U802 ( .A1(G2067), .A2(n735), .ZN(n718) );
  NAND2_X1 U803 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U804 ( .A(KEYINPUT106), .B(n720), .ZN(n721) );
  NAND2_X1 U805 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U806 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U807 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U808 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U809 ( .A1(G299), .A2(n729), .ZN(n730) );
  XNOR2_X1 U810 ( .A(n730), .B(KEYINPUT28), .ZN(n731) );
  NAND2_X1 U811 ( .A1(n732), .A2(n731), .ZN(n734) );
  XOR2_X1 U812 ( .A(KEYINPUT108), .B(KEYINPUT29), .Z(n733) );
  XNOR2_X1 U813 ( .A(n734), .B(n733), .ZN(n739) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NAND2_X1 U815 ( .A1(n735), .A2(n956), .ZN(n737) );
  INV_X1 U816 ( .A(G1961), .ZN(n1019) );
  NAND2_X1 U817 ( .A1(n1019), .A2(n747), .ZN(n736) );
  NAND2_X1 U818 ( .A1(n737), .A2(n736), .ZN(n743) );
  NAND2_X1 U819 ( .A1(n743), .A2(G171), .ZN(n738) );
  NAND2_X1 U820 ( .A1(n739), .A2(n738), .ZN(n760) );
  NAND2_X1 U821 ( .A1(G8), .A2(n747), .ZN(n819) );
  NOR2_X1 U822 ( .A1(G1966), .A2(n819), .ZN(n762) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n747), .ZN(n758) );
  NOR2_X1 U824 ( .A1(n762), .A2(n758), .ZN(n740) );
  NAND2_X1 U825 ( .A1(G8), .A2(n740), .ZN(n741) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n741), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G168), .A2(n742), .ZN(n745) );
  NOR2_X1 U828 ( .A1(G171), .A2(n743), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n746), .Z(n759) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n819), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n750), .A2(G303), .ZN(n752) );
  AND2_X1 U835 ( .A1(n759), .A2(n752), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n760), .A2(n751), .ZN(n755) );
  INV_X1 U837 ( .A(n752), .ZN(n753) );
  OR2_X1 U838 ( .A1(n753), .A2(G286), .ZN(n754) );
  AND2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U840 ( .A1(n756), .A2(G8), .ZN(n757) );
  NAND2_X1 U841 ( .A1(G8), .A2(n758), .ZN(n764) );
  AND2_X1 U842 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U843 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U845 ( .A1(n766), .A2(n765), .ZN(n815) );
  NOR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U847 ( .A1(G1971), .A2(G303), .ZN(n977) );
  XOR2_X1 U848 ( .A(n977), .B(KEYINPUT109), .Z(n767) );
  NOR2_X1 U849 ( .A1(n978), .A2(n767), .ZN(n769) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n768) );
  AND2_X1 U851 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U852 ( .A1(n815), .A2(n770), .ZN(n774) );
  INV_X1 U853 ( .A(n819), .ZN(n771) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n979) );
  AND2_X1 U855 ( .A1(n771), .A2(n979), .ZN(n772) );
  OR2_X1 U856 ( .A1(KEYINPUT33), .A2(n772), .ZN(n773) );
  NAND2_X1 U857 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U858 ( .A(n775), .B(KEYINPUT110), .ZN(n778) );
  NAND2_X1 U859 ( .A1(n978), .A2(KEYINPUT33), .ZN(n776) );
  NOR2_X1 U860 ( .A1(n819), .A2(n776), .ZN(n777) );
  NOR2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n811) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n991) );
  XNOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NAND2_X1 U864 ( .A1(n885), .A2(G140), .ZN(n779) );
  XOR2_X1 U865 ( .A(KEYINPUT99), .B(n779), .Z(n781) );
  NAND2_X1 U866 ( .A1(n884), .A2(G104), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U868 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G128), .A2(n880), .ZN(n784) );
  NAND2_X1 U870 ( .A1(G116), .A2(n881), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U872 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT36), .B(n788), .ZN(n868) );
  NOR2_X1 U875 ( .A1(n826), .A2(n868), .ZN(n932) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U877 ( .A(n791), .B(KEYINPUT98), .ZN(n837) );
  NAND2_X1 U878 ( .A1(n932), .A2(n837), .ZN(n834) );
  NAND2_X1 U879 ( .A1(n884), .A2(G105), .ZN(n793) );
  XNOR2_X1 U880 ( .A(KEYINPUT100), .B(KEYINPUT38), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n793), .B(n792), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G129), .A2(n880), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G117), .A2(n881), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G141), .A2(n885), .ZN(n796) );
  XNOR2_X1 U886 ( .A(KEYINPUT101), .B(n796), .ZN(n797) );
  NOR2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n867) );
  AND2_X1 U889 ( .A1(n867), .A2(G1996), .ZN(n931) );
  NAND2_X1 U890 ( .A1(G95), .A2(n884), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G119), .A2(n880), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G131), .A2(n885), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G107), .A2(n881), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n871) );
  AND2_X1 U897 ( .A1(n871), .A2(G1991), .ZN(n928) );
  OR2_X1 U898 ( .A1(n931), .A2(n928), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n837), .A2(n807), .ZN(n827) );
  NAND2_X1 U900 ( .A1(n834), .A2(n827), .ZN(n809) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n995) );
  AND2_X1 U902 ( .A1(n995), .A2(n837), .ZN(n808) );
  NOR2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n812) );
  AND2_X1 U904 ( .A1(n991), .A2(n812), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n825) );
  INV_X1 U906 ( .A(n812), .ZN(n823) );
  NOR2_X1 U907 ( .A1(G2090), .A2(G303), .ZN(n813) );
  NAND2_X1 U908 ( .A1(G8), .A2(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n819), .ZN(n821) );
  NOR2_X1 U911 ( .A1(G1981), .A2(G305), .ZN(n817) );
  XOR2_X1 U912 ( .A(n817), .B(KEYINPUT24), .Z(n818) );
  OR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  AND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  OR2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n840) );
  NAND2_X1 U917 ( .A1(n826), .A2(n868), .ZN(n943) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n867), .ZN(n925) );
  INV_X1 U919 ( .A(n827), .ZN(n831) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n871), .ZN(n927) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U922 ( .A1(n927), .A2(n828), .ZN(n829) );
  XOR2_X1 U923 ( .A(KEYINPUT111), .B(n829), .Z(n830) );
  NOR2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U925 ( .A1(n925), .A2(n832), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n833), .B(KEYINPUT39), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U928 ( .A1(n943), .A2(n836), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U931 ( .A(KEYINPUT40), .B(n841), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U934 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n845), .A2(n844), .ZN(G188) );
  XOR2_X1 U937 ( .A(G286), .B(n846), .Z(n847) );
  XOR2_X1 U938 ( .A(n988), .B(n847), .Z(n848) );
  XOR2_X1 U939 ( .A(n848), .B(G171), .Z(n849) );
  NOR2_X1 U940 ( .A1(G37), .A2(n849), .ZN(G397) );
  NAND2_X1 U941 ( .A1(n880), .A2(G124), .ZN(n850) );
  XNOR2_X1 U942 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U943 ( .A1(G136), .A2(n885), .ZN(n851) );
  NAND2_X1 U944 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U945 ( .A(n853), .B(KEYINPUT115), .ZN(n855) );
  NAND2_X1 U946 ( .A1(G100), .A2(n884), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U948 ( .A1(n881), .A2(G112), .ZN(n856) );
  XOR2_X1 U949 ( .A(KEYINPUT116), .B(n856), .Z(n857) );
  NOR2_X1 U950 ( .A1(n858), .A2(n857), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G103), .A2(n884), .ZN(n860) );
  NAND2_X1 U952 ( .A1(G139), .A2(n885), .ZN(n859) );
  NAND2_X1 U953 ( .A1(n860), .A2(n859), .ZN(n866) );
  NAND2_X1 U954 ( .A1(G127), .A2(n880), .ZN(n862) );
  NAND2_X1 U955 ( .A1(G115), .A2(n881), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U957 ( .A(KEYINPUT47), .B(n863), .ZN(n864) );
  XNOR2_X1 U958 ( .A(KEYINPUT117), .B(n864), .ZN(n865) );
  NOR2_X1 U959 ( .A1(n866), .A2(n865), .ZN(n939) );
  XNOR2_X1 U960 ( .A(n939), .B(G162), .ZN(n870) );
  XOR2_X1 U961 ( .A(n868), .B(n867), .Z(n869) );
  XNOR2_X1 U962 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U963 ( .A(G164), .B(n871), .Z(n872) );
  XNOR2_X1 U964 ( .A(n872), .B(n930), .ZN(n873) );
  XOR2_X1 U965 ( .A(n874), .B(n873), .Z(n879) );
  XOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT119), .Z(n876) );
  XNOR2_X1 U967 ( .A(KEYINPUT120), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U968 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U969 ( .A(KEYINPUT118), .B(n877), .ZN(n878) );
  XNOR2_X1 U970 ( .A(n879), .B(n878), .ZN(n893) );
  NAND2_X1 U971 ( .A1(G130), .A2(n880), .ZN(n883) );
  NAND2_X1 U972 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U973 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U974 ( .A1(G106), .A2(n884), .ZN(n887) );
  NAND2_X1 U975 ( .A1(G142), .A2(n885), .ZN(n886) );
  NAND2_X1 U976 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  NOR2_X1 U978 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U979 ( .A(G160), .B(n891), .ZN(n892) );
  XNOR2_X1 U980 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U981 ( .A1(G37), .A2(n894), .ZN(G395) );
  INV_X1 U983 ( .A(G132), .ZN(G219) );
  INV_X1 U984 ( .A(G120), .ZN(G236) );
  INV_X1 U985 ( .A(G108), .ZN(G238) );
  INV_X1 U986 ( .A(G82), .ZN(G220) );
  INV_X1 U987 ( .A(G69), .ZN(G235) );
  NOR2_X1 U988 ( .A1(n896), .A2(n895), .ZN(G325) );
  INV_X1 U989 ( .A(G325), .ZN(G261) );
  XOR2_X1 U990 ( .A(KEYINPUT41), .B(G1976), .Z(n898) );
  XOR2_X1 U991 ( .A(n1019), .B(G1956), .Z(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U993 ( .A(n899), .B(KEYINPUT114), .Z(n901) );
  XNOR2_X1 U994 ( .A(G1996), .B(G1991), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U996 ( .A(G1981), .B(G1971), .Z(n903) );
  XNOR2_X1 U997 ( .A(G1986), .B(G1966), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U999 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1000 ( .A(KEYINPUT113), .B(G2474), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(G229) );
  XOR2_X1 U1002 ( .A(G2096), .B(KEYINPUT43), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G2090), .B(G2678), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n910), .B(KEYINPUT112), .Z(n912) );
  XNOR2_X1 U1006 ( .A(G2067), .B(G2072), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1008 ( .A(KEYINPUT42), .B(G2100), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G2078), .B(G2084), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(G227) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G397), .A2(G395), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(KEYINPUT122), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n922), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n923), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n926), .Z(n938) );
  NOR2_X1 U1024 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n936) );
  XNOR2_X1 U1026 ( .A(G160), .B(G2084), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n946) );
  XOR2_X1 U1031 ( .A(G2072), .B(n939), .Z(n941) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n942), .B(KEYINPUT50), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n947), .ZN(n949) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(n950), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1041 ( .A(KEYINPUT124), .B(G34), .Z(n952) );
  XNOR2_X1 U1042 ( .A(G2084), .B(KEYINPUT54), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n952), .B(n951), .ZN(n969) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n967) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1048 ( .A(n955), .B(G32), .Z(n958) );
  XOR2_X1 U1049 ( .A(n956), .B(G27), .Z(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(KEYINPUT123), .B(n961), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n962), .A2(G28), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n965), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1059 ( .A(KEYINPUT55), .B(n970), .Z(n972) );
  INV_X1 U1060 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n973), .ZN(n1028) );
  XNOR2_X1 U1063 ( .A(KEYINPUT56), .B(KEYINPUT125), .ZN(n974) );
  XOR2_X1 U1064 ( .A(G16), .B(n974), .Z(n999) );
  XOR2_X1 U1065 ( .A(G301), .B(G1961), .Z(n976) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n982) );
  NOR2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1070 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1071 ( .A(G299), .B(G1956), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(n983), .B(G1341), .ZN(n984) );
  NOR2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1075 ( .A(G1348), .B(n988), .Z(n989) );
  NOR2_X1 U1076 ( .A1(n990), .A2(n989), .ZN(n997) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n993), .Z(n994) );
  NOR2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1081 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1082 ( .A1(n999), .A2(n998), .ZN(n1026) );
  INV_X1 U1083 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n1002) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(n1004), .B(KEYINPUT58), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1018) );
  XOR2_X1 U1092 ( .A(G1348), .B(KEYINPUT59), .Z(n1007) );
  XNOR2_X1 U1093 ( .A(G4), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G20), .B(G1956), .ZN(n1008) );
  NOR2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G1981), .B(G6), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1014), .B(KEYINPUT60), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(G21), .B(G1966), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(G5), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1108 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1110 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1031), .ZN(G150) );
  INV_X1 U1112 ( .A(G150), .ZN(G311) );
  INV_X1 U1113 ( .A(G303), .ZN(G166) );
endmodule

