//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  XOR2_X1   g000(.A(KEYINPUT24), .B(G110), .Z(new_n187));
  XNOR2_X1  g001(.A(G119), .B(G128), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT73), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(new_n191), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(G146), .B(new_n193), .C1(new_n197), .C2(new_n191), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT23), .B1(new_n203), .B2(G119), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G119), .ZN(new_n205));
  MUX2_X1   g019(.A(KEYINPUT23), .B(new_n204), .S(new_n205), .Z(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G110), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n190), .A2(new_n202), .A3(new_n207), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n206), .A2(G110), .B1(new_n188), .B2(new_n187), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n209), .B(new_n201), .C1(G146), .C2(new_n197), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT22), .B(G137), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n214));
  XOR2_X1   g028(.A(new_n212), .B(new_n214), .Z(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G902), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n208), .A2(new_n210), .A3(new_n215), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT74), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G217), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G234), .B2(new_n218), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT74), .B1(new_n220), .B2(new_n221), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n217), .A2(new_n219), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(G902), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n227), .A2(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT11), .B1(new_n237), .B2(G134), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(G134), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(G137), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n241), .A3(new_n236), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n241), .A3(new_n246), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT66), .A3(G131), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n235), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT65), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n199), .A2(KEYINPUT65), .A3(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT0), .B(G128), .Z(new_n262));
  AND2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n199), .A2(G143), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n259), .A3(G128), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT0), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n255), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n262), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(KEYINPUT69), .C1(new_n266), .C2(new_n265), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n251), .A2(G131), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(new_n248), .A3(new_n247), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT70), .A3(new_n252), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n254), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n264), .A2(new_n259), .A3(G128), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n257), .A2(G146), .ZN(new_n279));
  OAI21_X1  g093(.A(G128), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n261), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n244), .A2(G137), .ZN(new_n283));
  OAI21_X1  g097(.A(G131), .B1(new_n283), .B2(new_n239), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n247), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n275), .A2(KEYINPUT30), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G119), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G119), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT2), .B(G113), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(KEYINPUT0), .A2(new_n276), .B1(new_n261), .B2(new_n262), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n273), .A2(new_n295), .A3(new_n252), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n273), .A2(new_n295), .A3(new_n298), .A4(new_n252), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n247), .A2(new_n284), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT68), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n297), .A2(new_n299), .B1(new_n282), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n286), .B(new_n294), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  INV_X1    g120(.A(G101), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n308), .B(new_n309), .Z(new_n310));
  NAND3_X1  g124(.A1(new_n275), .A2(new_n293), .A3(new_n285), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n313));
  INV_X1    g127(.A(new_n310), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n315));
  NAND2_X1  g129(.A1(new_n297), .A2(new_n299), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n301), .A2(new_n282), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n294), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n319), .B2(new_n311), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n311), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n314), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT31), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n304), .A2(new_n325), .A3(new_n310), .A4(new_n311), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(G472), .A2(G902), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n327), .A2(KEYINPUT32), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT32), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n310), .B1(new_n320), .B2(new_n323), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n304), .A2(new_n314), .A3(new_n311), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n311), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n293), .B1(new_n275), .B2(new_n285), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT28), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n322), .A2(KEYINPUT72), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n311), .A2(new_n339), .A3(new_n321), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n337), .A2(new_n338), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n218), .ZN(new_n343));
  OAI21_X1  g157(.A(G472), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n234), .B1(new_n331), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n327), .A2(new_n328), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT32), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n327), .A2(KEYINPUT32), .A3(new_n328), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n344), .ZN(new_n352));
  INV_X1    g166(.A(new_n234), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT75), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n347), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G221), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT9), .B(G234), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n359), .B2(new_n218), .ZN(new_n360));
  INV_X1    g174(.A(G237), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n213), .A3(G214), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n257), .ZN(new_n363));
  AOI21_X1  g177(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n364));
  OAI211_X1 g178(.A(KEYINPUT17), .B(G131), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n200), .A2(new_n365), .A3(new_n201), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT89), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n363), .A2(new_n364), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n236), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  OAI21_X1  g184(.A(G131), .B1(new_n363), .B2(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT89), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n200), .A2(new_n365), .A3(new_n373), .A4(new_n201), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT18), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n368), .B1(new_n379), .B2(new_n236), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n197), .B(G146), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n380), .B(new_n381), .C1(new_n371), .C2(new_n379), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n369), .A2(new_n371), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n194), .A2(new_n196), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n386));
  AND2_X1   g200(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n199), .C1(new_n385), .C2(new_n386), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n384), .A2(new_n201), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n382), .ZN(new_n391));
  INV_X1    g205(.A(new_n378), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT90), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(G475), .B1(new_n383), .B2(new_n393), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT20), .A3(new_n218), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT20), .B1(new_n398), .B2(new_n218), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G475), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n394), .A2(new_n403), .A3(new_n218), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n397), .ZN(new_n406));
  INV_X1    g220(.A(new_n383), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n378), .B1(new_n375), .B2(new_n382), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n218), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n405), .A2(new_n406), .B1(new_n409), .B2(G475), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  AOI211_X1 g225(.A(G953), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n218), .B(new_n213), .C1(G234), .C2(G237), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT21), .B(G898), .Z(new_n416));
  OAI21_X1  g230(.A(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G116), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n289), .A2(KEYINPUT14), .A3(G122), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G107), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT91), .ZN(new_n423));
  XOR2_X1   g237(.A(G128), .B(G143), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G134), .ZN(new_n425));
  XNOR2_X1  g239(.A(G128), .B(G143), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n244), .ZN(new_n427));
  INV_X1    g241(.A(G107), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n425), .A2(new_n427), .B1(new_n428), .B2(new_n418), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT91), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n420), .A2(new_n430), .A3(G107), .A4(new_n421), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n423), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n418), .B(new_n428), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n257), .A3(G128), .ZN(new_n435));
  OAI211_X1 g249(.A(G134), .B(new_n435), .C1(new_n424), .C2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n436), .A3(new_n427), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n358), .A2(new_n225), .A3(G953), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n432), .A2(new_n437), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n218), .ZN(new_n444));
  INV_X1    g258(.A(G478), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n445), .A2(KEYINPUT15), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n444), .B(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n402), .A2(new_n410), .A3(new_n417), .A4(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n213), .A2(G227), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n449), .B(new_n450), .Z(new_n451));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n278), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n276), .A2(KEYINPUT78), .A3(new_n277), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n264), .A2(new_n259), .ZN(new_n455));
  INV_X1    g269(.A(new_n280), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT3), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n428), .A3(G104), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n377), .A2(G107), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n458), .A2(new_n460), .A3(new_n307), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n377), .A2(G107), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n428), .A2(G104), .ZN(new_n464));
  OAI21_X1  g278(.A(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT79), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n462), .B2(new_n465), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n282), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n457), .A2(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n252), .A3(new_n273), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n254), .A2(new_n274), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT76), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n462), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(new_n482), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n481), .A2(new_n485), .A3(G101), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n482), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT77), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n271), .B(new_n484), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n282), .B(KEYINPUT10), .C1(new_n470), .C2(new_n471), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n466), .A2(KEYINPUT79), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n469), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT10), .A4(new_n282), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n457), .A2(new_n467), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT10), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n495), .A2(new_n502), .A3(new_n478), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n451), .B1(new_n480), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(KEYINPUT81), .A3(new_n451), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT81), .B1(new_n506), .B2(new_n451), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n495), .A2(new_n505), .A3(new_n502), .ZN(new_n511));
  INV_X1    g325(.A(new_n478), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n512), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n507), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G469), .B1(new_n518), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(G469), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n451), .B1(new_n517), .B2(new_n506), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n506), .A2(new_n451), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n479), .B2(new_n477), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n520), .B(new_n218), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  AOI211_X1 g338(.A(new_n360), .B(new_n448), .C1(new_n519), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n291), .A2(new_n292), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n529), .A2(new_n288), .A3(new_n290), .ZN(new_n530));
  OAI21_X1  g344(.A(G113), .B1(new_n529), .B2(new_n288), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n472), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n492), .A2(KEYINPUT77), .A3(new_n493), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n483), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n533), .B1(new_n536), .B2(new_n294), .ZN(new_n537));
  XOR2_X1   g351(.A(G110), .B(G122), .Z(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n527), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n294), .B(new_n484), .C1(new_n491), .C2(new_n494), .ZN(new_n541));
  INV_X1    g355(.A(new_n533), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n473), .A2(new_n195), .ZN(new_n546));
  OAI21_X1  g360(.A(G125), .B1(new_n263), .B2(new_n267), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT85), .B(G224), .Z(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n213), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n548), .B(new_n550), .Z(new_n551));
  AOI211_X1 g365(.A(new_n293), .B(new_n483), .C1(new_n534), .C2(new_n535), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n527), .B(new_n538), .C1(new_n552), .C2(new_n533), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT84), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT84), .B1(new_n543), .B2(new_n527), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n545), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n548), .A2(KEYINPUT86), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n538), .B(KEYINPUT8), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT5), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n499), .B(new_n528), .C1(new_n531), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n532), .A2(new_n466), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT86), .B1(new_n548), .B2(new_n558), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n537), .A2(new_n539), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT7), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n557), .A2(new_n218), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G210), .B1(G237), .B2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n557), .A2(new_n218), .A3(new_n572), .A4(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G214), .B1(G237), .B2(G902), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n526), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  AOI211_X1 g393(.A(KEYINPUT87), .B(new_n579), .C1(new_n574), .C2(new_n575), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n525), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n356), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n307), .ZN(G3));
  AOI21_X1  g397(.A(new_n360), .B1(new_n519), .B2(new_n524), .ZN(new_n584));
  INV_X1    g398(.A(G472), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n327), .B2(new_n218), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n327), .B2(new_n328), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n587), .A3(new_n353), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n579), .B1(new_n574), .B2(new_n575), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n402), .A2(new_n410), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT33), .B1(new_n439), .B2(KEYINPUT92), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n443), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n441), .B2(new_n442), .ZN(new_n596));
  OAI21_X1  g410(.A(G478), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n443), .A2(new_n445), .A3(new_n218), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n445), .A2(new_n218), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n590), .A2(new_n417), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n589), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT93), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT34), .B(G104), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  NAND2_X1  g421(.A1(new_n404), .A2(new_n396), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n409), .A2(G475), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n399), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n610), .A2(new_n447), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n417), .B(KEYINPUT94), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n590), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  OAI211_X1 g431(.A(new_n525), .B(new_n587), .C1(new_n578), .C2(new_n580), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n216), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n211), .B(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n227), .A2(new_n229), .B1(new_n233), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT37), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  NAND2_X1  g440(.A1(new_n519), .A2(new_n524), .ZN(new_n627));
  INV_X1    g441(.A(new_n360), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n352), .A2(new_n627), .A3(new_n628), .A4(new_n622), .ZN(new_n629));
  INV_X1    g443(.A(G900), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n412), .B1(new_n414), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n590), .A2(new_n611), .A3(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n203), .ZN(G30));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n576), .B(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n592), .A2(new_n447), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n637), .A2(new_n579), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n631), .B(KEYINPUT39), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n584), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n643), .A2(KEYINPUT40), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n304), .A2(new_n311), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n310), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n335), .A2(new_n336), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n647), .B2(new_n314), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n585), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n329), .A2(new_n330), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n622), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n643), .A2(KEYINPUT40), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n640), .A2(new_n644), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G143), .ZN(G45));
  NAND2_X1  g468(.A1(new_n553), .A2(new_n554), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n543), .A2(KEYINPUT84), .A3(new_n527), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n655), .A2(new_n656), .B1(new_n544), .B2(new_n540), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n551), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n572), .B1(new_n658), .B2(new_n570), .ZN(new_n659));
  INV_X1    g473(.A(new_n575), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n577), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n601), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n406), .B1(new_n608), .B2(new_n399), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n609), .B1(new_n404), .B2(new_n397), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n662), .B(new_n632), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT95), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n591), .A2(new_n667), .A3(new_n662), .A4(new_n632), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n623), .B1(new_n331), .B2(new_n344), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n670), .A2(KEYINPUT96), .A3(new_n584), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT96), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n576), .A2(new_n577), .A3(new_n666), .A4(new_n668), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n629), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AND3_X1   g491(.A1(new_n511), .A2(KEYINPUT82), .A3(new_n512), .ZN(new_n678));
  AOI21_X1  g492(.A(KEYINPUT82), .B1(new_n511), .B2(new_n512), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n506), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n451), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n523), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(G469), .B1(new_n682), .B2(G902), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT97), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n524), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g499(.A(KEYINPUT97), .B(G469), .C1(new_n682), .C2(G902), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT98), .B1(new_n687), .B2(new_n628), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT98), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n689), .B(new_n360), .C1(new_n685), .C2(new_n686), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n603), .B(new_n345), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  OAI211_X1 g507(.A(new_n345), .B(new_n614), .C1(new_n688), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT99), .B(G116), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G18));
  AOI21_X1  g510(.A(new_n360), .B1(new_n685), .B2(new_n686), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n590), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n352), .A2(new_n622), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n448), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  AND2_X1   g516(.A1(new_n338), .A2(new_n340), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n310), .B1(new_n703), .B2(new_n337), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n313), .A2(new_n326), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n328), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n707), .A2(new_n234), .A3(new_n586), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n661), .A2(new_n639), .A3(new_n612), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n708), .B(new_n709), .C1(new_n688), .C2(new_n690), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT100), .B(G122), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  INV_X1    g526(.A(new_n586), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n622), .A3(new_n706), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n669), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n666), .A2(new_n668), .A3(KEYINPUT101), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n590), .A3(new_n697), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  NAND3_X1  g534(.A1(new_n574), .A2(new_n577), .A3(new_n575), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n584), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n354), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n716), .A2(new_n717), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n724), .A2(KEYINPUT42), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  NAND3_X1  g545(.A1(new_n724), .A2(new_n611), .A3(new_n632), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  INV_X1    g547(.A(KEYINPUT102), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n601), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n597), .A2(KEYINPUT102), .A3(new_n598), .A4(new_n600), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n402), .A3(new_n410), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n592), .A2(KEYINPUT43), .A3(new_n662), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n587), .A2(new_n623), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(KEYINPUT44), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT104), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT44), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n510), .A2(new_n517), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n507), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n518), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(G469), .A2(G902), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n524), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT46), .B1(new_n755), .B2(new_n756), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n628), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n641), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n748), .A2(new_n722), .A3(new_n750), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n760), .B(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n669), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n766), .A3(new_n722), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n331), .A2(new_n344), .A3(new_n234), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n192), .ZN(G42));
  XOR2_X1   g584(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n591), .A2(new_n447), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n613), .B(new_n773), .C1(new_n578), .C2(new_n580), .ZN(new_n774));
  OAI22_X1  g588(.A1(new_n623), .A2(new_n618), .B1(new_n774), .B2(new_n588), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n582), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI221_X1 g591(.A(KEYINPUT108), .B1(new_n618), .B2(new_n623), .C1(new_n588), .C2(new_n774), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n602), .B(new_n613), .C1(new_n578), .C2(new_n580), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n589), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n777), .A2(new_n778), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n691), .A2(new_n694), .A3(new_n710), .A4(new_n701), .ZN(new_n785));
  INV_X1    g599(.A(new_n634), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n661), .A2(new_n639), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n651), .A3(new_n584), .A4(new_n632), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n676), .A2(new_n786), .A3(new_n719), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(KEYINPUT52), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n447), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n610), .A2(new_n791), .A3(new_n631), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n699), .B1(KEYINPUT109), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n723), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT110), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n718), .A2(new_n794), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n795), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n732), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n634), .B1(new_n698), .B2(new_n718), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n676), .A4(new_n788), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n730), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n784), .A2(new_n790), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n790), .A2(new_n808), .A3(new_n806), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n807), .B1(KEYINPUT53), .B2(new_n809), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n691), .A2(new_n694), .A3(new_n710), .A4(new_n701), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n730), .A4(new_n805), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n777), .A2(new_n778), .A3(new_n783), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n801), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT53), .B1(new_n813), .B2(KEYINPUT111), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n772), .B1(new_n810), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n353), .A2(new_n713), .A3(new_n412), .A4(new_n706), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n743), .B2(new_n744), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n722), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n687), .B(KEYINPUT106), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n628), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n826), .A2(new_n827), .B1(KEYINPUT113), .B2(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n824), .A2(new_n579), .A3(new_n637), .A4(new_n697), .ZN(new_n833));
  XOR2_X1   g647(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT115), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT50), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n839), .A3(new_n834), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n697), .A2(new_n412), .A3(new_n722), .ZN(new_n842));
  INV_X1    g656(.A(new_n714), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n745), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n234), .A2(new_n591), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n842), .A2(new_n601), .A3(new_n650), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n841), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n822), .B1(new_n832), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n841), .A2(new_n844), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n722), .B(new_n824), .C1(new_n765), .C2(new_n829), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n842), .A2(new_n345), .A3(new_n745), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT48), .Z(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n411), .A3(G953), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n842), .A2(new_n353), .A3(new_n602), .A4(new_n650), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n848), .A2(new_n851), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n698), .A2(new_n824), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n818), .A2(new_n821), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(G952), .A2(G953), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT116), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n828), .B(KEYINPUT49), .Z(new_n862));
  NAND4_X1  g676(.A1(new_n845), .A2(new_n577), .A3(new_n628), .A4(new_n662), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT105), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n637), .A3(new_n650), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(G75));
  NOR2_X1   g684(.A1(new_n213), .A2(G952), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n810), .A2(new_n817), .A3(new_n218), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(G210), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n873), .B(new_n874), .C1(KEYINPUT118), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n657), .B(new_n551), .Z(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(KEYINPUT119), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n873), .B(new_n875), .C1(KEYINPUT118), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n871), .B1(new_n879), .B2(new_n881), .ZN(G51));
  XOR2_X1   g696(.A(new_n756), .B(KEYINPUT57), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n815), .A2(new_n816), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n807), .A2(KEYINPUT53), .A3(new_n809), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n771), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n771), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT120), .ZN(new_n889));
  INV_X1    g703(.A(new_n682), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n755), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n872), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n871), .B1(new_n893), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n872), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n394), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n871), .ZN(G60));
  AND2_X1   g715(.A1(new_n819), .A2(new_n820), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n887), .B1(new_n902), .B2(KEYINPUT54), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n599), .B(KEYINPUT59), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n903), .A2(new_n904), .B1(new_n596), .B2(new_n594), .ZN(new_n905));
  INV_X1    g719(.A(new_n871), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n594), .A2(new_n596), .ZN(new_n907));
  INV_X1    g721(.A(new_n904), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n907), .B(new_n908), .C1(new_n886), .C2(new_n887), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT60), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n884), .A2(new_n885), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n871), .B1(new_n913), .B2(new_n231), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n621), .B2(new_n913), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT61), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(G66));
  AOI21_X1  g733(.A(new_n213), .B1(new_n549), .B2(new_n416), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n814), .A2(new_n785), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(new_n213), .ZN(new_n923));
  INV_X1    g737(.A(G898), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n657), .B1(new_n924), .B2(G953), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n923), .B(new_n925), .ZN(G69));
  OAI21_X1  g740(.A(new_n286), .B1(new_n302), .B2(new_n303), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n773), .A2(new_n602), .A3(KEYINPUT122), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n356), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n602), .A2(new_n773), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n643), .B1(KEYINPUT122), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n722), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n762), .B(new_n936), .C1(new_n767), .C2(new_n768), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n653), .A2(new_n676), .A3(new_n803), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT62), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n930), .B1(new_n940), .B2(G953), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT123), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n762), .B(new_n732), .C1(new_n767), .C2(new_n768), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n730), .A2(new_n676), .A3(new_n803), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n761), .A2(new_n345), .A3(new_n787), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n213), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(G900), .A2(G953), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n929), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT123), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n930), .C1(new_n940), .C2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n942), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n942), .A2(new_n949), .A3(new_n954), .A4(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n213), .B1(G227), .B2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n953), .A2(new_n957), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  XOR2_X1   g775(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n585), .A2(new_n218), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n922), .ZN(new_n966));
  INV_X1    g780(.A(new_n333), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n871), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n940), .A2(new_n921), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n964), .ZN(new_n971));
  INV_X1    g785(.A(new_n646), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI211_X1 g787(.A(KEYINPUT126), .B(new_n646), .C1(new_n970), .C2(new_n964), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n902), .A2(new_n333), .A3(new_n646), .A4(new_n964), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT127), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n646), .B1(new_n970), .B2(new_n964), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n969), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n968), .A4(new_n976), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n978), .A2(new_n982), .ZN(G57));
endmodule


