

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n714), .A2(n971), .ZN(n719) );
  NOR2_X1 U551 ( .A1(G164), .A2(G1384), .ZN(n706) );
  AND2_X1 U552 ( .A1(n768), .A2(n767), .ZN(n770) );
  AND2_X1 U553 ( .A1(n752), .A2(n751), .ZN(n757) );
  NAND2_X1 U554 ( .A1(n706), .A2(n705), .ZN(n738) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n525) );
  NOR2_X1 U557 ( .A1(n792), .A2(n777), .ZN(n514) );
  AND2_X1 U558 ( .A1(n722), .A2(G1996), .ZN(n711) );
  BUF_X1 U559 ( .A(n738), .Z(n761) );
  NAND2_X1 U560 ( .A1(n749), .A2(n748), .ZN(n759) );
  XNOR2_X1 U561 ( .A(KEYINPUT100), .B(KEYINPUT32), .ZN(n769) );
  XNOR2_X1 U562 ( .A(n770), .B(n769), .ZN(n771) );
  INV_X1 U563 ( .A(G2105), .ZN(n519) );
  AND2_X2 U564 ( .A1(n519), .A2(G2104), .ZN(n856) );
  NOR2_X2 U565 ( .A1(G2104), .A2(n519), .ZN(n851) );
  NOR2_X1 U566 ( .A1(G651), .A2(n621), .ZN(n639) );
  XNOR2_X1 U567 ( .A(n526), .B(n525), .ZN(n527) );
  OR2_X1 U568 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U569 ( .A(n524), .B(KEYINPUT81), .ZN(G164) );
  NAND2_X1 U570 ( .A1(G126), .A2(n851), .ZN(n516) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n852) );
  NAND2_X1 U572 ( .A1(G114), .A2(n852), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U574 ( .A(KEYINPUT80), .B(n517), .ZN(n523) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n518), .Z(n855) );
  NAND2_X1 U576 ( .A1(G138), .A2(n855), .ZN(n521) );
  NAND2_X1 U577 ( .A1(G102), .A2(n856), .ZN(n520) );
  NAND2_X1 U578 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n855), .A2(G137), .ZN(n528) );
  NAND2_X1 U580 ( .A1(G101), .A2(n856), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G125), .A2(n851), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G113), .A2(n852), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(G160) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U587 ( .A(G57), .ZN(G237) );
  INV_X1 U588 ( .A(G651), .ZN(n537) );
  NOR2_X1 U589 ( .A1(G543), .A2(n537), .ZN(n534) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n534), .B(n533), .ZN(n632) );
  NAND2_X1 U592 ( .A1(G64), .A2(n632), .ZN(n536) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  NAND2_X1 U594 ( .A1(G52), .A2(n639), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U596 ( .A1(n621), .A2(n537), .ZN(n635) );
  NAND2_X1 U597 ( .A1(G77), .A2(n635), .ZN(n539) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U599 ( .A1(G90), .A2(n631), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U602 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U603 ( .A1(G75), .A2(n635), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G88), .A2(n631), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G62), .A2(n632), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G50), .A2(n639), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n548), .A2(n547), .ZN(G166) );
  NAND2_X1 U610 ( .A1(n635), .A2(G76), .ZN(n549) );
  XNOR2_X1 U611 ( .A(KEYINPUT70), .B(n549), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(KEYINPUT4), .Z(n551) );
  NAND2_X1 U613 ( .A1(G89), .A2(n631), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G63), .A2(n632), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G51), .A2(n639), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U622 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U626 ( .A(G223), .ZN(n826) );
  NAND2_X1 U627 ( .A1(n826), .A2(G567), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT11), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT67), .B(n563), .ZN(G234) );
  NAND2_X1 U630 ( .A1(G56), .A2(n632), .ZN(n564) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n564), .Z(n571) );
  NAND2_X1 U632 ( .A1(n631), .A2(G81), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT12), .B(n565), .Z(n568) );
  NAND2_X1 U634 ( .A1(n635), .A2(G68), .ZN(n566) );
  XOR2_X1 U635 ( .A(KEYINPUT68), .B(n566), .Z(n567) );
  NOR2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(KEYINPUT13), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n639), .A2(G43), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n971) );
  INV_X1 U641 ( .A(G860), .ZN(n592) );
  OR2_X1 U642 ( .A1(n971), .A2(n592), .ZN(G153) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G79), .A2(n635), .ZN(n575) );
  NAND2_X1 U646 ( .A1(G66), .A2(n632), .ZN(n574) );
  NAND2_X1 U647 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G92), .A2(n631), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G54), .A2(n639), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n580), .Z(n968) );
  OR2_X1 U653 ( .A1(n968), .A2(G868), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G78), .A2(n635), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G65), .A2(n632), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n631), .A2(G91), .ZN(n585) );
  XOR2_X1 U659 ( .A(KEYINPUT66), .B(n585), .Z(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n639), .A2(G53), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G299) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n591) );
  INV_X1 U664 ( .A(G868), .ZN(n653) );
  NOR2_X1 U665 ( .A1(G286), .A2(n653), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n592), .A2(G559), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n593), .A2(n968), .ZN(n594) );
  XNOR2_X1 U669 ( .A(n594), .B(KEYINPUT71), .ZN(n595) );
  XOR2_X1 U670 ( .A(KEYINPUT16), .B(n595), .Z(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n971), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G868), .A2(n968), .ZN(n596) );
  NOR2_X1 U673 ( .A1(G559), .A2(n596), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(G282) );
  NAND2_X1 U675 ( .A1(n851), .A2(G123), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT18), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G111), .A2(n852), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G135), .A2(n855), .ZN(n603) );
  NAND2_X1 U680 ( .A1(G99), .A2(n856), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n918) );
  XNOR2_X1 U683 ( .A(n918), .B(G2096), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT72), .ZN(n608) );
  INV_X1 U685 ( .A(G2100), .ZN(n607) );
  NAND2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n968), .A2(G559), .ZN(n650) );
  XNOR2_X1 U688 ( .A(n971), .B(n650), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n609), .A2(G860), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G80), .A2(n635), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G67), .A2(n632), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G93), .A2(n631), .ZN(n613) );
  NAND2_X1 U694 ( .A1(G55), .A2(n639), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n652) );
  XNOR2_X1 U697 ( .A(n616), .B(n652), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G49), .A2(n639), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U701 ( .A1(n632), .A2(n619), .ZN(n620) );
  XOR2_X1 U702 ( .A(KEYINPUT73), .B(n620), .Z(n623) );
  NAND2_X1 U703 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U705 ( .A1(G72), .A2(n635), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G85), .A2(n631), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT64), .B(n626), .Z(n630) );
  NAND2_X1 U709 ( .A1(G60), .A2(n632), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G47), .A2(n639), .ZN(n627) );
  AND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(G290) );
  NAND2_X1 U713 ( .A1(G86), .A2(n631), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G61), .A2(n632), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n639), .A2(G48), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(G305) );
  XOR2_X1 U721 ( .A(G290), .B(G305), .Z(n642) );
  XNOR2_X1 U722 ( .A(G288), .B(n642), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n644) );
  INV_X1 U724 ( .A(G299), .ZN(n961) );
  XNOR2_X1 U725 ( .A(n961), .B(KEYINPUT19), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U727 ( .A(n646), .B(n645), .Z(n648) );
  XNOR2_X1 U728 ( .A(G166), .B(n652), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(n971), .ZN(n876) );
  XNOR2_X1 U731 ( .A(n876), .B(n650), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n653), .A2(n651), .ZN(n655) );
  AND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U734 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n657) );
  XOR2_X1 U736 ( .A(KEYINPUT76), .B(KEYINPUT20), .Z(n656) );
  XNOR2_X1 U737 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(G2090), .ZN(n659) );
  XOR2_X1 U739 ( .A(KEYINPUT77), .B(n659), .Z(n660) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G132), .A2(G82), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n662), .B(KEYINPUT78), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n663), .B(KEYINPUT22), .ZN(n664) );
  NOR2_X1 U746 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U747 ( .A1(G96), .A2(n665), .ZN(n831) );
  NAND2_X1 U748 ( .A1(G2106), .A2(n831), .ZN(n666) );
  XOR2_X1 U749 ( .A(KEYINPUT79), .B(n666), .Z(n670) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U751 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G108), .A2(n668), .ZN(n832) );
  NAND2_X1 U753 ( .A1(G567), .A2(n832), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n902) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n902), .A2(n671), .ZN(n830) );
  NAND2_X1 U757 ( .A1(n830), .A2(G36), .ZN(G176) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  NAND2_X1 U759 ( .A1(G140), .A2(n855), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G104), .A2(n856), .ZN(n672) );
  NAND2_X1 U761 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U762 ( .A(KEYINPUT34), .B(n674), .ZN(n679) );
  NAND2_X1 U763 ( .A1(G128), .A2(n851), .ZN(n676) );
  NAND2_X1 U764 ( .A1(G116), .A2(n852), .ZN(n675) );
  NAND2_X1 U765 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U766 ( .A(n677), .B(KEYINPUT35), .Z(n678) );
  NOR2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U768 ( .A(KEYINPUT36), .B(n680), .Z(n681) );
  XNOR2_X1 U769 ( .A(KEYINPUT85), .B(n681), .ZN(n869) );
  XNOR2_X1 U770 ( .A(KEYINPUT37), .B(G2067), .ZN(n801) );
  NOR2_X1 U771 ( .A1(n869), .A2(n801), .ZN(n916) );
  NAND2_X1 U772 ( .A1(G40), .A2(G160), .ZN(n704) );
  XOR2_X1 U773 ( .A(KEYINPUT83), .B(n704), .Z(n682) );
  NOR2_X1 U774 ( .A1(n706), .A2(n682), .ZN(n811) );
  NAND2_X1 U775 ( .A1(n916), .A2(n811), .ZN(n683) );
  XNOR2_X1 U776 ( .A(n683), .B(KEYINPUT86), .ZN(n807) );
  NAND2_X1 U777 ( .A1(G129), .A2(n851), .ZN(n685) );
  NAND2_X1 U778 ( .A1(G141), .A2(n855), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n856), .A2(G105), .ZN(n686) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n686), .Z(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n852), .A2(G117), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n842) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n842), .ZN(n700) );
  NAND2_X1 U786 ( .A1(G131), .A2(n855), .ZN(n692) );
  NAND2_X1 U787 ( .A1(G95), .A2(n856), .ZN(n691) );
  NAND2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U789 ( .A(KEYINPUT88), .B(n693), .ZN(n696) );
  NAND2_X1 U790 ( .A1(G107), .A2(n852), .ZN(n694) );
  XNOR2_X1 U791 ( .A(KEYINPUT87), .B(n694), .ZN(n695) );
  NOR2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U793 ( .A1(n851), .A2(G119), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n872) );
  NAND2_X1 U795 ( .A1(G1991), .A2(n872), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U797 ( .A(KEYINPUT89), .B(n701), .ZN(n921) );
  INV_X1 U798 ( .A(n811), .ZN(n702) );
  NOR2_X1 U799 ( .A1(n921), .A2(n702), .ZN(n804) );
  INV_X1 U800 ( .A(n804), .ZN(n703) );
  NAND2_X1 U801 ( .A1(n807), .A2(n703), .ZN(n796) );
  XNOR2_X1 U802 ( .A(n704), .B(KEYINPUT83), .ZN(n705) );
  NAND2_X1 U803 ( .A1(G8), .A2(n738), .ZN(n792) );
  NOR2_X1 U804 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NAND2_X1 U805 ( .A1(n774), .A2(KEYINPUT33), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n792), .A2(n707), .ZN(n781) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n944) );
  NOR2_X1 U808 ( .A1(n944), .A2(n761), .ZN(n708) );
  XOR2_X1 U809 ( .A(KEYINPUT93), .B(n708), .Z(n710) );
  NOR2_X1 U810 ( .A1(n722), .A2(G1961), .ZN(n709) );
  NOR2_X1 U811 ( .A1(n710), .A2(n709), .ZN(n744) );
  OR2_X1 U812 ( .A1(n744), .A2(G301), .ZN(n737) );
  INV_X1 U813 ( .A(n738), .ZN(n722) );
  XOR2_X1 U814 ( .A(n711), .B(KEYINPUT26), .Z(n713) );
  NAND2_X1 U815 ( .A1(n761), .A2(G1341), .ZN(n712) );
  NAND2_X1 U816 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U817 ( .A1(n719), .A2(n968), .ZN(n718) );
  NOR2_X1 U818 ( .A1(G2067), .A2(n761), .ZN(n716) );
  NOR2_X1 U819 ( .A1(n722), .A2(G1348), .ZN(n715) );
  NOR2_X1 U820 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U821 ( .A1(n718), .A2(n717), .ZN(n721) );
  OR2_X1 U822 ( .A1(n968), .A2(n719), .ZN(n720) );
  NAND2_X1 U823 ( .A1(n721), .A2(n720), .ZN(n728) );
  NAND2_X1 U824 ( .A1(G2072), .A2(n722), .ZN(n723) );
  XNOR2_X1 U825 ( .A(n723), .B(KEYINPUT27), .ZN(n724) );
  XNOR2_X1 U826 ( .A(n724), .B(KEYINPUT94), .ZN(n726) );
  AND2_X1 U827 ( .A1(G1956), .A2(n761), .ZN(n725) );
  NOR2_X1 U828 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U829 ( .A1(n729), .A2(n961), .ZN(n727) );
  NAND2_X1 U830 ( .A1(n728), .A2(n727), .ZN(n734) );
  NOR2_X1 U831 ( .A1(n729), .A2(n961), .ZN(n732) );
  XNOR2_X1 U832 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n730) );
  XNOR2_X1 U833 ( .A(n730), .B(KEYINPUT28), .ZN(n731) );
  XNOR2_X1 U834 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U836 ( .A(KEYINPUT29), .B(n735), .Z(n736) );
  NAND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n749) );
  NOR2_X1 U838 ( .A1(G1966), .A2(n792), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G2084), .A2(n738), .ZN(n739) );
  XNOR2_X1 U840 ( .A(KEYINPUT91), .B(n739), .ZN(n753) );
  NAND2_X1 U841 ( .A1(G8), .A2(n753), .ZN(n740) );
  NOR2_X1 U842 ( .A1(n750), .A2(n740), .ZN(n741) );
  XOR2_X1 U843 ( .A(KEYINPUT30), .B(n741), .Z(n742) );
  NOR2_X1 U844 ( .A1(G168), .A2(n742), .ZN(n743) );
  XNOR2_X1 U845 ( .A(n743), .B(KEYINPUT97), .ZN(n746) );
  NAND2_X1 U846 ( .A1(n744), .A2(G301), .ZN(n745) );
  NAND2_X1 U847 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U848 ( .A(KEYINPUT31), .B(n747), .ZN(n748) );
  XNOR2_X1 U849 ( .A(n759), .B(KEYINPUT98), .ZN(n752) );
  INV_X1 U850 ( .A(n750), .ZN(n751) );
  INV_X1 U851 ( .A(n753), .ZN(n754) );
  NAND2_X1 U852 ( .A1(n754), .A2(G8), .ZN(n755) );
  XNOR2_X1 U853 ( .A(n755), .B(KEYINPUT92), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n757), .A2(n756), .ZN(n772) );
  AND2_X1 U855 ( .A1(G286), .A2(G8), .ZN(n758) );
  NAND2_X1 U856 ( .A1(n759), .A2(n758), .ZN(n768) );
  INV_X1 U857 ( .A(G8), .ZN(n766) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n792), .ZN(n760) );
  XNOR2_X1 U859 ( .A(KEYINPUT99), .B(n760), .ZN(n764) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U861 ( .A1(G166), .A2(n762), .ZN(n763) );
  NAND2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n765) );
  OR2_X1 U863 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n965) );
  XOR2_X1 U867 ( .A(n965), .B(KEYINPUT101), .Z(n775) );
  NAND2_X1 U868 ( .A1(n785), .A2(n775), .ZN(n776) );
  XNOR2_X1 U869 ( .A(n776), .B(KEYINPUT102), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n964) );
  INV_X1 U871 ( .A(n964), .ZN(n777) );
  AND2_X1 U872 ( .A1(n778), .A2(n514), .ZN(n779) );
  NOR2_X1 U873 ( .A1(n779), .A2(KEYINPUT33), .ZN(n780) );
  NOR2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U875 ( .A(G1981), .B(G305), .Z(n958) );
  NAND2_X1 U876 ( .A1(n782), .A2(n958), .ZN(n788) );
  NOR2_X1 U877 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U878 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n786), .A2(n792), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n794) );
  NOR2_X1 U882 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U883 ( .A(n789), .B(KEYINPUT90), .Z(n790) );
  XNOR2_X1 U884 ( .A(KEYINPUT24), .B(n790), .ZN(n791) );
  NOR2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT82), .B(G1986), .ZN(n797) );
  XNOR2_X1 U889 ( .A(n797), .B(G290), .ZN(n977) );
  NAND2_X1 U890 ( .A1(n977), .A2(n811), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT84), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n814) );
  NAND2_X1 U893 ( .A1(n869), .A2(n801), .ZN(n910) );
  NOR2_X1 U894 ( .A1(G1996), .A2(n842), .ZN(n913) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n872), .ZN(n917) );
  NOR2_X1 U897 ( .A1(n802), .A2(n917), .ZN(n803) );
  NOR2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U899 ( .A1(n913), .A2(n805), .ZN(n806) );
  XNOR2_X1 U900 ( .A(KEYINPUT39), .B(n806), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n910), .A2(n809), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT103), .B(n812), .Z(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U906 ( .A(n815), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U907 ( .A(G2430), .B(G2435), .ZN(n824) );
  XNOR2_X1 U908 ( .A(G2454), .B(KEYINPUT104), .ZN(n822) );
  XOR2_X1 U909 ( .A(G2451), .B(G2427), .Z(n817) );
  XNOR2_X1 U910 ( .A(G2438), .B(G2446), .ZN(n816) );
  XNOR2_X1 U911 ( .A(n817), .B(n816), .ZN(n818) );
  XOR2_X1 U912 ( .A(n818), .B(G2443), .Z(n820) );
  XNOR2_X1 U913 ( .A(G1348), .B(G1341), .ZN(n819) );
  XNOR2_X1 U914 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U916 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U917 ( .A1(n825), .A2(G14), .ZN(n905) );
  XNOR2_X1 U918 ( .A(KEYINPUT105), .B(n905), .ZN(G401) );
  NAND2_X1 U919 ( .A1(n826), .A2(G2106), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U922 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G188) );
  XNOR2_X1 U925 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U927 ( .A(G132), .ZN(G219) );
  INV_X1 U928 ( .A(G120), .ZN(G236) );
  INV_X1 U929 ( .A(G82), .ZN(G220) );
  INV_X1 U930 ( .A(G69), .ZN(G235) );
  NOR2_X1 U931 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  NAND2_X1 U933 ( .A1(G124), .A2(n851), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n833), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U935 ( .A1(G112), .A2(n852), .ZN(n834) );
  XOR2_X1 U936 ( .A(KEYINPUT113), .B(n834), .Z(n835) );
  NAND2_X1 U937 ( .A1(n836), .A2(n835), .ZN(n840) );
  NAND2_X1 U938 ( .A1(G136), .A2(n855), .ZN(n838) );
  NAND2_X1 U939 ( .A1(G100), .A2(n856), .ZN(n837) );
  NAND2_X1 U940 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U941 ( .A1(n840), .A2(n839), .ZN(G162) );
  XOR2_X1 U942 ( .A(G160), .B(G162), .Z(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n865) );
  NAND2_X1 U944 ( .A1(G127), .A2(n851), .ZN(n844) );
  NAND2_X1 U945 ( .A1(G115), .A2(n852), .ZN(n843) );
  NAND2_X1 U946 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n845), .B(KEYINPUT47), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G139), .A2(n855), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n856), .A2(G103), .ZN(n848) );
  XOR2_X1 U951 ( .A(KEYINPUT114), .B(n848), .Z(n849) );
  NOR2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n922) );
  XNOR2_X1 U953 ( .A(n922), .B(n918), .ZN(n863) );
  NAND2_X1 U954 ( .A1(G130), .A2(n851), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G118), .A2(n852), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G142), .A2(n855), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G106), .A2(n856), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(KEYINPUT45), .B(n859), .Z(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n871) );
  XOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n867) );
  XNOR2_X1 U965 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n871), .B(n870), .ZN(n874) );
  XOR2_X1 U969 ( .A(n872), .B(G164), .Z(n873) );
  XNOR2_X1 U970 ( .A(n874), .B(n873), .ZN(n875) );
  NOR2_X1 U971 ( .A1(G37), .A2(n875), .ZN(G395) );
  XOR2_X1 U972 ( .A(KEYINPUT117), .B(n876), .Z(n878) );
  XNOR2_X1 U973 ( .A(G171), .B(n968), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U975 ( .A(G286), .B(n879), .Z(n880) );
  NOR2_X1 U976 ( .A1(G37), .A2(n880), .ZN(G397) );
  XOR2_X1 U977 ( .A(G1976), .B(G1966), .Z(n882) );
  XNOR2_X1 U978 ( .A(G1986), .B(G1971), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U980 ( .A(n883), .B(KEYINPUT41), .Z(n885) );
  XNOR2_X1 U981 ( .A(G1996), .B(G1991), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n889) );
  XOR2_X1 U983 ( .A(G2474), .B(G1981), .Z(n887) );
  XNOR2_X1 U984 ( .A(G1961), .B(G1956), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(G229) );
  XOR2_X1 U987 ( .A(G2096), .B(G2072), .Z(n891) );
  XNOR2_X1 U988 ( .A(G2067), .B(G2090), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n901) );
  XOR2_X1 U990 ( .A(KEYINPUT112), .B(G2678), .Z(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT111), .B(KEYINPUT109), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U993 ( .A(G2100), .B(KEYINPUT43), .Z(n895) );
  XNOR2_X1 U994 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U997 ( .A(G2078), .B(G2084), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(G227) );
  XOR2_X1 U1000 ( .A(KEYINPUT108), .B(n902), .Z(G319) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G397), .A2(n906), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n907), .A2(G319), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G395), .A2(n908), .ZN(G308) );
  INV_X1 U1007 ( .A(G308), .ZN(G225) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1009 ( .A(G160), .B(G2084), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n909), .B(KEYINPUT118), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n931) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n912) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(n914), .B(KEYINPUT51), .ZN(n915) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n929) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT119), .B(n919), .Z(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1022 ( .A(KEYINPUT50), .B(n925), .Z(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1026 ( .A(KEYINPUT52), .B(n932), .Z(n933) );
  NAND2_X1 U1027 ( .A1(G29), .A2(n933), .ZN(n1012) );
  XOR2_X1 U1028 ( .A(G2090), .B(G35), .Z(n950) );
  XNOR2_X1 U1029 ( .A(KEYINPUT53), .B(KEYINPUT122), .ZN(n934) );
  XNOR2_X1 U1030 ( .A(n934), .B(KEYINPUT123), .ZN(n948) );
  XNOR2_X1 U1031 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n943) );
  XOR2_X1 U1034 ( .A(G1991), .B(G25), .Z(n937) );
  NAND2_X1 U1035 ( .A1(n937), .A2(G28), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT120), .ZN(n941) );
  XOR2_X1 U1037 ( .A(G1996), .B(KEYINPUT121), .Z(n939) );
  XNOR2_X1 U1038 ( .A(G32), .B(n939), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G27), .B(n944), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G34), .B(G2084), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(n954), .B(KEYINPUT124), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(G29), .A2(n955), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT55), .B(n956), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n957), .A2(G11), .ZN(n1010) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n981) );
  XNOR2_X1 U1053 ( .A(G168), .B(G1966), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT57), .ZN(n979) );
  XNOR2_X1 U1056 ( .A(G1956), .B(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(G1971), .A2(G303), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n967) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n975) );
  XNOR2_X1 U1061 ( .A(G1348), .B(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(G1341), .B(n971), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n1008) );
  INV_X1 U1070 ( .A(G16), .ZN(n1006) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1074 ( .A(KEYINPUT126), .B(n984), .Z(n986) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(KEYINPUT58), .B(n987), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1961), .B(G5), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G21), .B(G1966), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n1002) );
  XNOR2_X1 U1082 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(n992), .B(G4), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G1348), .B(n993), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G1956), .B(G20), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT61), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT127), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT62), .B(n1013), .Z(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

