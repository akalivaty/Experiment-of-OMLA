

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777;

  XNOR2_X1 U377 ( .A(n540), .B(KEYINPUT40), .ZN(n664) );
  OR2_X1 U378 ( .A1(n698), .A2(n424), .ZN(n422) );
  BUF_X1 U379 ( .A(G128), .Z(n372) );
  XNOR2_X1 U380 ( .A(G143), .B(G128), .ZN(n374) );
  XNOR2_X1 U381 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n431) );
  OR2_X4 U383 ( .A1(n734), .A2(G902), .ZN(n442) );
  NOR2_X1 U384 ( .A1(n524), .A2(n710), .ZN(n528) );
  BUF_X2 U385 ( .A(n634), .Z(n771) );
  NOR2_X1 U386 ( .A1(n544), .A2(n543), .ZN(n407) );
  XNOR2_X2 U387 ( .A(G146), .B(G125), .ZN(n505) );
  XOR2_X1 U388 ( .A(G143), .B(G128), .Z(n358) );
  NOR2_X1 U389 ( .A1(n658), .A2(G902), .ZN(n382) );
  INV_X1 U390 ( .A(G953), .ZN(n403) );
  XNOR2_X1 U391 ( .A(n542), .B(KEYINPUT85), .ZN(n561) );
  NOR2_X2 U392 ( .A1(n725), .A2(n544), .ZN(n537) );
  NAND2_X2 U393 ( .A1(n421), .A2(n420), .ZN(n725) );
  XNOR2_X2 U394 ( .A(KEYINPUT78), .B(KEYINPUT89), .ZN(n504) );
  XNOR2_X2 U395 ( .A(G137), .B(KEYINPUT94), .ZN(n415) );
  XNOR2_X2 U396 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n508) );
  NAND2_X2 U397 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X2 U398 ( .A(n591), .B(n590), .ZN(n696) );
  NOR2_X2 U399 ( .A1(n609), .A2(n383), .ZN(n591) );
  AND2_X1 U400 ( .A1(n399), .A2(n414), .ZN(n413) );
  XNOR2_X1 U401 ( .A(n561), .B(KEYINPUT19), .ZN(n573) );
  INV_X1 U402 ( .A(KEYINPUT102), .ZN(n417) );
  AND2_X1 U403 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U404 ( .A1(n604), .A2(n355), .ZN(n605) );
  XNOR2_X1 U405 ( .A(n587), .B(n586), .ZN(n599) );
  NAND2_X1 U406 ( .A1(n593), .A2(n592), .ZN(n594) );
  AND2_X1 U407 ( .A1(n423), .A2(n422), .ZN(n421) );
  OR2_X1 U408 ( .A1(n573), .A2(n411), .ZN(n410) );
  XNOR2_X1 U409 ( .A(n418), .B(n417), .ZN(n546) );
  BUF_X1 U410 ( .A(n620), .Z(n383) );
  NOR2_X1 U411 ( .A1(n554), .A2(n367), .ZN(n418) );
  XNOR2_X1 U412 ( .A(n498), .B(n368), .ZN(n367) );
  XOR2_X1 U413 ( .A(n665), .B(KEYINPUT59), .Z(n666) );
  XNOR2_X1 U414 ( .A(n401), .B(KEYINPUT75), .ZN(n484) );
  XNOR2_X1 U415 ( .A(n419), .B(n443), .ZN(n766) );
  XNOR2_X1 U416 ( .A(n449), .B(KEYINPUT8), .ZN(n490) );
  AND2_X1 U417 ( .A1(G234), .A2(n506), .ZN(n449) );
  INV_X1 U418 ( .A(G953), .ZN(n506) );
  XNOR2_X1 U419 ( .A(n594), .B(KEYINPUT35), .ZN(n355) );
  XNOR2_X2 U420 ( .A(n648), .B(n647), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n648), .B(n647), .ZN(n744) );
  NAND2_X2 U422 ( .A1(n646), .A2(n645), .ZN(n648) );
  INV_X1 U423 ( .A(G104), .ZN(n435) );
  INV_X1 U424 ( .A(KEYINPUT68), .ZN(n434) );
  XNOR2_X1 U425 ( .A(n761), .B(n471), .ZN(n518) );
  INV_X1 U426 ( .A(n367), .ZN(n553) );
  NAND2_X1 U427 ( .A1(n579), .A2(KEYINPUT0), .ZN(n414) );
  NAND2_X1 U428 ( .A1(n580), .A2(n412), .ZN(n411) );
  INV_X1 U429 ( .A(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U430 ( .A(G110), .B(KEYINPUT24), .ZN(n444) );
  XOR2_X1 U431 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n443) );
  XNOR2_X2 U432 ( .A(G146), .B(G125), .ZN(n380) );
  XNOR2_X1 U433 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U434 ( .A1(n405), .A2(n404), .ZN(n547) );
  INV_X1 U435 ( .A(n544), .ZN(n404) );
  NOR2_X1 U436 ( .A1(n543), .A2(n406), .ZN(n405) );
  XOR2_X1 U437 ( .A(KEYINPUT5), .B(G146), .Z(n472) );
  NAND2_X1 U438 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U439 ( .A(G902), .B(KEYINPUT15), .ZN(n631) );
  NAND2_X1 U440 ( .A1(n358), .A2(n377), .ZN(n379) );
  INV_X1 U441 ( .A(n431), .ZN(n377) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n456) );
  OR2_X1 U443 ( .A1(n622), .A2(n672), .ZN(n623) );
  XNOR2_X1 U444 ( .A(n569), .B(n568), .ZN(n641) );
  NAND2_X1 U445 ( .A1(n424), .A2(n697), .ZN(n426) );
  NAND2_X1 U446 ( .A1(n359), .A2(n531), .ZN(n423) );
  INV_X1 U447 ( .A(n697), .ZN(n427) );
  NAND2_X1 U448 ( .A1(n520), .A2(G214), .ZN(n697) );
  INV_X1 U449 ( .A(G472), .ZN(n381) );
  XOR2_X1 U450 ( .A(G122), .B(G107), .Z(n494) );
  XNOR2_X1 U451 ( .A(G113), .B(G143), .ZN(n479) );
  XNOR2_X1 U452 ( .A(n471), .B(G146), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n594), .B(KEYINPUT35), .ZN(n603) );
  NOR2_X1 U454 ( .A1(n741), .A2(G902), .ZN(n498) );
  XNOR2_X1 U455 ( .A(n487), .B(G475), .ZN(n488) );
  XNOR2_X1 U456 ( .A(n393), .B(n470), .ZN(n761) );
  XNOR2_X1 U457 ( .A(n469), .B(KEYINPUT88), .ZN(n393) );
  XNOR2_X1 U458 ( .A(G116), .B(G113), .ZN(n469) );
  XNOR2_X1 U459 ( .A(n409), .B(n408), .ZN(n745) );
  XNOR2_X1 U460 ( .A(n766), .B(n450), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n357), .B(n448), .ZN(n408) );
  AND2_X1 U462 ( .A1(n653), .A2(G953), .ZN(n748) );
  BUF_X1 U463 ( .A(n599), .Z(n670) );
  XOR2_X1 U464 ( .A(n447), .B(n446), .Z(n357) );
  OR2_X1 U465 ( .A1(n700), .A2(n427), .ZN(n359) );
  XNOR2_X1 U466 ( .A(KEYINPUT81), .B(n695), .ZN(n360) );
  XOR2_X1 U467 ( .A(n483), .B(n482), .Z(n361) );
  OR2_X1 U468 ( .A1(n700), .A2(n709), .ZN(n362) );
  AND2_X1 U469 ( .A1(n520), .A2(G210), .ZN(n363) );
  INV_X1 U470 ( .A(G237), .ZN(n402) );
  INV_X1 U471 ( .A(n531), .ZN(n424) );
  XOR2_X1 U472 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n364) );
  NAND2_X1 U473 ( .A1(n546), .A2(n545), .ZN(n701) );
  NOR2_X1 U474 ( .A1(n365), .A2(n366), .ZN(n672) );
  NAND2_X1 U475 ( .A1(n621), .A2(n383), .ZN(n365) );
  OR2_X1 U476 ( .A1(n706), .A2(n710), .ZN(n366) );
  XNOR2_X1 U477 ( .A(KEYINPUT101), .B(G478), .ZN(n368) );
  BUF_X1 U478 ( .A(n664), .Z(n369) );
  INV_X1 U479 ( .A(n608), .ZN(n370) );
  NOR2_X1 U480 ( .A1(n385), .A2(n696), .ZN(n371) );
  XNOR2_X1 U481 ( .A(n371), .B(KEYINPUT34), .ZN(n593) );
  XNOR2_X1 U482 ( .A(n416), .B(KEYINPUT39), .ZN(n539) );
  XNOR2_X1 U483 ( .A(n361), .B(n486), .ZN(n665) );
  XNOR2_X1 U484 ( .A(n485), .B(n766), .ZN(n486) );
  BUF_X1 U485 ( .A(n541), .Z(n551) );
  NAND2_X1 U486 ( .A1(n539), .A2(n685), .ZN(n540) );
  XOR2_X1 U487 ( .A(G137), .B(KEYINPUT71), .Z(n433) );
  XNOR2_X1 U488 ( .A(n767), .B(n396), .ZN(n734) );
  XNOR2_X1 U489 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U490 ( .A(n516), .B(n435), .ZN(n436) );
  AND2_X2 U491 ( .A1(n556), .A2(n592), .ZN(n682) );
  NAND2_X1 U492 ( .A1(n378), .A2(n379), .ZN(n373) );
  NAND2_X1 U493 ( .A1(n378), .A2(n379), .ZN(n511) );
  XNOR2_X1 U494 ( .A(n391), .B(n529), .ZN(n375) );
  XNOR2_X1 U495 ( .A(n391), .B(n529), .ZN(n550) );
  NOR2_X1 U496 ( .A1(n557), .A2(n682), .ZN(n558) );
  BUF_X1 U497 ( .A(n658), .Z(n376) );
  NAND2_X1 U498 ( .A1(n374), .A2(n431), .ZN(n378) );
  XNOR2_X1 U499 ( .A(n439), .B(n436), .ZN(n398) );
  XNOR2_X1 U500 ( .A(n400), .B(n364), .ZN(n566) );
  NOR2_X2 U501 ( .A1(n384), .A2(n362), .ZN(n581) );
  XNOR2_X2 U502 ( .A(n382), .B(n381), .ZN(n712) );
  NAND2_X1 U503 ( .A1(n413), .A2(n410), .ZN(n384) );
  NAND2_X1 U504 ( .A1(n413), .A2(n410), .ZN(n385) );
  NAND2_X1 U505 ( .A1(n510), .A2(n509), .ZN(n388) );
  NAND2_X1 U506 ( .A1(n386), .A2(n387), .ZN(n389) );
  NAND2_X1 U507 ( .A1(n389), .A2(n388), .ZN(n512) );
  INV_X1 U508 ( .A(n510), .ZN(n386) );
  INV_X1 U509 ( .A(n509), .ZN(n387) );
  XNOR2_X1 U510 ( .A(n390), .B(n518), .ZN(n658) );
  XNOR2_X1 U511 ( .A(n475), .B(n394), .ZN(n390) );
  NAND2_X2 U512 ( .A1(n527), .A2(n528), .ZN(n391) );
  NAND2_X1 U513 ( .A1(n392), .A2(n549), .ZN(n557) );
  NAND2_X1 U514 ( .A1(n548), .A2(n407), .ZN(n392) );
  XOR2_X1 U515 ( .A(n701), .B(KEYINPUT80), .Z(n619) );
  XNOR2_X1 U516 ( .A(n495), .B(n429), .ZN(n497) );
  NAND2_X1 U517 ( .A1(n595), .A2(n596), .ZN(n598) );
  NAND2_X1 U518 ( .A1(n360), .A2(n645), .ZN(n731) );
  XNOR2_X1 U519 ( .A(n395), .B(n474), .ZN(n394) );
  XNOR2_X1 U520 ( .A(n473), .B(n472), .ZN(n395) );
  XNOR2_X2 U521 ( .A(n511), .B(n432), .ZN(n475) );
  XNOR2_X2 U522 ( .A(n475), .B(n433), .ZN(n767) );
  NAND2_X1 U523 ( .A1(n573), .A2(KEYINPUT0), .ZN(n399) );
  NAND2_X1 U524 ( .A1(n664), .A2(n777), .ZN(n400) );
  XNOR2_X1 U525 ( .A(n537), .B(n536), .ZN(n777) );
  INV_X1 U526 ( .A(n701), .ZN(n406) );
  NAND2_X1 U527 ( .A1(n407), .A2(n689), .ZN(n680) );
  NAND2_X1 U528 ( .A1(n407), .A2(n685), .ZN(n684) );
  XNOR2_X1 U529 ( .A(n415), .B(KEYINPUT74), .ZN(n473) );
  INV_X1 U530 ( .A(n539), .ZN(n538) );
  NAND2_X1 U531 ( .A1(n375), .A2(n698), .ZN(n416) );
  XNOR2_X2 U532 ( .A(n489), .B(n488), .ZN(n554) );
  XNOR2_X1 U533 ( .A(n380), .B(G140), .ZN(n419) );
  NAND2_X1 U534 ( .A1(n425), .A2(n698), .ZN(n420) );
  XNOR2_X2 U535 ( .A(n530), .B(KEYINPUT38), .ZN(n698) );
  NAND2_X1 U536 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U537 ( .A1(n700), .A2(n426), .ZN(n425) );
  NOR2_X1 U538 ( .A1(n385), .A2(n428), .ZN(n616) );
  OR2_X1 U539 ( .A1(n615), .A2(n709), .ZN(n428) );
  XNOR2_X2 U540 ( .A(n581), .B(KEYINPUT22), .ZN(n621) );
  AND2_X1 U541 ( .A1(n599), .A2(n589), .ZN(n596) );
  INV_X2 U542 ( .A(n551), .ZN(n530) );
  XOR2_X1 U543 ( .A(n494), .B(n493), .Z(n429) );
  XOR2_X1 U544 ( .A(n651), .B(n650), .Z(n430) );
  NOR2_X1 U545 ( .A1(n476), .A2(n620), .ZN(n477) );
  XNOR2_X1 U546 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U547 ( .A(KEYINPUT30), .ZN(n525) );
  XNOR2_X1 U548 ( .A(n572), .B(n571), .ZN(n634) );
  INV_X1 U549 ( .A(n748), .ZN(n654) );
  XNOR2_X1 U550 ( .A(G134), .B(G131), .ZN(n432) );
  XNOR2_X1 U551 ( .A(n434), .B(G101), .ZN(n471) );
  XOR2_X2 U552 ( .A(G110), .B(G107), .Z(n516) );
  NAND2_X1 U553 ( .A1(G227), .A2(n403), .ZN(n438) );
  INV_X1 U554 ( .A(G140), .ZN(n437) );
  INV_X1 U555 ( .A(G902), .ZN(n440) );
  XNOR2_X2 U556 ( .A(n442), .B(G469), .ZN(n613) );
  XNOR2_X2 U557 ( .A(n613), .B(KEYINPUT1), .ZN(n706) );
  XOR2_X1 U558 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n445) );
  XNOR2_X1 U559 ( .A(n445), .B(n444), .ZN(n448) );
  XNOR2_X1 U560 ( .A(G119), .B(n372), .ZN(n447) );
  XNOR2_X1 U561 ( .A(G137), .B(KEYINPUT71), .ZN(n446) );
  NAND2_X1 U562 ( .A1(G221), .A2(n490), .ZN(n450) );
  NOR2_X1 U563 ( .A1(G902), .A2(n745), .ZN(n455) );
  NAND2_X1 U564 ( .A1(G234), .A2(n631), .ZN(n451) );
  XNOR2_X1 U565 ( .A(KEYINPUT20), .B(n451), .ZN(n463) );
  NAND2_X1 U566 ( .A1(G217), .A2(n463), .ZN(n453) );
  XNOR2_X1 U567 ( .A(KEYINPUT25), .B(KEYINPUT77), .ZN(n452) );
  XNOR2_X2 U568 ( .A(n455), .B(n454), .ZN(n710) );
  XOR2_X1 U569 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n457) );
  XNOR2_X1 U570 ( .A(n457), .B(n456), .ZN(n459) );
  NAND2_X1 U571 ( .A1(n459), .A2(G952), .ZN(n458) );
  XNOR2_X1 U572 ( .A(n458), .B(KEYINPUT90), .ZN(n724) );
  NOR2_X1 U573 ( .A1(n724), .A2(G953), .ZN(n578) );
  NAND2_X1 U574 ( .A1(G902), .A2(n459), .ZN(n574) );
  NOR2_X1 U575 ( .A1(G900), .A2(n574), .ZN(n460) );
  NAND2_X1 U576 ( .A1(G953), .A2(n460), .ZN(n461) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(n461), .Z(n462) );
  OR2_X1 U578 ( .A1(n578), .A2(n462), .ZN(n468) );
  NAND2_X1 U579 ( .A1(G221), .A2(n463), .ZN(n466) );
  INV_X1 U580 ( .A(KEYINPUT93), .ZN(n464) );
  XNOR2_X1 U581 ( .A(n464), .B(KEYINPUT21), .ZN(n465) );
  XNOR2_X1 U582 ( .A(n466), .B(n465), .ZN(n709) );
  INV_X1 U583 ( .A(n709), .ZN(n467) );
  AND2_X1 U584 ( .A1(n468), .A2(n467), .ZN(n523) );
  AND2_X1 U585 ( .A1(n710), .A2(n523), .ZN(n532) );
  INV_X1 U586 ( .A(n532), .ZN(n476) );
  XOR2_X1 U587 ( .A(KEYINPUT3), .B(G119), .Z(n470) );
  NAND2_X1 U588 ( .A1(n484), .A2(G210), .ZN(n474) );
  XNOR2_X1 U589 ( .A(n712), .B(KEYINPUT6), .ZN(n620) );
  XNOR2_X1 U590 ( .A(n477), .B(KEYINPUT107), .ZN(n499) );
  INV_X1 U591 ( .A(G122), .ZN(n478) );
  XNOR2_X1 U592 ( .A(n478), .B(G104), .ZN(n514) );
  XNOR2_X1 U593 ( .A(n514), .B(n479), .ZN(n483) );
  XOR2_X1 U594 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n481) );
  XNOR2_X1 U595 ( .A(G131), .B(KEYINPUT11), .ZN(n480) );
  XNOR2_X1 U596 ( .A(n481), .B(n480), .ZN(n482) );
  AND2_X1 U597 ( .A1(n484), .A2(G214), .ZN(n485) );
  NOR2_X1 U598 ( .A1(G902), .A2(n665), .ZN(n489) );
  XNOR2_X1 U599 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n487) );
  NAND2_X1 U600 ( .A1(n490), .A2(G217), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n374), .B(KEYINPUT100), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n492), .B(n491), .ZN(n495) );
  XNOR2_X1 U603 ( .A(G116), .B(G134), .ZN(n493) );
  XNOR2_X1 U604 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n496) );
  XNOR2_X1 U605 ( .A(n497), .B(n496), .ZN(n741) );
  NOR2_X2 U606 ( .A1(n499), .A2(n546), .ZN(n559) );
  NAND2_X1 U607 ( .A1(n440), .A2(n402), .ZN(n520) );
  NAND2_X1 U608 ( .A1(n559), .A2(n697), .ZN(n500) );
  XNOR2_X1 U609 ( .A(KEYINPUT108), .B(n500), .ZN(n501) );
  NOR2_X1 U610 ( .A1(n706), .A2(n501), .ZN(n503) );
  INV_X1 U611 ( .A(KEYINPUT43), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n503), .B(n502), .ZN(n522) );
  XNOR2_X1 U613 ( .A(n505), .B(n504), .ZN(n510) );
  NAND2_X1 U614 ( .A1(n506), .A2(G224), .ZN(n507) );
  XNOR2_X1 U615 ( .A(n512), .B(n373), .ZN(n517) );
  INV_X1 U616 ( .A(KEYINPUT16), .ZN(n513) );
  XNOR2_X1 U617 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U618 ( .A(n516), .B(n515), .ZN(n759) );
  XNOR2_X1 U619 ( .A(n517), .B(n759), .ZN(n519) );
  XNOR2_X1 U620 ( .A(n519), .B(n518), .ZN(n649) );
  NAND2_X1 U621 ( .A1(n649), .A2(n631), .ZN(n521) );
  XNOR2_X2 U622 ( .A(n521), .B(n363), .ZN(n541) );
  NAND2_X1 U623 ( .A1(n522), .A2(n530), .ZN(n639) );
  XNOR2_X1 U624 ( .A(n639), .B(G140), .ZN(G42) );
  NAND2_X1 U625 ( .A1(n523), .A2(n613), .ZN(n524) );
  NAND2_X1 U626 ( .A1(n712), .A2(n697), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U628 ( .A(KEYINPUT76), .ZN(n529) );
  AND2_X1 U629 ( .A1(n554), .A2(n367), .ZN(n689) );
  INV_X1 U630 ( .A(n689), .ZN(n545) );
  OR2_X1 U631 ( .A1(n538), .A2(n545), .ZN(n636) );
  XNOR2_X1 U632 ( .A(n636), .B(G134), .ZN(G36) );
  NAND2_X1 U633 ( .A1(n554), .A2(n553), .ZN(n700) );
  XNOR2_X1 U634 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n531) );
  NAND2_X1 U635 ( .A1(n532), .A2(n712), .ZN(n534) );
  XOR2_X1 U636 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n533) );
  XNOR2_X1 U637 ( .A(n534), .B(n533), .ZN(n535) );
  NAND2_X1 U638 ( .A1(n535), .A2(n613), .ZN(n544) );
  INV_X1 U639 ( .A(KEYINPUT42), .ZN(n536) );
  INV_X1 U640 ( .A(n546), .ZN(n685) );
  NAND2_X1 U641 ( .A1(n541), .A2(n697), .ZN(n542) );
  BUF_X1 U642 ( .A(n573), .Z(n543) );
  NAND2_X1 U643 ( .A1(n547), .A2(KEYINPUT47), .ZN(n549) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(n619), .ZN(n548) );
  NAND2_X1 U645 ( .A1(n550), .A2(n551), .ZN(n552) );
  XNOR2_X1 U646 ( .A(n552), .B(KEYINPUT109), .ZN(n556) );
  NOR2_X1 U647 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U648 ( .A(n555), .B(KEYINPUT105), .Z(n592) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT72), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n559), .B(KEYINPUT112), .ZN(n560) );
  AND2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U652 ( .A(n562), .B(KEYINPUT36), .ZN(n563) );
  XNOR2_X1 U653 ( .A(n706), .B(KEYINPUT86), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n563), .A2(n582), .ZN(n692) );
  AND2_X1 U655 ( .A1(n564), .A2(n692), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n566), .A2(n565), .ZN(n569) );
  INV_X1 U657 ( .A(KEYINPUT84), .ZN(n567) );
  XNOR2_X1 U658 ( .A(n567), .B(KEYINPUT48), .ZN(n568) );
  AND2_X1 U659 ( .A1(n639), .A2(n636), .ZN(n570) );
  NAND2_X1 U660 ( .A1(n641), .A2(n570), .ZN(n572) );
  INV_X1 U661 ( .A(KEYINPUT83), .ZN(n571) );
  NOR2_X1 U662 ( .A1(n634), .A2(n631), .ZN(n627) );
  INV_X1 U663 ( .A(n574), .ZN(n575) );
  NOR2_X1 U664 ( .A1(G898), .A2(n403), .ZN(n763) );
  NAND2_X1 U665 ( .A1(n575), .A2(n763), .ZN(n576) );
  XNOR2_X1 U666 ( .A(n576), .B(KEYINPUT91), .ZN(n577) );
  NOR2_X1 U667 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U668 ( .A(n579), .ZN(n580) );
  AND2_X1 U669 ( .A1(n582), .A2(n710), .ZN(n583) );
  AND2_X1 U670 ( .A1(n383), .A2(n583), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n621), .A2(n584), .ZN(n587) );
  INV_X1 U672 ( .A(KEYINPUT67), .ZN(n585) );
  XNOR2_X1 U673 ( .A(n585), .B(KEYINPUT32), .ZN(n586) );
  INV_X1 U674 ( .A(n712), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n710), .A2(n608), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n706), .A2(n588), .ZN(n600) );
  NAND2_X1 U677 ( .A1(n621), .A2(n600), .ZN(n589) );
  NOR2_X1 U678 ( .A1(n709), .A2(n710), .ZN(n707) );
  NAND2_X1 U679 ( .A1(n707), .A2(n706), .ZN(n609) );
  XNOR2_X1 U680 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT69), .ZN(n595) );
  INV_X1 U682 ( .A(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n607) );
  AND2_X1 U684 ( .A1(n621), .A2(n600), .ZN(n679) );
  INV_X1 U685 ( .A(KEYINPUT69), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n601), .A2(KEYINPUT44), .ZN(n602) );
  OR2_X1 U687 ( .A1(n679), .A2(n602), .ZN(n604) );
  NAND2_X1 U688 ( .A1(n670), .A2(n605), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n625) );
  OR2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n716) );
  NOR2_X1 U691 ( .A1(n384), .A2(n716), .ZN(n612) );
  XNOR2_X1 U692 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n610) );
  XNOR2_X1 U693 ( .A(n610), .B(KEYINPUT31), .ZN(n611) );
  XNOR2_X1 U694 ( .A(n612), .B(n611), .ZN(n688) );
  INV_X1 U695 ( .A(KEYINPUT95), .ZN(n617) );
  NOR2_X1 U696 ( .A1(n710), .A2(n370), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n617), .B(n616), .ZN(n674) );
  NOR2_X1 U699 ( .A1(n688), .A2(n674), .ZN(n618) );
  NOR2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT103), .ZN(n624) );
  XNOR2_X2 U702 ( .A(n626), .B(KEYINPUT45), .ZN(n749) );
  NAND2_X1 U703 ( .A1(n627), .A2(n749), .ZN(n630) );
  OR2_X1 U704 ( .A1(n631), .A2(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n628), .A2(KEYINPUT2), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n631), .A2(KEYINPUT82), .ZN(n632) );
  AND2_X2 U708 ( .A1(n633), .A2(n632), .ZN(n646) );
  INV_X1 U709 ( .A(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n771), .A2(n635), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n636), .A2(KEYINPUT2), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT79), .ZN(n638) );
  AND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  AND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n749), .A2(n642), .ZN(n643) );
  INV_X1 U716 ( .A(KEYINPUT66), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n356), .A2(G210), .ZN(n652) );
  BUF_X1 U718 ( .A(n649), .Z(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n652), .B(n430), .ZN(n655) );
  INV_X1 U721 ( .A(G952), .ZN(n653) );
  AND2_X2 U722 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U723 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U724 ( .A1(n744), .A2(G472), .ZN(n660) );
  XOR2_X1 U725 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n657) );
  XNOR2_X1 U726 ( .A(n376), .B(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X2 U728 ( .A1(n661), .A2(n748), .ZN(n663) );
  XNOR2_X1 U729 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(G57) );
  XNOR2_X1 U731 ( .A(n369), .B(G131), .ZN(G33) );
  NAND2_X1 U732 ( .A1(n744), .A2(G475), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X2 U734 ( .A1(n668), .A2(n748), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U736 ( .A(G119), .B(KEYINPUT127), .ZN(n671) );
  XOR2_X1 U737 ( .A(n671), .B(n670), .Z(G21) );
  XOR2_X1 U738 ( .A(G101), .B(n672), .Z(G3) );
  NAND2_X1 U739 ( .A1(n685), .A2(n674), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n673), .B(G104), .ZN(G6) );
  XNOR2_X1 U741 ( .A(G107), .B(KEYINPUT27), .ZN(n678) );
  XOR2_X1 U742 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n676) );
  NAND2_X1 U743 ( .A1(n674), .A2(n689), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U745 ( .A(n678), .B(n677), .ZN(G9) );
  XOR2_X1 U746 ( .A(G110), .B(n679), .Z(G12) );
  XOR2_X1 U747 ( .A(n372), .B(KEYINPUT29), .Z(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(n680), .ZN(G30) );
  XNOR2_X1 U749 ( .A(n682), .B(G143), .ZN(n683) );
  XNOR2_X1 U750 ( .A(n683), .B(KEYINPUT115), .ZN(G45) );
  XNOR2_X1 U751 ( .A(n684), .B(G146), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n688), .A2(n685), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n686), .B(KEYINPUT116), .ZN(n687) );
  XNOR2_X1 U754 ( .A(G113), .B(n687), .ZN(G15) );
  XOR2_X1 U755 ( .A(G116), .B(KEYINPUT117), .Z(n691) );
  NAND2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U757 ( .A(n691), .B(n690), .ZN(G18) );
  BUF_X1 U758 ( .A(n692), .Z(n694) );
  XOR2_X1 U759 ( .A(G125), .B(KEYINPUT37), .Z(n693) );
  XNOR2_X1 U760 ( .A(n694), .B(n693), .ZN(G27) );
  XNOR2_X1 U761 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n733) );
  NOR2_X1 U762 ( .A1(n749), .A2(KEYINPUT2), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U764 ( .A1(n700), .A2(n699), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n406), .A2(n702), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n696), .A2(n705), .ZN(n721) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U769 ( .A(KEYINPUT50), .B(n708), .Z(n715) );
  NAND2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U771 ( .A(n711), .B(KEYINPUT49), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n713), .A2(n370), .ZN(n714) );
  NAND2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U775 ( .A(KEYINPUT51), .B(n718), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n725), .A2(n719), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT52), .ZN(n723) );
  NOR2_X1 U779 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n696), .A2(n725), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U782 ( .A(KEYINPUT118), .B(n728), .Z(n729) );
  NOR2_X1 U783 ( .A1(G953), .A2(n729), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(G75) );
  XNOR2_X1 U786 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n737) );
  BUF_X1 U787 ( .A(n734), .Z(n735) );
  XNOR2_X1 U788 ( .A(n735), .B(KEYINPUT57), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n737), .B(n736), .ZN(n739) );
  NAND2_X1 U790 ( .A1(n356), .A2(G469), .ZN(n738) );
  XOR2_X1 U791 ( .A(n739), .B(n738), .Z(n740) );
  NOR2_X1 U792 ( .A1(n748), .A2(n740), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n356), .A2(G478), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n748), .A2(n743), .ZN(G63) );
  NAND2_X1 U796 ( .A1(n356), .A2(G217), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(G66) );
  INV_X1 U799 ( .A(n749), .ZN(n750) );
  NOR2_X1 U800 ( .A1(n750), .A2(G953), .ZN(n757) );
  XOR2_X1 U801 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n752) );
  NAND2_X1 U802 ( .A1(G224), .A2(G953), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U804 ( .A(KEYINPUT121), .B(n753), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n754), .A2(G898), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n755), .B(KEYINPUT123), .ZN(n756) );
  NOR2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n765) );
  XOR2_X1 U808 ( .A(G101), .B(KEYINPUT124), .Z(n758) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n760) );
  XOR2_X1 U810 ( .A(n761), .B(n760), .Z(n762) );
  NOR2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U812 ( .A(n765), .B(n764), .Z(G69) );
  XNOR2_X1 U813 ( .A(n767), .B(n766), .ZN(n772) );
  XOR2_X1 U814 ( .A(G227), .B(n772), .Z(n768) );
  NAND2_X1 U815 ( .A1(n768), .A2(G900), .ZN(n769) );
  XOR2_X1 U816 ( .A(KEYINPUT125), .B(n769), .Z(n770) );
  NAND2_X1 U817 ( .A1(G953), .A2(n770), .ZN(n775) );
  XOR2_X1 U818 ( .A(n771), .B(n772), .Z(n773) );
  NAND2_X1 U819 ( .A1(n773), .A2(n403), .ZN(n774) );
  NAND2_X1 U820 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U821 ( .A(n776), .B(KEYINPUT126), .ZN(G72) );
  XOR2_X1 U822 ( .A(n355), .B(G122), .Z(G24) );
  XNOR2_X1 U823 ( .A(G137), .B(n777), .ZN(G39) );
endmodule

