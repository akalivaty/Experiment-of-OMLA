//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .A4(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT65), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n194), .A2(new_n195), .A3(new_n191), .A4(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT66), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT66), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n197), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT11), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G134), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n209), .B2(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(KEYINPUT64), .A3(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n206), .A2(G137), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n209), .A2(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n188), .A2(new_n190), .A3(G128), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n188), .A2(new_n190), .B1(KEYINPUT0), .B2(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT0), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(G128), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n207), .A2(new_n210), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n214), .A2(new_n215), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n226), .A2(G131), .A3(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n206), .A2(KEYINPUT64), .A3(G137), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT64), .B1(new_n206), .B2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n212), .B1(new_n231), .B2(new_n211), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n224), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G116), .ZN(new_n235));
  INV_X1    g049(.A(G116), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G119), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n235), .B2(new_n237), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n237), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(new_n240), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n221), .A2(new_n233), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT71), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n228), .A2(new_n232), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n224), .A2(new_n225), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n193), .A2(new_n196), .B1(new_n202), .B2(new_n203), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n216), .A2(new_n219), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n248), .B1(new_n258), .B2(new_n247), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n249), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n251), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT29), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(G902), .B1(new_n262), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n221), .A2(new_n246), .A3(new_n233), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n246), .B1(new_n221), .B2(new_n233), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT28), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n250), .B1(new_n275), .B2(KEYINPUT68), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(KEYINPUT28), .C1(new_n273), .C2(new_n274), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n276), .A2(new_n277), .A3(new_n268), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n256), .A2(KEYINPUT30), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n221), .A2(new_n233), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n273), .B1(new_n285), .B2(new_n257), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n286), .B2(new_n268), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n221), .A2(new_n283), .A3(new_n233), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n283), .B1(new_n221), .B2(new_n233), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n257), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n247), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT70), .A3(new_n269), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n280), .A2(new_n270), .A3(new_n287), .A4(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n275), .A2(KEYINPUT68), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(new_n268), .A3(new_n279), .A4(new_n249), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n272), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G472), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n276), .A2(new_n279), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n268), .A3(new_n247), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n290), .A2(KEYINPUT31), .A3(new_n268), .A4(new_n247), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n269), .A2(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT32), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n303), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n249), .B1(new_n259), .B2(new_n278), .ZN(new_n309));
  INV_X1    g123(.A(new_n279), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n269), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(new_n305), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n298), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n298), .B2(new_n315), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT25), .ZN(new_n320));
  INV_X1    g134(.A(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT24), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G110), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(new_n324), .A3(KEYINPUT74), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT74), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n198), .A2(G119), .A3(new_n199), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  INV_X1    g143(.A(G128), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G119), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n199), .ZN(new_n338));
  NOR2_X1   g152(.A1(KEYINPUT66), .A2(G128), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(new_n234), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT73), .B1(new_n340), .B2(new_n331), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT75), .A3(new_n327), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n346));
  AND2_X1   g160(.A1(KEYINPUT76), .A2(G140), .ZN(new_n347));
  NOR2_X1   g161(.A1(KEYINPUT76), .A2(G140), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(G125), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  OR2_X1    g164(.A1(KEYINPUT76), .A2(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT76), .A2(G140), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT77), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n349), .B(KEYINPUT16), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(new_n350), .A2(G140), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT16), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G146), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n187), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n234), .B2(G128), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n332), .C1(new_n328), .C2(new_n364), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G110), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n345), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  OAI22_X1  g182(.A1(new_n343), .A2(new_n327), .B1(new_n366), .B2(G110), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n357), .A2(new_n354), .A3(new_n187), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n361), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G137), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n372), .B(new_n373), .Z(new_n374));
  AND3_X1   g188(.A1(new_n368), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n368), .B2(new_n371), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n375), .A2(new_n376), .A3(G902), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n319), .B(new_n320), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  INV_X1    g194(.A(G902), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(G234), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT25), .B1(new_n377), .B2(new_n319), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n368), .A2(new_n371), .ZN(new_n384));
  INV_X1    g198(.A(new_n374), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n368), .A2(new_n371), .A3(new_n374), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n381), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT79), .B1(new_n388), .B2(KEYINPUT78), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n379), .B(new_n382), .C1(new_n383), .C2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n382), .A2(G902), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n375), .A2(new_n376), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(KEYINPUT80), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(KEYINPUT80), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n317), .A2(new_n318), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n263), .A2(new_n264), .A3(G214), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(new_n189), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G131), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n399), .B(G143), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n212), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(KEYINPUT17), .A3(G131), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n405), .A2(new_n361), .A3(new_n362), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n400), .B(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n349), .B(G146), .C1(new_n353), .C2(new_n355), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n370), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G113), .B(G122), .ZN(new_n413));
  INV_X1    g227(.A(G104), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n407), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n349), .B(KEYINPUT19), .C1(new_n353), .C2(new_n355), .ZN(new_n417));
  OR2_X1    g231(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n357), .A2(new_n354), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n187), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n401), .A2(new_n403), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n361), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n415), .B1(new_n424), .B2(new_n412), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n398), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT20), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n416), .A2(new_n425), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n398), .ZN(new_n430));
  INV_X1    g244(.A(G475), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n415), .B1(new_n407), .B2(new_n412), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n381), .B1(new_n416), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n433), .B2(KEYINPUT94), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT94), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n381), .C1(new_n416), .C2(new_n432), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n427), .A2(new_n430), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n189), .A2(G128), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT13), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n198), .A2(G143), .A3(new_n199), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G134), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G122), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n236), .A2(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(G107), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n206), .A3(new_n438), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n443), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT81), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(new_n380), .A3(G953), .ZN(new_n453));
  INV_X1    g267(.A(G107), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n445), .B2(KEYINPUT14), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n447), .ZN(new_n457));
  INV_X1    g271(.A(new_n449), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n206), .B1(new_n441), .B2(new_n438), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n450), .A2(new_n453), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n453), .B1(new_n460), .B2(new_n450), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n381), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT95), .B(new_n381), .C1(new_n461), .C2(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n463), .A2(new_n467), .ZN(new_n470));
  INV_X1    g284(.A(G952), .ZN(new_n471));
  AOI211_X1 g285(.A(G953), .B(new_n471), .C1(G234), .C2(G237), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n381), .B(new_n264), .C1(G234), .C2(G237), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n469), .A2(new_n470), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT96), .B1(new_n437), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n430), .A2(new_n427), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n434), .A2(new_n436), .ZN(new_n480));
  AND4_X1   g294(.A1(KEYINPUT96), .A2(new_n479), .A3(new_n480), .A4(new_n477), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G221), .ZN(new_n483));
  INV_X1    g297(.A(new_n452), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n381), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n487));
  XNOR2_X1  g301(.A(G110), .B(G140), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n264), .A2(G227), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n252), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT3), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n414), .B2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n454), .A2(KEYINPUT3), .A3(G104), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G101), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT82), .B1(new_n454), .B2(G104), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n414), .A3(G107), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n496), .A2(new_n497), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n414), .B2(G107), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n414), .A2(G107), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n454), .A2(KEYINPUT84), .A3(G104), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G101), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n254), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n201), .A2(KEYINPUT85), .ZN(new_n511));
  OAI21_X1  g325(.A(G128), .B1(new_n201), .B2(KEYINPUT85), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n203), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n197), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n492), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n197), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n501), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n509), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT12), .A3(new_n492), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n498), .A2(new_n500), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n497), .B1(new_n525), .B2(new_n496), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT83), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G101), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT83), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT4), .A4(new_n501), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n253), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT4), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n534), .A3(G101), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n508), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n520), .A2(new_n537), .B1(new_n205), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n252), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n491), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n205), .A2(new_n519), .A3(KEYINPUT10), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n514), .B2(KEYINPUT10), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n535), .A2(new_n224), .A3(new_n225), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n527), .B2(new_n531), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n492), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n540), .A2(new_n491), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n487), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT12), .B1(new_n521), .B2(new_n492), .ZN(new_n549));
  AOI211_X1 g363(.A(new_n516), .B(new_n252), .C1(new_n520), .C2(new_n509), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n543), .A2(new_n545), .A3(new_n492), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n490), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n546), .A3(new_n491), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT86), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n548), .A2(G469), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G469), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n551), .A2(new_n552), .A3(new_n490), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n491), .B1(new_n540), .B2(new_n546), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n557), .B(new_n381), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(G469), .A2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n486), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n482), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G210), .B1(G237), .B2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G110), .B(G122), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT89), .B(KEYINPUT6), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT5), .B1(new_n239), .B2(new_n242), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT5), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n234), .A3(G116), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n574), .A2(G113), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n245), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n519), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n535), .B1(new_n243), .B2(new_n245), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n527), .B2(new_n531), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n577), .B1(new_n579), .B2(KEYINPUT87), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT87), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n581), .B(new_n578), .C1(new_n531), .C2(new_n527), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n570), .B(new_n571), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n254), .A2(new_n350), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n533), .B2(new_n350), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT90), .B(G224), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G953), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n586), .B(new_n588), .Z(new_n589));
  OAI21_X1  g403(.A(new_n570), .B1(new_n580), .B2(new_n582), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n527), .A2(new_n531), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n581), .B1(new_n591), .B2(new_n578), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n579), .A2(KEYINPUT87), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n569), .A3(new_n593), .A4(new_n577), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n594), .A3(KEYINPUT6), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT88), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT88), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n590), .A2(new_n594), .A3(new_n597), .A4(KEYINPUT6), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n584), .B(new_n589), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT7), .B1(new_n587), .B2(G953), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n586), .B(new_n600), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n569), .B(KEYINPUT8), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n575), .B1(new_n573), .B2(new_n244), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n519), .B(new_n603), .C1(new_n240), .C2(new_n244), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n604), .A2(KEYINPUT91), .B1(new_n519), .B2(new_n576), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n604), .A2(KEYINPUT91), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n594), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n381), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n609), .B1(new_n608), .B2(new_n381), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n568), .B1(new_n599), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n589), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT6), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n592), .A2(new_n593), .A3(new_n577), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n570), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n597), .B1(new_n618), .B2(new_n594), .ZN(new_n619));
  INV_X1    g433(.A(new_n598), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n583), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n608), .A2(new_n381), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT92), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n610), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n624), .A3(new_n567), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n566), .B1(new_n614), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n564), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n397), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  AND3_X1   g443(.A1(new_n621), .A2(new_n567), .A3(new_n624), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n567), .B1(new_n621), .B2(new_n624), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n565), .B(new_n476), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n461), .A2(new_n462), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT33), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n466), .A2(G902), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n465), .A2(new_n468), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT97), .B(G478), .Z(new_n637));
  AOI22_X1  g451(.A1(new_n634), .A2(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n437), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n308), .B2(new_n311), .ZN(new_n642));
  INV_X1    g456(.A(G472), .ZN(new_n643));
  OAI22_X1  g457(.A1(new_n642), .A2(new_n643), .B1(new_n304), .B2(new_n306), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n396), .A2(new_n563), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G104), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT98), .B(KEYINPUT34), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NOR2_X1   g463(.A1(new_n427), .A2(KEYINPUT99), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n436), .B2(new_n434), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n469), .A2(new_n470), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n430), .A2(KEYINPUT99), .A3(new_n427), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n645), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  NAND2_X1  g472(.A1(new_n564), .A2(new_n626), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n660));
  INV_X1    g474(.A(new_n382), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n319), .B1(new_n377), .B2(new_n378), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n320), .B1(new_n388), .B2(KEYINPUT79), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n385), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n384), .B(new_n665), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n664), .A2(new_n379), .B1(new_n391), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n660), .B1(new_n667), .B2(new_n644), .ZN(new_n668));
  INV_X1    g482(.A(new_n644), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n666), .A2(new_n391), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n390), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n669), .A2(KEYINPUT100), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n659), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT101), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G12));
  NOR2_X1   g491(.A1(new_n317), .A2(new_n318), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n473), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n472), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n651), .A2(new_n652), .A3(new_n653), .A4(new_n682), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n566), .B(new_n683), .C1(new_n614), .C2(new_n625), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n667), .A2(new_n563), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n678), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  INV_X1    g501(.A(new_n562), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n548), .A2(G469), .A3(new_n555), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n485), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n682), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT40), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n614), .A2(new_n625), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT38), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT38), .B1(new_n614), .B2(new_n625), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n286), .A2(new_n269), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n258), .A2(new_n269), .A3(new_n247), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n381), .ZN(new_n702));
  OAI21_X1  g516(.A(G472), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n315), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n652), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n437), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n667), .A2(new_n565), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n694), .A2(new_n699), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n189), .ZN(G45));
  NAND2_X1  g524(.A1(new_n479), .A2(new_n480), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n636), .A2(new_n637), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n633), .B(KEYINPUT33), .Z(new_n713));
  INV_X1    g527(.A(new_n635), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n715), .A3(new_n682), .ZN(new_n716));
  AOI211_X1 g530(.A(new_n566), .B(new_n716), .C1(new_n614), .C2(new_n625), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n313), .B1(new_n312), .B2(new_n305), .ZN(new_n718));
  AOI211_X1 g532(.A(KEYINPUT32), .B(new_n306), .C1(new_n308), .C2(new_n311), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT70), .B1(new_n291), .B2(new_n269), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n281), .B(new_n268), .C1(new_n290), .C2(new_n247), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n270), .A3(new_n724), .A4(new_n280), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n643), .B1(new_n725), .B2(new_n272), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT72), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n298), .A2(new_n315), .A3(new_n316), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n717), .A2(new_n727), .A3(new_n728), .A4(new_n685), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  NAND3_X1  g544(.A1(new_n626), .A2(new_n476), .A3(new_n639), .ZN(new_n731));
  INV_X1    g545(.A(new_n396), .ZN(new_n732));
  INV_X1    g546(.A(new_n560), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n523), .A2(new_n540), .A3(new_n491), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n540), .A2(new_n546), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n491), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n557), .B1(new_n736), .B2(new_n381), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n733), .A2(new_n737), .A3(new_n485), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n727), .A2(new_n732), .A3(new_n728), .A4(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT41), .B(G113), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND3_X1  g556(.A1(new_n397), .A2(new_n655), .A3(new_n738), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  INV_X1    g558(.A(new_n482), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n727), .A2(new_n745), .A3(new_n728), .A4(new_n671), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n626), .A2(new_n738), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n234), .ZN(G21));
  INV_X1    g563(.A(new_n642), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(G472), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n308), .B1(new_n268), .B2(new_n262), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n305), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n733), .A2(new_n737), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n486), .A3(new_n476), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n754), .A2(new_n756), .A3(new_n396), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n626), .A3(new_n706), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NOR3_X1   g573(.A1(new_n754), .A2(new_n667), .A3(new_n716), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n626), .A3(new_n738), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT102), .B(G125), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G27));
  NAND3_X1  g577(.A1(new_n614), .A2(new_n565), .A3(new_n625), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n561), .B(KEYINPUT103), .Z(new_n765));
  NAND2_X1  g579(.A1(new_n553), .A2(new_n554), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n560), .B(new_n765), .C1(new_n557), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n486), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n298), .A2(new_n315), .ZN(new_n771));
  INV_X1    g585(.A(new_n716), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n732), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n397), .A2(new_n769), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n212), .ZN(G33));
  INV_X1    g592(.A(new_n683), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n397), .A2(new_n779), .A3(new_n769), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  NAND2_X1  g595(.A1(new_n437), .A2(new_n715), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT43), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n671), .A2(new_n644), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT105), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n671), .A2(new_n644), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n764), .B1(new_n788), .B2(KEYINPUT44), .ZN(new_n789));
  INV_X1    g603(.A(new_n691), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n548), .B2(new_n555), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n766), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT46), .B(new_n765), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n560), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT46), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n765), .B1(new_n791), .B2(new_n793), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n795), .A2(KEYINPUT104), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT104), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n799), .A3(new_n560), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n485), .B(new_n790), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n783), .ZN(new_n802));
  INV_X1    g616(.A(new_n787), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n786), .B1(new_n671), .B2(new_n644), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n789), .A2(new_n801), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  XNOR2_X1  g623(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n795), .A2(KEYINPUT104), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n797), .A2(new_n796), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n812), .A2(new_n800), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n814), .B2(new_n485), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n798), .A2(new_n800), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n486), .A3(new_n810), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n772), .A2(new_n396), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n678), .A2(new_n764), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NOR4_X1   g635(.A1(new_n783), .A2(new_n396), .A3(new_n754), .A4(new_n681), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(G952), .B(new_n264), .C1(new_n823), .C2(new_n747), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n704), .A2(new_n732), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n738), .A2(new_n472), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n825), .A2(new_n764), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n824), .B1(new_n639), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n764), .A2(new_n783), .A3(new_n826), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n732), .A3(new_n771), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n737), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n566), .A3(new_n486), .A4(new_n560), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n697), .B2(new_n698), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n836), .B(KEYINPUT110), .C1(new_n697), .C2(new_n698), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT50), .B1(new_n841), .B2(new_n822), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n843), .B(new_n823), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n754), .A2(new_n667), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n829), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n829), .A2(new_n846), .A3(new_n847), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n827), .A2(new_n437), .A3(new_n638), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n815), .A2(new_n817), .B1(new_n485), .B2(new_n755), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n823), .A2(new_n764), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n851), .B(new_n852), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n845), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n829), .A2(new_n846), .A3(new_n847), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n852), .B1(new_n858), .B2(new_n848), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n815), .A2(new_n817), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n755), .A2(new_n485), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n862), .B2(new_n854), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n863), .B(new_n864), .C1(new_n842), .C2(new_n844), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n832), .B1(new_n857), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n727), .A2(new_n728), .A3(new_n685), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n651), .A2(new_n653), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n705), .A2(new_n682), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n764), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n868), .A2(new_n871), .B1(new_n760), .B2(new_n769), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n774), .A3(new_n776), .A4(new_n780), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n668), .A2(new_n672), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n627), .B1(new_n397), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n397), .A2(new_n641), .A3(new_n738), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n743), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n640), .B1(new_n711), .B2(new_n705), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n645), .A2(new_n878), .ZN(new_n879));
  OAI221_X1 g693(.A(new_n758), .B1(new_n879), .B2(new_n632), .C1(new_n747), .C2(new_n746), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n873), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n678), .B(new_n685), .C1(new_n684), .C2(new_n717), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n682), .B(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n767), .A2(new_n486), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n704), .A2(new_n671), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n626), .A3(new_n706), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n761), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT108), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n882), .A2(new_n886), .A3(KEYINPUT52), .A4(new_n761), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n887), .A2(KEYINPUT108), .A3(new_n888), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n881), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n877), .A2(new_n880), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n774), .A2(new_n776), .A3(new_n780), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n897), .A3(new_n872), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n889), .A2(new_n891), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(KEYINPUT54), .C1(new_n900), .C2(new_n893), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n893), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n881), .A2(new_n892), .A3(KEYINPUT53), .A4(new_n894), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n866), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n471), .A2(new_n264), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n755), .B(KEYINPUT49), .Z(new_n909));
  NAND4_X1  g723(.A1(new_n437), .A2(new_n715), .A3(new_n565), .A4(new_n486), .ZN(new_n910));
  OR4_X1    g724(.A1(new_n699), .A2(new_n825), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(KEYINPUT112), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n264), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n902), .A2(new_n904), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(G210), .A3(G902), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n583), .B1(new_n619), .B2(new_n620), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n615), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n924), .B(new_n925), .Z(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT115), .Z(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n922), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT114), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT114), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n922), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n931), .B2(new_n933), .ZN(G51));
  INV_X1    g748(.A(new_n905), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n903), .B1(new_n902), .B2(new_n904), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n765), .B(KEYINPUT57), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n736), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n791), .A2(new_n793), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT116), .Z(new_n941));
  NAND3_X1  g755(.A1(new_n919), .A2(G902), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n917), .B1(new_n939), .B2(new_n942), .ZN(G54));
  AND4_X1   g757(.A1(KEYINPUT58), .A2(new_n919), .A3(G475), .A4(G902), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n918), .B1(new_n944), .B2(new_n428), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n428), .B2(new_n944), .ZN(G60));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n947));
  INV_X1    g761(.A(new_n936), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n905), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n466), .A2(new_n381), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n713), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n947), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n947), .B(new_n953), .C1(new_n935), .C2(new_n936), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n901), .B2(new_n905), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n918), .B1(new_n957), .B2(new_n634), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n954), .A2(new_n956), .A3(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  NAND3_X1  g775(.A1(new_n919), .A2(new_n666), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n919), .A2(new_n961), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n393), .A2(new_n394), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n918), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT61), .B1(new_n962), .B2(KEYINPUT119), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G66));
  NOR2_X1   g781(.A1(new_n587), .A2(new_n474), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n264), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT120), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n877), .B2(new_n880), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n758), .B1(new_n746), .B2(new_n747), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n879), .A2(new_n632), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n727), .A2(new_n732), .A3(new_n728), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n659), .B1(new_n975), .B2(new_n673), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n740), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT120), .A4(new_n743), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n969), .B1(new_n979), .B2(new_n264), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n923), .B1(G898), .B2(new_n264), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT121), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n980), .B(new_n982), .ZN(G69));
  NAND2_X1  g797(.A1(G900), .A2(G953), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n285), .B(new_n421), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n732), .A2(new_n626), .A3(new_n771), .A4(new_n706), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n486), .A3(new_n816), .A4(new_n691), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n774), .A2(new_n987), .A3(new_n776), .A4(new_n780), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n626), .A2(new_n779), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n626), .A2(new_n772), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n867), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n761), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT123), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT123), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n686), .A2(new_n729), .A3(new_n994), .A4(new_n761), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n988), .A2(new_n808), .A3(new_n820), .A4(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n984), .B(new_n985), .C1(new_n997), .C2(G953), .ZN(new_n998));
  INV_X1    g812(.A(new_n692), .ZN(new_n999));
  INV_X1    g813(.A(new_n764), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n397), .A2(new_n999), .A3(new_n1000), .A4(new_n878), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n820), .A2(new_n808), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n709), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT123), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n994), .B1(new_n882), .B2(new_n761), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1002), .B1(new_n1006), .B2(KEYINPUT62), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  AND4_X1   g822(.A1(KEYINPUT124), .A2(new_n996), .A3(new_n1008), .A4(new_n1003), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n709), .B1(new_n993), .B2(new_n995), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT124), .B1(new_n1010), .B2(new_n1008), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1007), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1012), .A2(new_n264), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n985), .B(KEYINPUT122), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n998), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n997), .B2(new_n979), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1020), .A2(new_n269), .A3(new_n286), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1019), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n723), .B2(new_n300), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n895), .B(new_n1023), .C1(new_n900), .C2(new_n893), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1021), .A2(new_n1024), .A3(new_n918), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT125), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n971), .A2(new_n978), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1007), .B(new_n1027), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1019), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1026), .B1(new_n1029), .B2(new_n700), .ZN(new_n1030));
  INV_X1    g844(.A(new_n700), .ZN(new_n1031));
  AOI211_X1 g845(.A(KEYINPUT125), .B(new_n1031), .C1(new_n1028), .C2(new_n1019), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1025), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT126), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n1025), .B(KEYINPUT126), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(G57));
endmodule


