

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U549 ( .A1(G8), .A2(n741), .ZN(n793) );
  NOR2_X1 U550 ( .A1(n635), .A2(n527), .ZN(n640) );
  NAND2_X2 U551 ( .A1(n709), .A2(n708), .ZN(n741) );
  NOR2_X2 U552 ( .A1(G2104), .A2(n517), .ZN(n871) );
  XNOR2_X1 U553 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n514) );
  OR2_X1 U554 ( .A1(n721), .A2(n720), .ZN(n718) );
  INV_X1 U555 ( .A(n914), .ZN(n775) );
  NAND2_X1 U556 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U557 ( .A1(G1966), .A2(n793), .ZN(n767) );
  XNOR2_X1 U558 ( .A(n762), .B(n514), .ZN(n769) );
  NOR2_X1 U559 ( .A1(n769), .A2(n768), .ZN(n778) );
  AND2_X1 U560 ( .A1(G160), .A2(G40), .ZN(n709) );
  INV_X1 U561 ( .A(KEYINPUT105), .ZN(n798) );
  NOR2_X1 U562 ( .A1(n635), .A2(G651), .ZN(n638) );
  NOR2_X1 U563 ( .A1(n591), .A2(n590), .ZN(n593) );
  NOR2_X1 U564 ( .A1(n525), .A2(n524), .ZN(G160) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n516) );
  INV_X1 U566 ( .A(G2105), .ZN(n517) );
  AND2_X2 U567 ( .A1(n517), .A2(G2104), .ZN(n875) );
  NAND2_X1 U568 ( .A1(G101), .A2(n875), .ZN(n515) );
  XNOR2_X1 U569 ( .A(n516), .B(n515), .ZN(n520) );
  NAND2_X1 U570 ( .A1(G125), .A2(n871), .ZN(n518) );
  XOR2_X1 U571 ( .A(KEYINPUT65), .B(n518), .Z(n519) );
  NAND2_X1 U572 ( .A1(n520), .A2(n519), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U574 ( .A(KEYINPUT17), .B(n521), .Z(n876) );
  NAND2_X1 U575 ( .A1(G137), .A2(n876), .ZN(n523) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U577 ( .A1(G113), .A2(n872), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  INV_X1 U579 ( .A(G651), .ZN(n527) );
  NOR2_X1 U580 ( .A1(G543), .A2(n527), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n526), .Z(n639) );
  NAND2_X1 U582 ( .A1(G65), .A2(n639), .ZN(n529) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  NAND2_X1 U584 ( .A1(G78), .A2(n640), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n638), .A2(G53), .ZN(n532) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n530) );
  XNOR2_X1 U588 ( .A(n530), .B(KEYINPUT64), .ZN(n643) );
  NAND2_X1 U589 ( .A1(G91), .A2(n643), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(G299) );
  NAND2_X1 U592 ( .A1(G72), .A2(n640), .ZN(n536) );
  NAND2_X1 U593 ( .A1(G85), .A2(n643), .ZN(n535) );
  NAND2_X1 U594 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G60), .A2(n639), .ZN(n538) );
  NAND2_X1 U596 ( .A1(G47), .A2(n638), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U598 ( .A1(n540), .A2(n539), .ZN(G290) );
  NAND2_X1 U599 ( .A1(G64), .A2(n639), .ZN(n542) );
  NAND2_X1 U600 ( .A1(G52), .A2(n638), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U602 ( .A(KEYINPUT67), .B(n543), .Z(n548) );
  NAND2_X1 U603 ( .A1(G77), .A2(n640), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G90), .A2(n643), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(G171) );
  NAND2_X1 U608 ( .A1(G99), .A2(n875), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n549), .B(KEYINPUT82), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G123), .A2(n871), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT18), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n551), .B(KEYINPUT80), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G135), .A2(n876), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n553), .A2(n552), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G111), .A2(n872), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT81), .B(n554), .ZN(n555) );
  NOR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n937) );
  XNOR2_X1 U619 ( .A(G2096), .B(n937), .ZN(n559) );
  OR2_X1 U620 ( .A1(G2100), .A2(n559), .ZN(G156) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G132), .ZN(G219) );
  NAND2_X1 U623 ( .A1(G102), .A2(n875), .ZN(n561) );
  NAND2_X1 U624 ( .A1(G138), .A2(n876), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G126), .A2(n871), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G114), .A2(n872), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n565), .A2(n564), .ZN(G164) );
  NAND2_X1 U630 ( .A1(n643), .A2(G89), .ZN(n566) );
  XOR2_X1 U631 ( .A(KEYINPUT75), .B(n566), .Z(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G76), .A2(n640), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT5), .ZN(n577) );
  XNOR2_X1 U636 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n639), .A2(G63), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT76), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G51), .A2(n638), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G94), .A2(G452), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT68), .B(n579), .Z(G173) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U649 ( .A(G223), .B(KEYINPUT70), .Z(n816) );
  NAND2_X1 U650 ( .A1(n816), .A2(G567), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n581), .Z(G234) );
  NAND2_X1 U652 ( .A1(n639), .A2(G56), .ZN(n582) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n582), .Z(n591) );
  NAND2_X1 U654 ( .A1(n640), .A2(G68), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n583), .B(KEYINPUT72), .ZN(n587) );
  XOR2_X1 U656 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n585) );
  NAND2_X1 U657 ( .A1(G81), .A2(n643), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n585), .B(n584), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U660 ( .A(KEYINPUT13), .B(n588), .ZN(n589) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n589), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n638), .A2(G43), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n921) );
  INV_X1 U664 ( .A(G860), .ZN(n606) );
  OR2_X1 U665 ( .A1(n921), .A2(n606), .ZN(G153) );
  INV_X1 U666 ( .A(G171), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G54), .A2(n638), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G66), .A2(n639), .ZN(n595) );
  NAND2_X1 U670 ( .A1(G79), .A2(n640), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n643), .A2(G92), .ZN(n596) );
  XOR2_X1 U673 ( .A(KEYINPUT74), .B(n596), .Z(n597) );
  NOR2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n601), .B(KEYINPUT15), .ZN(n720) );
  INV_X1 U677 ( .A(n720), .ZN(n908) );
  INV_X1 U678 ( .A(G868), .ZN(n658) );
  NAND2_X1 U679 ( .A1(n908), .A2(n658), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U682 ( .A1(G286), .A2(n658), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n607), .A2(n720), .ZN(n608) );
  XNOR2_X1 U686 ( .A(n608), .B(KEYINPUT78), .ZN(n609) );
  XNOR2_X1 U687 ( .A(KEYINPUT16), .B(n609), .ZN(G148) );
  NOR2_X1 U688 ( .A1(G559), .A2(n658), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n720), .A2(n610), .ZN(n611) );
  XNOR2_X1 U690 ( .A(n611), .B(KEYINPUT79), .ZN(n613) );
  NOR2_X1 U691 ( .A1(n921), .A2(G868), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G80), .A2(n640), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G93), .A2(n643), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U696 ( .A(KEYINPUT84), .B(n616), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G67), .A2(n639), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G55), .A2(n638), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n659) );
  NAND2_X1 U701 ( .A1(n720), .A2(G559), .ZN(n656) );
  XOR2_X1 U702 ( .A(KEYINPUT83), .B(n921), .Z(n621) );
  XNOR2_X1 U703 ( .A(n656), .B(n621), .ZN(n622) );
  NOR2_X1 U704 ( .A1(G860), .A2(n622), .ZN(n623) );
  XOR2_X1 U705 ( .A(n659), .B(n623), .Z(G145) );
  NAND2_X1 U706 ( .A1(G61), .A2(n639), .ZN(n625) );
  NAND2_X1 U707 ( .A1(G86), .A2(n643), .ZN(n624) );
  NAND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n640), .A2(G73), .ZN(n626) );
  XOR2_X1 U710 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n638), .A2(G48), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G49), .A2(n638), .ZN(n632) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U716 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U717 ( .A1(n639), .A2(n633), .ZN(n634) );
  XOR2_X1 U718 ( .A(KEYINPUT85), .B(n634), .Z(n637) );
  NAND2_X1 U719 ( .A1(n635), .A2(G87), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G50), .A2(n638), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G62), .A2(n639), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G75), .A2(n640), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n643), .A2(G88), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT86), .B(n644), .Z(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U728 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(KEYINPUT87), .ZN(G166) );
  XOR2_X1 U730 ( .A(G290), .B(G305), .Z(n650) );
  XNOR2_X1 U731 ( .A(n921), .B(n650), .ZN(n653) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(G299), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n651), .B(G288), .ZN(n652) );
  XOR2_X1 U734 ( .A(n653), .B(n652), .Z(n655) );
  XOR2_X1 U735 ( .A(G166), .B(n659), .Z(n654) );
  XNOR2_X1 U736 ( .A(n655), .B(n654), .ZN(n888) );
  XOR2_X1 U737 ( .A(n888), .B(n656), .Z(n657) );
  NAND2_X1 U738 ( .A1(G868), .A2(n657), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U747 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U748 ( .A1(G219), .A2(G220), .ZN(n667) );
  XNOR2_X1 U749 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n668), .A2(G96), .ZN(n669) );
  NOR2_X1 U752 ( .A1(G218), .A2(n669), .ZN(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT89), .B(n670), .ZN(n822) );
  NAND2_X1 U754 ( .A1(n822), .A2(G2106), .ZN(n675) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n672), .A2(G108), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n673), .B(KEYINPUT90), .ZN(n823) );
  NAND2_X1 U759 ( .A1(G567), .A2(n823), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n824) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U762 ( .A1(n824), .A2(n676), .ZN(n819) );
  NAND2_X1 U763 ( .A1(n819), .A2(G36), .ZN(G176) );
  XNOR2_X1 U764 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n708) );
  NAND2_X1 U766 ( .A1(G160), .A2(G40), .ZN(n677) );
  NOR2_X1 U767 ( .A1(n708), .A2(n677), .ZN(n811) );
  XNOR2_X1 U768 ( .A(G2067), .B(KEYINPUT37), .ZN(n809) );
  NAND2_X1 U769 ( .A1(G104), .A2(n875), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G140), .A2(n876), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U772 ( .A(KEYINPUT34), .B(n680), .ZN(n686) );
  NAND2_X1 U773 ( .A1(G128), .A2(n871), .ZN(n682) );
  NAND2_X1 U774 ( .A1(G116), .A2(n872), .ZN(n681) );
  NAND2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U776 ( .A(KEYINPUT35), .B(n683), .Z(n684) );
  XNOR2_X1 U777 ( .A(KEYINPUT92), .B(n684), .ZN(n685) );
  NOR2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U779 ( .A(KEYINPUT36), .B(n687), .ZN(n866) );
  NOR2_X1 U780 ( .A1(n809), .A2(n866), .ZN(n948) );
  NAND2_X1 U781 ( .A1(n811), .A2(n948), .ZN(n807) );
  NAND2_X1 U782 ( .A1(G129), .A2(n871), .ZN(n689) );
  NAND2_X1 U783 ( .A1(G117), .A2(n872), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n875), .A2(G105), .ZN(n690) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(n690), .Z(n691) );
  NOR2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U788 ( .A(KEYINPUT93), .B(n693), .Z(n695) );
  NAND2_X1 U789 ( .A1(n876), .A2(G141), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n862) );
  AND2_X1 U791 ( .A1(n862), .A2(G1996), .ZN(n703) );
  NAND2_X1 U792 ( .A1(G95), .A2(n875), .ZN(n697) );
  NAND2_X1 U793 ( .A1(G131), .A2(n876), .ZN(n696) );
  NAND2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U795 ( .A1(G119), .A2(n871), .ZN(n699) );
  NAND2_X1 U796 ( .A1(G107), .A2(n872), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U798 ( .A1(n701), .A2(n700), .ZN(n884) );
  INV_X1 U799 ( .A(G1991), .ZN(n992) );
  NOR2_X1 U800 ( .A1(n884), .A2(n992), .ZN(n702) );
  NOR2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n933) );
  INV_X1 U802 ( .A(n811), .ZN(n704) );
  NOR2_X1 U803 ( .A1(n933), .A2(n704), .ZN(n804) );
  INV_X1 U804 ( .A(n804), .ZN(n705) );
  NAND2_X1 U805 ( .A1(n807), .A2(n705), .ZN(n797) );
  NOR2_X1 U806 ( .A1(G2090), .A2(G303), .ZN(n706) );
  XOR2_X1 U807 ( .A(KEYINPUT103), .B(n706), .Z(n707) );
  NAND2_X1 U808 ( .A1(G8), .A2(n707), .ZN(n771) );
  INV_X1 U809 ( .A(G1996), .ZN(n987) );
  NOR2_X1 U810 ( .A1(n741), .A2(n987), .ZN(n711) );
  INV_X1 U811 ( .A(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U812 ( .A(n711), .B(n710), .ZN(n713) );
  BUF_X1 U813 ( .A(n741), .Z(n753) );
  NAND2_X1 U814 ( .A1(n753), .A2(G1341), .ZN(n712) );
  NAND2_X1 U815 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U816 ( .A1(n921), .A2(n714), .ZN(n719) );
  NAND2_X1 U817 ( .A1(G1348), .A2(n741), .ZN(n716) );
  INV_X1 U818 ( .A(n741), .ZN(n724) );
  NAND2_X1 U819 ( .A1(G2067), .A2(n724), .ZN(n715) );
  NAND2_X1 U820 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U821 ( .A(KEYINPUT97), .B(n717), .ZN(n721) );
  NAND2_X1 U822 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U823 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n724), .A2(G2072), .ZN(n726) );
  INV_X1 U826 ( .A(KEYINPUT27), .ZN(n725) );
  XNOR2_X1 U827 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U828 ( .A1(G1956), .A2(n753), .ZN(n727) );
  NAND2_X1 U829 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U830 ( .A1(G299), .A2(n731), .ZN(n729) );
  NOR2_X1 U831 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U832 ( .A1(G299), .A2(n731), .ZN(n732) );
  XOR2_X1 U833 ( .A(KEYINPUT28), .B(n732), .Z(n733) );
  NOR2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U835 ( .A(n735), .B(KEYINPUT29), .ZN(n740) );
  XNOR2_X1 U836 ( .A(KEYINPUT25), .B(G2078), .ZN(n995) );
  NAND2_X1 U837 ( .A1(n724), .A2(n995), .ZN(n736) );
  XNOR2_X1 U838 ( .A(n736), .B(KEYINPUT96), .ZN(n738) );
  XNOR2_X1 U839 ( .A(G1961), .B(KEYINPUT95), .ZN(n962) );
  NAND2_X1 U840 ( .A1(n962), .A2(n753), .ZN(n737) );
  NAND2_X1 U841 ( .A1(n738), .A2(n737), .ZN(n746) );
  NAND2_X1 U842 ( .A1(G171), .A2(n746), .ZN(n739) );
  NAND2_X1 U843 ( .A1(n740), .A2(n739), .ZN(n752) );
  NOR2_X1 U844 ( .A1(G2084), .A2(n741), .ZN(n763) );
  NOR2_X1 U845 ( .A1(n767), .A2(n763), .ZN(n742) );
  NAND2_X1 U846 ( .A1(G8), .A2(n742), .ZN(n743) );
  XNOR2_X1 U847 ( .A(n743), .B(KEYINPUT30), .ZN(n744) );
  NOR2_X1 U848 ( .A1(n744), .A2(G168), .ZN(n745) );
  XNOR2_X1 U849 ( .A(n745), .B(KEYINPUT98), .ZN(n748) );
  NOR2_X1 U850 ( .A1(n746), .A2(G171), .ZN(n747) );
  NOR2_X1 U851 ( .A1(n748), .A2(n747), .ZN(n750) );
  INV_X1 U852 ( .A(KEYINPUT31), .ZN(n749) );
  XNOR2_X1 U853 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U854 ( .A1(n752), .A2(n751), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(G286), .ZN(n761) );
  INV_X1 U856 ( .A(G8), .ZN(n759) );
  NOR2_X1 U857 ( .A1(G1971), .A2(n793), .ZN(n755) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n753), .ZN(n754) );
  NOR2_X1 U859 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U860 ( .A(KEYINPUT99), .B(n756), .Z(n757) );
  NAND2_X1 U861 ( .A1(n757), .A2(G303), .ZN(n758) );
  OR2_X1 U862 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U863 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U864 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U865 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U866 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U867 ( .A(n778), .ZN(n770) );
  NAND2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U869 ( .A1(n772), .A2(n793), .ZN(n773) );
  XNOR2_X1 U870 ( .A(KEYINPUT104), .B(n773), .ZN(n789) );
  NOR2_X1 U871 ( .A1(G1971), .A2(G303), .ZN(n774) );
  XNOR2_X1 U872 ( .A(n774), .B(KEYINPUT101), .ZN(n776) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n914) );
  OR2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U875 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U876 ( .A(n915), .ZN(n779) );
  NOR2_X1 U877 ( .A1(n793), .A2(n779), .ZN(n780) );
  AND2_X1 U878 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U879 ( .A1(n782), .A2(KEYINPUT33), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n914), .A2(KEYINPUT33), .ZN(n783) );
  NOR2_X1 U881 ( .A1(n783), .A2(n793), .ZN(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U883 ( .A(G1981), .B(G305), .Z(n924) );
  NAND2_X1 U884 ( .A1(n786), .A2(n924), .ZN(n787) );
  XNOR2_X1 U885 ( .A(n787), .B(KEYINPUT102), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n795) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U888 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  XNOR2_X1 U889 ( .A(KEYINPUT94), .B(n791), .ZN(n792) );
  NOR2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n799) );
  XNOR2_X1 U893 ( .A(n799), .B(n798), .ZN(n801) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n918) );
  NAND2_X1 U895 ( .A1(n918), .A2(n811), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n814) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n862), .ZN(n940) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n802) );
  AND2_X1 U899 ( .A1(n992), .A2(n884), .ZN(n936) );
  NOR2_X1 U900 ( .A1(n802), .A2(n936), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n940), .A2(n805), .ZN(n806) );
  XNOR2_X1 U903 ( .A(n806), .B(KEYINPUT39), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n809), .A2(n866), .ZN(n945) );
  NAND2_X1 U906 ( .A1(n810), .A2(n945), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(KEYINPUT40), .B(n815), .ZN(G329) );
  NAND2_X1 U910 ( .A1(n816), .A2(G2106), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U913 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT107), .B(n821), .Z(G188) );
  XOR2_X1 U917 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(G325) );
  XNOR2_X1 U919 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(n824), .ZN(G319) );
  XOR2_X1 U924 ( .A(G2100), .B(G2096), .Z(n826) );
  XNOR2_X1 U925 ( .A(KEYINPUT42), .B(G2678), .ZN(n825) );
  XNOR2_X1 U926 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U927 ( .A(KEYINPUT43), .B(G2072), .Z(n828) );
  XNOR2_X1 U928 ( .A(G2067), .B(G2090), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U930 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U931 ( .A(G2078), .B(G2084), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U933 ( .A(G1976), .B(G1966), .Z(n834) );
  XNOR2_X1 U934 ( .A(G1961), .B(G1956), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n844) );
  XOR2_X1 U936 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n836) );
  XNOR2_X1 U937 ( .A(G1996), .B(KEYINPUT112), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U939 ( .A(G1971), .B(G1981), .Z(n838) );
  XNOR2_X1 U940 ( .A(G1991), .B(G1986), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U942 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U943 ( .A(KEYINPUT111), .B(G2474), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G100), .A2(n875), .ZN(n846) );
  NAND2_X1 U947 ( .A1(G112), .A2(n872), .ZN(n845) );
  NAND2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n871), .A2(G124), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U951 ( .A1(G136), .A2(n876), .ZN(n848) );
  NAND2_X1 U952 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(KEYINPUT113), .B(n850), .Z(n851) );
  NOR2_X1 U954 ( .A1(n852), .A2(n851), .ZN(G162) );
  NAND2_X1 U955 ( .A1(n871), .A2(G127), .ZN(n853) );
  XOR2_X1 U956 ( .A(KEYINPUT115), .B(n853), .Z(n855) );
  NAND2_X1 U957 ( .A1(n872), .A2(G115), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n856), .B(KEYINPUT47), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G139), .A2(n876), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n875), .A2(G103), .ZN(n859) );
  XOR2_X1 U963 ( .A(KEYINPUT114), .B(n859), .Z(n860) );
  NOR2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n950) );
  XNOR2_X1 U965 ( .A(n950), .B(G162), .ZN(n870) );
  XOR2_X1 U966 ( .A(KEYINPUT46), .B(KEYINPUT116), .Z(n864) );
  XOR2_X1 U967 ( .A(n862), .B(KEYINPUT48), .Z(n863) );
  XNOR2_X1 U968 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n868) );
  XNOR2_X1 U970 ( .A(G164), .B(G160), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n886) );
  NAND2_X1 U973 ( .A1(G130), .A2(n871), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G118), .A2(n872), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n881) );
  NAND2_X1 U976 ( .A1(G106), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G142), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n879), .B(KEYINPUT45), .Z(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(n937), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U984 ( .A1(G37), .A2(n887), .ZN(G395) );
  XNOR2_X1 U985 ( .A(n888), .B(n908), .ZN(n890) );
  XOR2_X1 U986 ( .A(G171), .B(G286), .Z(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U988 ( .A1(G37), .A2(n891), .ZN(G397) );
  XOR2_X1 U989 ( .A(G2451), .B(G2430), .Z(n893) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2443), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n899) );
  XOR2_X1 U992 ( .A(G2435), .B(G2454), .Z(n895) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U995 ( .A(G2446), .B(G2427), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U998 ( .A1(G14), .A2(n900), .ZN(n907) );
  NAND2_X1 U999 ( .A1(G319), .A2(n907), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n901) );
  XOR2_X1 U1001 ( .A(KEYINPUT117), .B(n901), .Z(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(KEYINPUT49), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G108), .ZN(G238) );
  INV_X1 U1008 ( .A(n907), .ZN(G401) );
  XOR2_X1 U1009 ( .A(KEYINPUT56), .B(G16), .Z(n932) );
  XOR2_X1 U1010 ( .A(G303), .B(G1971), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G301), .B(G1961), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n908), .B(G1348), .ZN(n909) );
  NOR2_X1 U1013 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1014 ( .A(KEYINPUT124), .B(n911), .ZN(n912) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n930) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n775), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT125), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G1956), .B(G299), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(G1341), .B(n921), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(G168), .B(G1966), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT57), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n1014) );
  XNOR2_X1 U1029 ( .A(KEYINPUT52), .B(KEYINPUT121), .ZN(n958) );
  XNOR2_X1 U1030 ( .A(G160), .B(G2084), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n944) );
  XOR2_X1 U1034 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT51), .B(n941), .Z(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT118), .B(n942), .Z(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT119), .B(n949), .Z(n956) );
  XOR2_X1 U1042 ( .A(G2072), .B(n950), .Z(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT120), .B(n951), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n954), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(n958), .B(n957), .ZN(n960) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1051 ( .A1(n961), .A2(G29), .ZN(n1012) );
  XNOR2_X1 U1052 ( .A(G5), .B(n962), .ZN(n975) );
  XOR2_X1 U1053 ( .A(G1956), .B(G20), .Z(n967) );
  XNOR2_X1 U1054 ( .A(G1981), .B(G6), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G1341), .B(G19), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(KEYINPUT126), .B(n965), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n970) );
  XOR2_X1 U1059 ( .A(KEYINPUT59), .B(G1348), .Z(n968) );
  XNOR2_X1 U1060 ( .A(G4), .B(n968), .ZN(n969) );
  NOR2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(KEYINPUT60), .B(n971), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n982) );
  XNOR2_X1 U1066 ( .A(G1971), .B(G22), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G23), .B(G1976), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G1986), .B(G24), .Z(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT58), .B(n980), .ZN(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(KEYINPUT61), .B(n983), .ZN(n985) );
  INV_X1 U1074 ( .A(G16), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n986), .A2(G11), .ZN(n1010) );
  XOR2_X1 U1077 ( .A(G2067), .B(G26), .Z(n989) );
  XNOR2_X1 U1078 ( .A(n987), .B(G32), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G33), .B(G2072), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(n992), .B(G25), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n993), .A2(G28), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT122), .ZN(n997) );
  XOR2_X1 U1085 ( .A(G27), .B(n995), .Z(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT53), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(G2084), .B(G34), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(KEYINPUT54), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G35), .B(G2090), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT55), .B(n1006), .Z(n1007) );
  NOR2_X1 U1095 ( .A1(G29), .A2(n1007), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(KEYINPUT123), .B(n1008), .Z(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT127), .B(n1015), .Z(n1016) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1016), .ZN(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

