

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766;

  NOR2_X1 U375 ( .A1(G953), .A2(n732), .ZN(n733) );
  AND2_X1 U376 ( .A1(n424), .A2(n423), .ZN(n637) );
  OR2_X1 U377 ( .A1(n647), .A2(n717), .ZN(n648) );
  NOR2_X1 U378 ( .A1(n647), .A2(n629), .ZN(n375) );
  NOR2_X1 U379 ( .A1(n625), .A2(n624), .ZN(n627) );
  XNOR2_X1 U380 ( .A(n623), .B(KEYINPUT1), .ZN(n708) );
  XNOR2_X1 U381 ( .A(n493), .B(n492), .ZN(n665) );
  XNOR2_X1 U382 ( .A(n422), .B(G143), .ZN(n526) );
  XNOR2_X2 U383 ( .A(n352), .B(n524), .ZN(n611) );
  XNOR2_X2 U384 ( .A(G110), .B(G107), .ZN(n449) );
  AND2_X2 U385 ( .A1(n687), .A2(KEYINPUT2), .ZN(n654) );
  XNOR2_X2 U386 ( .A(n523), .B(n522), .ZN(n352) );
  XNOR2_X2 U387 ( .A(n448), .B(G101), .ZN(n450) );
  INV_X1 U388 ( .A(G953), .ZN(n752) );
  INV_X2 U389 ( .A(G104), .ZN(n448) );
  XOR2_X2 U390 ( .A(KEYINPUT10), .B(n527), .Z(n748) );
  NOR2_X1 U391 ( .A1(n766), .A2(n764), .ZN(n650) );
  NOR2_X1 U392 ( .A1(n762), .A2(n571), .ZN(n600) );
  NAND2_X2 U393 ( .A1(n442), .A2(n439), .ZN(n706) );
  AND2_X1 U394 ( .A1(n381), .A2(n380), .ZN(n379) );
  AND2_X1 U395 ( .A1(n765), .A2(n590), .ZN(n380) );
  XNOR2_X1 U396 ( .A(n596), .B(KEYINPUT102), .ZN(n765) );
  AND2_X1 U397 ( .A1(n600), .A2(n366), .ZN(n601) );
  NAND2_X1 U398 ( .A1(n371), .A2(n595), .ZN(n596) );
  XNOR2_X1 U399 ( .A(n593), .B(KEYINPUT79), .ZN(n371) );
  INV_X1 U400 ( .A(n594), .ZN(n373) );
  NOR2_X1 U401 ( .A1(n702), .A2(n542), .ZN(n543) );
  AND2_X1 U402 ( .A1(n433), .A2(n359), .ZN(n442) );
  XNOR2_X1 U403 ( .A(n731), .B(n730), .ZN(n732) );
  BUF_X1 U404 ( .A(n744), .Z(n353) );
  XNOR2_X1 U405 ( .A(n570), .B(n569), .ZN(n762) );
  XNOR2_X1 U406 ( .A(n565), .B(KEYINPUT103), .ZN(n571) );
  XNOR2_X1 U407 ( .A(n622), .B(KEYINPUT109), .ZN(n759) );
  NOR2_X1 U408 ( .A1(n618), .A2(n617), .ZN(n619) );
  AND2_X1 U409 ( .A1(n572), .A2(n400), .ZN(n581) );
  XNOR2_X1 U410 ( .A(n543), .B(KEYINPUT66), .ZN(n572) );
  BUF_X1 U411 ( .A(n548), .Z(n638) );
  XNOR2_X1 U412 ( .A(n513), .B(n512), .ZN(n542) );
  NOR2_X1 U413 ( .A1(n745), .A2(G902), .ZN(n513) );
  XNOR2_X1 U414 ( .A(KEYINPUT16), .B(G122), .ZN(n522) );
  XNOR2_X1 U415 ( .A(G137), .B(G140), .ZN(n503) );
  AND2_X2 U416 ( .A1(n420), .A2(n355), .ZN(n744) );
  XNOR2_X2 U417 ( .A(n562), .B(KEYINPUT22), .ZN(n592) );
  XNOR2_X1 U418 ( .A(n750), .B(G146), .ZN(n493) );
  NAND2_X1 U419 ( .A1(n763), .A2(KEYINPUT80), .ZN(n378) );
  XNOR2_X1 U420 ( .A(n408), .B(KEYINPUT88), .ZN(n407) );
  INV_X1 U421 ( .A(KEYINPUT24), .ZN(n408) );
  XNOR2_X1 U422 ( .A(G128), .B(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U423 ( .A(G119), .B(KEYINPUT23), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n580), .B(KEYINPUT101), .ZN(n698) );
  NAND2_X1 U425 ( .A1(n694), .A2(n438), .ZN(n437) );
  INV_X1 U426 ( .A(KEYINPUT30), .ZN(n438) );
  XNOR2_X1 U427 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n453) );
  XNOR2_X1 U428 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n529) );
  INV_X1 U429 ( .A(G128), .ZN(n422) );
  INV_X1 U430 ( .A(G237), .ZN(n517) );
  INV_X1 U431 ( .A(n572), .ZN(n401) );
  NOR2_X1 U432 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U433 ( .A1(n436), .A2(n434), .ZN(n430) );
  NOR2_X1 U434 ( .A1(n442), .A2(n437), .ZN(n429) );
  NAND2_X1 U435 ( .A1(n435), .A2(KEYINPUT30), .ZN(n434) );
  NAND2_X1 U436 ( .A1(n358), .A2(n442), .ZN(n431) );
  OR2_X1 U437 ( .A1(n665), .A2(n440), .ZN(n439) );
  INV_X1 U438 ( .A(KEYINPUT68), .ZN(n487) );
  XOR2_X1 U439 ( .A(KEYINPUT9), .B(G122), .Z(n459) );
  XNOR2_X1 U440 ( .A(G107), .B(G116), .ZN(n458) );
  XNOR2_X1 U441 ( .A(n526), .B(G134), .ZN(n457) );
  NOR2_X1 U442 ( .A1(n690), .A2(n689), .ZN(n691) );
  INV_X1 U443 ( .A(KEYINPUT71), .ZN(n421) );
  XNOR2_X1 U444 ( .A(n465), .B(n464), .ZN(n578) );
  NAND2_X1 U445 ( .A1(n744), .A2(G472), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n451), .B(n447), .ZN(n394) );
  INV_X1 U447 ( .A(n759), .ZN(n423) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n496) );
  INV_X1 U449 ( .A(n694), .ZN(n435) );
  OR2_X1 U450 ( .A1(n437), .A2(n440), .ZN(n432) );
  NAND2_X1 U451 ( .A1(n441), .A2(n518), .ZN(n440) );
  INV_X1 U452 ( .A(n494), .ZN(n441) );
  XOR2_X1 U453 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n481) );
  XNOR2_X1 U454 ( .A(G101), .B(G137), .ZN(n483) );
  AND2_X1 U455 ( .A1(n378), .A2(KEYINPUT44), .ZN(n415) );
  XNOR2_X1 U456 ( .A(n404), .B(n403), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n407), .B(n406), .ZN(n405) );
  XNOR2_X1 U458 ( .A(KEYINPUT90), .B(KEYINPUT69), .ZN(n404) );
  XNOR2_X1 U459 ( .A(G104), .B(G143), .ZN(n466) );
  XOR2_X1 U460 ( .A(G131), .B(G140), .Z(n467) );
  XNOR2_X1 U461 ( .A(G113), .B(G122), .ZN(n468) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n469) );
  NOR2_X1 U463 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U464 ( .A(n457), .B(n444), .ZN(n750) );
  XNOR2_X1 U465 ( .A(KEYINPUT4), .B(G131), .ZN(n444) );
  XNOR2_X1 U466 ( .A(n645), .B(n644), .ZN(n697) );
  INV_X1 U467 ( .A(KEYINPUT107), .ZN(n644) );
  XNOR2_X1 U468 ( .A(n638), .B(n377), .ZN(n643) );
  INV_X1 U469 ( .A(KEYINPUT38), .ZN(n377) );
  NAND2_X1 U470 ( .A1(n574), .A2(n388), .ZN(n384) );
  NAND2_X1 U471 ( .A1(n373), .A2(n357), .ZN(n624) );
  XNOR2_X1 U472 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U473 ( .A(n530), .B(n529), .ZN(n531) );
  NAND2_X1 U474 ( .A1(n534), .A2(G214), .ZN(n694) );
  NOR2_X1 U475 ( .A1(n708), .A2(n401), .ZN(n585) );
  NOR2_X1 U476 ( .A1(n541), .A2(n540), .ZN(n544) );
  XNOR2_X1 U477 ( .A(n579), .B(KEYINPUT100), .ZN(n671) );
  XNOR2_X1 U478 ( .A(n462), .B(n461), .ZN(n740) );
  XNOR2_X1 U479 ( .A(n457), .B(n460), .ZN(n461) );
  NAND2_X1 U480 ( .A1(n729), .A2(n728), .ZN(n731) );
  NOR2_X1 U481 ( .A1(n692), .A2(n586), .ZN(n389) );
  INV_X1 U482 ( .A(KEYINPUT75), .ZN(n374) );
  INV_X1 U483 ( .A(n671), .ZN(n682) );
  NAND2_X1 U484 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U485 ( .A(n393), .B(n361), .ZN(n392) );
  INV_X1 U486 ( .A(KEYINPUT124), .ZN(n409) );
  NAND2_X1 U487 ( .A1(n411), .A2(n391), .ZN(n410) );
  XNOR2_X1 U488 ( .A(n412), .B(n363), .ZN(n411) );
  INV_X1 U489 ( .A(KEYINPUT60), .ZN(n416) );
  NAND2_X1 U490 ( .A1(n418), .A2(n391), .ZN(n417) );
  XNOR2_X1 U491 ( .A(n419), .B(n362), .ZN(n418) );
  XNOR2_X1 U492 ( .A(n735), .B(n376), .ZN(n737) );
  XNOR2_X1 U493 ( .A(n736), .B(n734), .ZN(n376) );
  INV_X1 U494 ( .A(KEYINPUT56), .ZN(n368) );
  AND2_X1 U495 ( .A1(n578), .A2(n558), .ZN(n354) );
  AND2_X1 U496 ( .A1(n660), .A2(n659), .ZN(n355) );
  XNOR2_X1 U497 ( .A(n452), .B(G469), .ZN(n623) );
  INV_X1 U498 ( .A(n623), .ZN(n400) );
  NOR2_X1 U499 ( .A1(n556), .A2(n555), .ZN(n356) );
  NOR2_X1 U500 ( .A1(n702), .A2(n541), .ZN(n357) );
  AND2_X1 U501 ( .A1(n439), .A2(KEYINPUT30), .ZN(n358) );
  NAND2_X1 U502 ( .A1(n494), .A2(G902), .ZN(n359) );
  XOR2_X1 U503 ( .A(n557), .B(KEYINPUT0), .Z(n360) );
  XOR2_X1 U504 ( .A(n666), .B(KEYINPUT62), .Z(n361) );
  XOR2_X1 U505 ( .A(n739), .B(n738), .Z(n362) );
  XNOR2_X1 U506 ( .A(n394), .B(n493), .ZN(n736) );
  XOR2_X1 U507 ( .A(n745), .B(n746), .Z(n363) );
  XOR2_X1 U508 ( .A(n663), .B(n662), .Z(n364) );
  NAND2_X1 U509 ( .A1(n598), .A2(KEYINPUT80), .ZN(n365) );
  AND2_X1 U510 ( .A1(n599), .A2(KEYINPUT80), .ZN(n366) );
  NOR2_X1 U511 ( .A1(n752), .A2(G952), .ZN(n747) );
  INV_X1 U512 ( .A(n747), .ZN(n391) );
  XOR2_X1 U513 ( .A(KEYINPUT63), .B(KEYINPUT111), .Z(n367) );
  XNOR2_X1 U514 ( .A(n369), .B(n368), .ZN(G51) );
  NAND2_X1 U515 ( .A1(n370), .A2(n391), .ZN(n369) );
  XNOR2_X1 U516 ( .A(n664), .B(n364), .ZN(n370) );
  XNOR2_X2 U517 ( .A(n372), .B(KEYINPUT45), .ZN(n686) );
  NAND2_X1 U518 ( .A1(n379), .A2(n604), .ZN(n372) );
  XNOR2_X1 U519 ( .A(n405), .B(n402), .ZN(n507) );
  INV_X1 U520 ( .A(n503), .ZN(n502) );
  XNOR2_X1 U521 ( .A(n375), .B(n374), .ZN(n678) );
  NAND2_X1 U522 ( .A1(n630), .A2(KEYINPUT47), .ZN(n427) );
  NAND2_X1 U523 ( .A1(n693), .A2(n694), .ZN(n645) );
  XNOR2_X2 U524 ( .A(n576), .B(KEYINPUT35), .ZN(n763) );
  NAND2_X1 U525 ( .A1(n414), .A2(n365), .ZN(n381) );
  NAND2_X1 U526 ( .A1(n383), .A2(n382), .ZN(n692) );
  NAND2_X1 U527 ( .A1(n387), .A2(n386), .ZN(n382) );
  AND2_X1 U528 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n708), .A2(n388), .ZN(n385) );
  INV_X1 U530 ( .A(n574), .ZN(n386) );
  NOR2_X1 U531 ( .A1(n708), .A2(n388), .ZN(n387) );
  INV_X1 U532 ( .A(KEYINPUT33), .ZN(n388) );
  XNOR2_X1 U533 ( .A(n389), .B(KEYINPUT34), .ZN(n575) );
  XNOR2_X1 U534 ( .A(n390), .B(n367), .ZN(G57) );
  AND2_X2 U535 ( .A1(n395), .A2(n443), .ZN(n687) );
  XNOR2_X1 U536 ( .A(n397), .B(n396), .ZN(n395) );
  INV_X1 U537 ( .A(KEYINPUT48), .ZN(n396) );
  NAND2_X1 U538 ( .A1(n399), .A2(n398), .ZN(n397) );
  XNOR2_X1 U539 ( .A(n650), .B(KEYINPUT46), .ZN(n398) );
  AND2_X2 U540 ( .A1(n637), .A2(n636), .ZN(n399) );
  NAND2_X1 U541 ( .A1(n708), .A2(n401), .ZN(n709) );
  XNOR2_X1 U542 ( .A(n410), .B(n409), .ZN(G66) );
  NAND2_X1 U543 ( .A1(n744), .A2(G217), .ZN(n412) );
  NOR2_X2 U544 ( .A1(n629), .A2(n356), .ZN(n413) );
  XNOR2_X2 U545 ( .A(n616), .B(n552), .ZN(n629) );
  XNOR2_X2 U546 ( .A(n413), .B(n360), .ZN(n586) );
  NAND2_X1 U547 ( .A1(n415), .A2(n600), .ZN(n414) );
  XNOR2_X1 U548 ( .A(n417), .B(n416), .ZN(G60) );
  NAND2_X1 U549 ( .A1(n744), .A2(G475), .ZN(n419) );
  XNOR2_X2 U550 ( .A(n551), .B(n550), .ZN(n616) );
  XNOR2_X2 U551 ( .A(n538), .B(n537), .ZN(n548) );
  XNOR2_X2 U552 ( .A(n450), .B(n449), .ZN(n523) );
  NAND2_X1 U553 ( .A1(n691), .A2(n420), .ZN(n729) );
  XNOR2_X2 U554 ( .A(n655), .B(n421), .ZN(n420) );
  XNOR2_X1 U555 ( .A(n425), .B(KEYINPUT77), .ZN(n424) );
  NAND2_X1 U556 ( .A1(n427), .A2(n426), .ZN(n425) );
  XNOR2_X1 U557 ( .A(n634), .B(n633), .ZN(n426) );
  NAND2_X1 U558 ( .A1(n431), .A2(n428), .ZN(n540) );
  OR2_X1 U559 ( .A1(n665), .A2(n432), .ZN(n436) );
  NAND2_X1 U560 ( .A1(n665), .A2(n494), .ZN(n433) );
  OR2_X1 U561 ( .A1(n639), .A2(n547), .ZN(n631) );
  XOR2_X2 U562 ( .A(G125), .B(G146), .Z(n527) );
  AND2_X1 U563 ( .A1(n653), .A2(n652), .ZN(n443) );
  INV_X1 U564 ( .A(KEYINPUT76), .ZN(n633) );
  XNOR2_X1 U565 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U566 ( .A(n485), .B(n484), .ZN(n491) );
  XNOR2_X1 U567 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U568 ( .A(n463), .B(G478), .ZN(n464) );
  INV_X1 U569 ( .A(KEYINPUT121), .ZN(n730) );
  XNOR2_X1 U570 ( .A(n649), .B(n648), .ZN(n764) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n521) );
  NAND2_X1 U572 ( .A1(G227), .A2(n752), .ZN(n446) );
  INV_X1 U573 ( .A(KEYINPUT73), .ZN(n445) );
  XOR2_X1 U574 ( .A(KEYINPUT87), .B(n502), .Z(n749) );
  XNOR2_X1 U575 ( .A(n523), .B(n749), .ZN(n451) );
  NOR2_X1 U576 ( .A1(G902), .A2(n736), .ZN(n452) );
  INV_X1 U577 ( .A(n708), .ZN(n620) );
  XOR2_X1 U578 ( .A(KEYINPUT7), .B(KEYINPUT97), .Z(n456) );
  NAND2_X1 U579 ( .A1(n752), .A2(G234), .ZN(n454) );
  XNOR2_X1 U580 ( .A(n454), .B(n453), .ZN(n505) );
  NAND2_X1 U581 ( .A1(G217), .A2(n505), .ZN(n455) );
  XNOR2_X1 U582 ( .A(n456), .B(n455), .ZN(n462) );
  XNOR2_X1 U583 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U584 ( .A1(G902), .A2(n740), .ZN(n465) );
  XNOR2_X1 U585 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U586 ( .A(n467), .B(n466), .ZN(n471) );
  XNOR2_X1 U587 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U588 ( .A(n471), .B(n470), .Z(n473) );
  NAND2_X1 U589 ( .A1(n479), .A2(G214), .ZN(n472) );
  XNOR2_X1 U590 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n748), .B(n474), .ZN(n739) );
  NOR2_X1 U592 ( .A1(G902), .A2(n739), .ZN(n478) );
  XOR2_X1 U593 ( .A(KEYINPUT13), .B(KEYINPUT96), .Z(n476) );
  XNOR2_X1 U594 ( .A(KEYINPUT95), .B(G475), .ZN(n475) );
  XOR2_X1 U595 ( .A(n476), .B(n475), .Z(n477) );
  XNOR2_X1 U596 ( .A(n478), .B(n477), .ZN(n577) );
  NOR2_X1 U597 ( .A1(n578), .A2(n577), .ZN(n680) );
  NAND2_X1 U598 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U599 ( .A(n481), .B(n480), .ZN(n485) );
  INV_X1 U600 ( .A(KEYINPUT93), .ZN(n482) );
  XNOR2_X1 U601 ( .A(G119), .B(G116), .ZN(n486) );
  XNOR2_X1 U602 ( .A(n486), .B(KEYINPUT3), .ZN(n489) );
  XNOR2_X1 U603 ( .A(n487), .B(G113), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n489), .B(n488), .ZN(n524) );
  INV_X1 U605 ( .A(n524), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U607 ( .A(KEYINPUT70), .B(G472), .ZN(n494) );
  INV_X1 U608 ( .A(KEYINPUT6), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n706), .B(n495), .ZN(n573) );
  INV_X1 U610 ( .A(n573), .ZN(n591) );
  XNOR2_X1 U611 ( .A(n496), .B(KEYINPUT14), .ZN(n498) );
  NAND2_X1 U612 ( .A1(G952), .A2(n498), .ZN(n497) );
  XNOR2_X1 U613 ( .A(n497), .B(KEYINPUT84), .ZN(n724) );
  NOR2_X1 U614 ( .A1(n724), .A2(G953), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G902), .A2(n498), .ZN(n553) );
  NOR2_X1 U616 ( .A1(G900), .A2(n553), .ZN(n499) );
  NAND2_X1 U617 ( .A1(G953), .A2(n499), .ZN(n500) );
  XOR2_X1 U618 ( .A(KEYINPUT104), .B(n500), .Z(n501) );
  NOR2_X1 U619 ( .A1(n556), .A2(n501), .ZN(n541) );
  XOR2_X1 U620 ( .A(G110), .B(n503), .Z(n504) );
  XNOR2_X1 U621 ( .A(n748), .B(n504), .ZN(n509) );
  NAND2_X1 U622 ( .A1(G221), .A2(n505), .ZN(n506) );
  XNOR2_X1 U623 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U624 ( .A(n509), .B(n508), .ZN(n745) );
  XNOR2_X1 U625 ( .A(G902), .B(KEYINPUT15), .ZN(n658) );
  NAND2_X1 U626 ( .A1(G234), .A2(n658), .ZN(n510) );
  XNOR2_X1 U627 ( .A(KEYINPUT20), .B(n510), .ZN(n514) );
  AND2_X1 U628 ( .A1(n514), .A2(G217), .ZN(n511) );
  XNOR2_X1 U629 ( .A(KEYINPUT25), .B(n511), .ZN(n512) );
  INV_X1 U630 ( .A(n542), .ZN(n594) );
  AND2_X1 U631 ( .A1(n514), .A2(G221), .ZN(n515) );
  XNOR2_X1 U632 ( .A(n515), .B(KEYINPUT21), .ZN(n559) );
  NOR2_X1 U633 ( .A1(n591), .A2(n624), .ZN(n516) );
  NAND2_X1 U634 ( .A1(n680), .A2(n516), .ZN(n618) );
  NOR2_X1 U635 ( .A1(n620), .A2(n618), .ZN(n519) );
  INV_X1 U636 ( .A(G902), .ZN(n518) );
  NAND2_X1 U637 ( .A1(n518), .A2(n517), .ZN(n534) );
  NAND2_X1 U638 ( .A1(n519), .A2(n694), .ZN(n520) );
  XNOR2_X1 U639 ( .A(n521), .B(n520), .ZN(n539) );
  XOR2_X1 U640 ( .A(n526), .B(n527), .Z(n532) );
  NAND2_X1 U641 ( .A1(n752), .A2(G224), .ZN(n528) );
  XNOR2_X1 U642 ( .A(n528), .B(KEYINPUT17), .ZN(n530) );
  XNOR2_X1 U643 ( .A(n611), .B(n533), .ZN(n661) );
  NAND2_X1 U644 ( .A1(n661), .A2(n658), .ZN(n538) );
  NAND2_X1 U645 ( .A1(n534), .A2(G210), .ZN(n536) );
  INV_X1 U646 ( .A(KEYINPUT83), .ZN(n535) );
  XNOR2_X1 U647 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U648 ( .A1(n539), .A2(n638), .ZN(n652) );
  XNOR2_X1 U649 ( .A(n652), .B(G140), .ZN(G42) );
  INV_X1 U650 ( .A(n559), .ZN(n702) );
  NAND2_X1 U651 ( .A1(n544), .A2(n581), .ZN(n545) );
  XNOR2_X1 U652 ( .A(KEYINPUT72), .B(n545), .ZN(n639) );
  INV_X1 U653 ( .A(n638), .ZN(n546) );
  INV_X1 U654 ( .A(n577), .ZN(n558) );
  NAND2_X1 U655 ( .A1(n546), .A2(n354), .ZN(n547) );
  XNOR2_X1 U656 ( .A(n631), .B(G143), .ZN(G45) );
  INV_X1 U657 ( .A(n548), .ZN(n549) );
  NAND2_X1 U658 ( .A1(n549), .A2(n694), .ZN(n551) );
  INV_X1 U659 ( .A(KEYINPUT82), .ZN(n550) );
  XNOR2_X1 U660 ( .A(KEYINPUT64), .B(KEYINPUT19), .ZN(n552) );
  XNOR2_X1 U661 ( .A(G898), .B(KEYINPUT85), .ZN(n608) );
  NAND2_X1 U662 ( .A1(G953), .A2(n608), .ZN(n612) );
  NOR2_X1 U663 ( .A1(n553), .A2(n612), .ZN(n554) );
  XNOR2_X1 U664 ( .A(n554), .B(KEYINPUT86), .ZN(n555) );
  INV_X1 U665 ( .A(KEYINPUT65), .ZN(n557) );
  OR2_X1 U666 ( .A1(n578), .A2(n558), .ZN(n696) );
  INV_X1 U667 ( .A(n696), .ZN(n560) );
  NAND2_X1 U668 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X2 U669 ( .A1(n586), .A2(n561), .ZN(n562) );
  NOR2_X1 U670 ( .A1(n706), .A2(n594), .ZN(n563) );
  AND2_X1 U671 ( .A1(n708), .A2(n563), .ZN(n564) );
  NAND2_X1 U672 ( .A1(n592), .A2(n564), .ZN(n565) );
  XOR2_X1 U673 ( .A(n571), .B(G110), .Z(G12) );
  NAND2_X1 U674 ( .A1(n591), .A2(n373), .ZN(n566) );
  NOR2_X1 U675 ( .A1(n708), .A2(n566), .ZN(n567) );
  XNOR2_X1 U676 ( .A(KEYINPUT74), .B(n567), .ZN(n568) );
  NAND2_X1 U677 ( .A1(n592), .A2(n568), .ZN(n570) );
  INV_X1 U678 ( .A(KEYINPUT32), .ZN(n569) );
  NAND2_X1 U679 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U680 ( .A1(n575), .A2(n354), .ZN(n576) );
  INV_X1 U681 ( .A(KEYINPUT44), .ZN(n598) );
  INV_X1 U682 ( .A(n680), .ZN(n641) );
  NAND2_X1 U683 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U684 ( .A1(n641), .A2(n671), .ZN(n580) );
  INV_X1 U685 ( .A(n581), .ZN(n582) );
  NOR2_X1 U686 ( .A1(n586), .A2(n582), .ZN(n583) );
  XNOR2_X1 U687 ( .A(n583), .B(KEYINPUT91), .ZN(n584) );
  NOR2_X1 U688 ( .A1(n706), .A2(n584), .ZN(n672) );
  XNOR2_X1 U689 ( .A(KEYINPUT31), .B(KEYINPUT94), .ZN(n588) );
  NAND2_X1 U690 ( .A1(n706), .A2(n585), .ZN(n713) );
  NOR2_X1 U691 ( .A1(n713), .A2(n586), .ZN(n587) );
  XOR2_X1 U692 ( .A(n588), .B(n587), .Z(n683) );
  NOR2_X1 U693 ( .A1(n672), .A2(n683), .ZN(n589) );
  OR2_X1 U694 ( .A1(n698), .A2(n589), .ZN(n590) );
  NAND2_X1 U695 ( .A1(n592), .A2(n591), .ZN(n593) );
  AND2_X1 U696 ( .A1(n708), .A2(n594), .ZN(n595) );
  OR2_X1 U697 ( .A1(n600), .A2(KEYINPUT81), .ZN(n603) );
  INV_X1 U698 ( .A(KEYINPUT81), .ZN(n597) );
  NAND2_X1 U699 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U700 ( .A1(n601), .A2(n763), .ZN(n602) );
  NAND2_X1 U701 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U702 ( .A1(n686), .A2(n752), .ZN(n605) );
  XNOR2_X1 U703 ( .A(n605), .B(KEYINPUT125), .ZN(n610) );
  NAND2_X1 U704 ( .A1(G953), .A2(G224), .ZN(n606) );
  XOR2_X1 U705 ( .A(KEYINPUT61), .B(n606), .Z(n607) );
  NOR2_X1 U706 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U707 ( .A1(n610), .A2(n609), .ZN(n615) );
  INV_X1 U708 ( .A(n611), .ZN(n613) );
  NAND2_X1 U709 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U710 ( .A(n615), .B(n614), .ZN(G69) );
  INV_X1 U711 ( .A(n616), .ZN(n617) );
  XNOR2_X1 U712 ( .A(n619), .B(KEYINPUT36), .ZN(n621) );
  NAND2_X1 U713 ( .A1(n621), .A2(n620), .ZN(n622) );
  INV_X1 U714 ( .A(n706), .ZN(n625) );
  XNOR2_X1 U715 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n626) );
  XNOR2_X1 U716 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U717 ( .A1(n400), .A2(n628), .ZN(n647) );
  INV_X1 U718 ( .A(n678), .ZN(n630) );
  NAND2_X1 U719 ( .A1(KEYINPUT47), .A2(n698), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n634) );
  NOR2_X1 U721 ( .A1(KEYINPUT47), .A2(n698), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n678), .A2(n635), .ZN(n636) );
  NOR2_X1 U723 ( .A1(n639), .A2(n643), .ZN(n640) );
  XNOR2_X1 U724 ( .A(n640), .B(KEYINPUT39), .ZN(n651) );
  NOR2_X1 U725 ( .A1(n641), .A2(n651), .ZN(n642) );
  XNOR2_X1 U726 ( .A(n642), .B(KEYINPUT40), .ZN(n766) );
  XOR2_X1 U727 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n649) );
  INV_X1 U728 ( .A(n643), .ZN(n693) );
  NOR2_X1 U729 ( .A1(n697), .A2(n696), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n646), .B(KEYINPUT41), .ZN(n717) );
  NOR2_X1 U731 ( .A1(n671), .A2(n651), .ZN(n685) );
  INV_X1 U732 ( .A(n685), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n686), .A2(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n686), .A2(n687), .ZN(n657) );
  INV_X1 U735 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n660) );
  INV_X1 U737 ( .A(n658), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n744), .A2(G210), .ZN(n664) );
  BUF_X1 U739 ( .A(n661), .Z(n663) );
  XNOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT110), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n672), .A2(n680), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(G104), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n669) );
  XNOR2_X1 U745 ( .A(G107), .B(KEYINPUT112), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U747 ( .A(KEYINPUT26), .B(n670), .Z(n674) );
  NAND2_X1 U748 ( .A1(n672), .A2(n682), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n674), .B(n673), .ZN(G9) );
  XOR2_X1 U750 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n676) );
  NAND2_X1 U751 ( .A1(n678), .A2(n682), .ZN(n675) );
  XNOR2_X1 U752 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U753 ( .A(G128), .B(n677), .ZN(G30) );
  NAND2_X1 U754 ( .A1(n678), .A2(n680), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(G146), .ZN(G48) );
  NAND2_X1 U756 ( .A1(n683), .A2(n680), .ZN(n681) );
  XNOR2_X1 U757 ( .A(n681), .B(G113), .ZN(G15) );
  NAND2_X1 U758 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n684), .B(G116), .ZN(G18) );
  XOR2_X1 U760 ( .A(G134), .B(n685), .Z(G36) );
  NOR2_X1 U761 ( .A1(n686), .A2(KEYINPUT2), .ZN(n690) );
  NOR2_X1 U762 ( .A1(n687), .A2(KEYINPUT2), .ZN(n688) );
  XNOR2_X1 U763 ( .A(n688), .B(KEYINPUT78), .ZN(n689) );
  NOR2_X1 U764 ( .A1(n693), .A2(n694), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n692), .A2(n701), .ZN(n720) );
  XNOR2_X1 U769 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n716) );
  XNOR2_X1 U770 ( .A(KEYINPUT49), .B(KEYINPUT115), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n373), .A2(n702), .ZN(n703) );
  XOR2_X1 U772 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n707), .B(KEYINPUT116), .ZN(n712) );
  XOR2_X1 U775 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n710) );
  XNOR2_X1 U776 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U779 ( .A(n716), .B(n715), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U782 ( .A(n721), .B(KEYINPUT52), .Z(n722) );
  XNOR2_X1 U783 ( .A(KEYINPUT119), .B(n722), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n724), .A2(n723), .ZN(n726) );
  NOR2_X1 U785 ( .A1(n717), .A2(n692), .ZN(n725) );
  NOR2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n727), .B(KEYINPUT120), .ZN(n728) );
  XNOR2_X1 U788 ( .A(KEYINPUT53), .B(n733), .ZN(G75) );
  NAND2_X1 U789 ( .A1(n353), .A2(G469), .ZN(n735) );
  XOR2_X1 U790 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n734) );
  NOR2_X1 U791 ( .A1(n747), .A2(n737), .ZN(G54) );
  INV_X1 U792 ( .A(KEYINPUT59), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n353), .A2(G478), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n740), .B(KEYINPUT122), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U796 ( .A1(n747), .A2(n743), .ZN(G63) );
  INV_X1 U797 ( .A(KEYINPUT123), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n748), .B(n749), .ZN(n751) );
  XOR2_X1 U799 ( .A(n750), .B(n751), .Z(n754) );
  XOR2_X1 U800 ( .A(n754), .B(n687), .Z(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(n752), .ZN(n758) );
  XNOR2_X1 U802 ( .A(G227), .B(n754), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(G953), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n758), .A2(n757), .ZN(G72) );
  XNOR2_X1 U806 ( .A(n759), .B(G125), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n760), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U808 ( .A(G119), .B(KEYINPUT126), .Z(n761) );
  XNOR2_X1 U809 ( .A(n762), .B(n761), .ZN(G21) );
  XOR2_X1 U810 ( .A(n763), .B(G122), .Z(G24) );
  XOR2_X1 U811 ( .A(G137), .B(n764), .Z(G39) );
  XNOR2_X1 U812 ( .A(n765), .B(G101), .ZN(G3) );
  XOR2_X1 U813 ( .A(G131), .B(n766), .Z(G33) );
endmodule

