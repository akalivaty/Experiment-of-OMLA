//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND4_X1   g002(.A1(G143), .A2(new_n187), .A3(new_n188), .A4(G214), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n191));
  OAI211_X1 g005(.A(KEYINPUT18), .B(G131), .C1(new_n189), .C2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT18), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n195), .B(new_n196), .C1(new_n197), .C2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n192), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT87), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT87), .B1(new_n202), .B2(new_n204), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n200), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n205), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n213), .A3(G146), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT17), .B(G131), .C1(new_n189), .C2(new_n191), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n189), .A2(new_n191), .A3(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n198), .B1(new_n195), .B2(new_n196), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n222));
  AOI22_X1  g036(.A1(KEYINPUT89), .A2(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT89), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n215), .A2(new_n217), .A3(new_n224), .A4(new_n216), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n211), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G113), .B(G122), .ZN(new_n227));
  INV_X1    g041(.A(G104), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n218), .A2(KEYINPUT89), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n222), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n225), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n210), .A2(new_n206), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n199), .A3(new_n192), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n229), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT90), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(KEYINPUT90), .A3(new_n235), .A4(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n230), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(G475), .B1(new_n240), .B2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G478), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(KEYINPUT15), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT73), .B(G217), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT9), .B(G234), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n246), .A2(G953), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT13), .B1(new_n250), .B2(G143), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(G128), .B(G143), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n253), .B(new_n254), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT92), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(G122), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n258), .A2(KEYINPUT93), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n262));
  INV_X1    g076(.A(G122), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(KEYINPUT92), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(KEYINPUT92), .ZN(new_n265));
  OAI21_X1  g079(.A(G116), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n266), .B2(new_n259), .ZN(new_n267));
  OAI21_X1  g081(.A(G107), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT93), .B1(new_n258), .B2(new_n260), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n262), .A3(new_n259), .ZN(new_n270));
  INV_X1    g084(.A(G107), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n255), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n259), .B(KEYINPUT14), .ZN(new_n274));
  OAI21_X1  g088(.A(G107), .B1(new_n274), .B2(new_n258), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n254), .B(new_n252), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n249), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n255), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n261), .A2(new_n267), .A3(G107), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n271), .B1(new_n269), .B2(new_n270), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n275), .A3(new_n276), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(new_n248), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n244), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n286), .B(new_n243), .C1(new_n278), .C2(new_n284), .ZN(new_n289));
  INV_X1    g103(.A(G234), .ZN(new_n290));
  OAI211_X1 g104(.A(G952), .B(new_n188), .C1(new_n290), .C2(new_n187), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT94), .Z(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n188), .B(new_n287), .C1(G234), .C2(G237), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT21), .B(G898), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n288), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT19), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n202), .A2(new_n204), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT88), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n209), .B2(KEYINPUT19), .ZN(new_n301));
  NOR4_X1   g115(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT88), .A4(new_n298), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n205), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n221), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n216), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n235), .ZN(new_n306));
  INV_X1    g120(.A(new_n229), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT90), .B1(new_n226), .B2(new_n229), .ZN(new_n309));
  INV_X1    g123(.A(new_n239), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT91), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT20), .ZN(new_n313));
  NOR2_X1   g127(.A1(G475), .A2(G902), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n229), .B1(new_n305), .B2(new_n235), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n238), .B2(new_n239), .ZN(new_n317));
  INV_X1    g131(.A(new_n314), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT20), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n312), .B1(new_n321), .B2(new_n313), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n241), .B(new_n297), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n326));
  XNOR2_X1  g140(.A(G110), .B(G122), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n271), .A2(KEYINPUT79), .A3(G104), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n271), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(G104), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n228), .A2(G107), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n329), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G113), .ZN(new_n340));
  INV_X1    g154(.A(G113), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT2), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT68), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n339), .A2(G113), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  XOR2_X1   g162(.A(G116), .B(G119), .Z(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n344), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n346), .ZN(new_n351));
  XNOR2_X1  g165(.A(G116), .B(G119), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n352), .B1(KEYINPUT68), .B2(new_n351), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n344), .B1(new_n355), .B2(new_n348), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n338), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n335), .A2(new_n329), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n332), .B2(new_n333), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n358), .B1(new_n362), .B2(new_n336), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n334), .A2(new_n335), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G101), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT80), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n357), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n271), .A2(G104), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n329), .B1(new_n370), .B2(new_n335), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(KEYINPUT5), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n257), .A2(KEYINPUT5), .A3(G119), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n341), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n374), .A2(new_n376), .B1(new_n351), .B2(new_n352), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n373), .B1(new_n372), .B2(new_n377), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n326), .B(new_n328), .C1(new_n369), .C2(new_n381), .ZN(new_n382));
  NOR4_X1   g196(.A1(new_n336), .A2(new_n358), .A3(new_n366), .A4(new_n360), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT80), .B1(new_n365), .B2(new_n367), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n327), .B(new_n380), .C1(new_n385), .C2(new_n357), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT6), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n343), .A2(new_n349), .ZN(new_n388));
  INV_X1    g202(.A(new_n348), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT69), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n353), .A3(new_n350), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n391), .B(new_n338), .C1(new_n383), .C2(new_n384), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n327), .B1(new_n392), .B2(new_n380), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n325), .B(new_n382), .C1(new_n387), .C2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n328), .B1(new_n369), .B2(new_n381), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n395), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n386), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G128), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n205), .A2(G143), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n194), .A2(G146), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(KEYINPUT64), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  XNOR2_X1  g218(.A(G143), .B(G146), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n398), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT0), .A3(G128), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n400), .A2(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n402), .A2(new_n410), .A3(G128), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n400), .B(new_n401), .C1(KEYINPUT1), .C2(new_n250), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n203), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n188), .A2(G224), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n397), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  AND2_X1   g234(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n416), .B1(KEYINPUT86), .B2(KEYINPUT7), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n415), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n414), .A4(new_n416), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n327), .B(KEYINPUT8), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n372), .A2(new_n377), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n372), .A2(new_n377), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n429), .B2(new_n386), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n420), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n417), .B1(new_n394), .B2(new_n396), .ZN(new_n433));
  INV_X1    g247(.A(new_n430), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G214), .B1(G237), .B2(G902), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n247), .B2(G902), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT78), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n408), .B1(new_n336), .B2(new_n337), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n383), .B2(new_n384), .ZN(new_n441));
  INV_X1    g255(.A(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(KEYINPUT11), .A3(G134), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n252), .A2(G137), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT11), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n252), .B2(G137), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n198), .A4(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(new_n443), .A3(new_n198), .A4(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT65), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n443), .A3(new_n444), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(new_n443), .A3(KEYINPUT66), .A4(new_n444), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(G131), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n453), .B1(new_n452), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n372), .A2(new_n412), .A3(new_n411), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT10), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n413), .A2(new_n360), .A3(new_n371), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT10), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n441), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(G110), .B(G140), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n188), .A2(G227), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n457), .A2(G131), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n473), .A2(new_n456), .B1(new_n449), .B2(new_n451), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n441), .B2(new_n467), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n452), .A2(new_n458), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n413), .B1(new_n360), .B2(new_n371), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n479), .B2(new_n464), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n462), .A2(new_n478), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n441), .A2(new_n461), .A3(new_n467), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n472), .A2(new_n476), .B1(new_n487), .B2(new_n471), .ZN(new_n488));
  OAI21_X1  g302(.A(G469), .B1(new_n488), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT83), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n477), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n483), .B2(new_n477), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n482), .A2(KEYINPUT83), .A3(new_n484), .ZN(new_n494));
  INV_X1    g308(.A(new_n471), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n486), .A4(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n471), .B1(new_n468), .B2(new_n475), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n287), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n439), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n324), .A2(new_n436), .A3(new_n437), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n408), .B1(new_n452), .B2(new_n458), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n252), .A2(G137), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n442), .A2(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n411), .A2(new_n506), .A3(new_n412), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n449), .B2(new_n451), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n391), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n354), .A2(new_n356), .ZN(new_n510));
  INV_X1    g324(.A(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n452), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n512), .C1(new_n408), .C2(new_n474), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n509), .A2(new_n513), .A3(KEYINPUT71), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n515), .B(new_n391), .C1(new_n503), .C2(new_n508), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(KEYINPUT28), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n190), .A2(G210), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT26), .B(G101), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n517), .A2(KEYINPUT29), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n511), .A2(new_n452), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n474), .B2(new_n408), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n508), .A2(new_n526), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n408), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n477), .A2(new_n531), .B1(new_n452), .B2(new_n511), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n510), .B1(new_n532), .B2(KEYINPUT30), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n521), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n513), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n391), .B1(new_n528), .B2(new_n529), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n532), .A2(KEYINPUT28), .A3(new_n510), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n523), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n521), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n524), .B(new_n287), .C1(new_n541), .C2(KEYINPUT29), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n535), .B1(new_n532), .B2(new_n510), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT31), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n526), .A2(new_n508), .B1(new_n477), .B2(new_n531), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n512), .A2(KEYINPUT67), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT30), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT30), .B(new_n512), .C1(new_n474), .C2(new_n408), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n391), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n546), .B(new_n547), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n513), .A2(new_n521), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n530), .B2(new_n533), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT70), .A3(new_n547), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n546), .B1(new_n550), .B2(new_n552), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n560), .A2(KEYINPUT31), .B1(new_n539), .B2(new_n535), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT32), .B(new_n545), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n553), .A2(new_n554), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT70), .B1(new_n557), .B2(new_n547), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n563), .B1(new_n566), .B2(new_n544), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n543), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT23), .B1(new_n250), .B2(G119), .ZN(new_n569));
  INV_X1    g383(.A(G119), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT75), .B1(new_n570), .B2(G128), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n569), .B(new_n571), .Z(new_n572));
  XNOR2_X1  g386(.A(G119), .B(G128), .ZN(new_n573));
  XOR2_X1   g387(.A(KEYINPUT24), .B(G110), .Z(new_n574));
  OAI22_X1  g388(.A1(new_n572), .A2(G110), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n216), .A3(new_n206), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n572), .A2(G110), .B1(new_n573), .B2(new_n574), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n215), .A2(new_n216), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n579), .A3(new_n584), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n286), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n245), .B1(new_n286), .B2(new_n290), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT74), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT77), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n586), .A2(new_n587), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n590), .A2(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n568), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n502), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n329), .ZN(G3));
  INV_X1    g416(.A(new_n437), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n431), .B2(new_n435), .ZN(new_n604));
  INV_X1    g418(.A(new_n296), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n285), .B(KEYINPUT33), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n286), .A2(new_n242), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n285), .A2(new_n287), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n606), .A2(new_n607), .B1(new_n242), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT91), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n319), .A3(new_n315), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n612), .B2(new_n241), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n604), .A2(new_n605), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n439), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n476), .A2(new_n486), .A3(new_n495), .ZN(new_n616));
  INV_X1    g430(.A(new_n487), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n495), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n499), .B1(new_n618), .B2(new_n594), .ZN(new_n619));
  AOI211_X1 g433(.A(G469), .B(new_n286), .C1(new_n496), .C2(new_n497), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n599), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n566), .B2(new_n287), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n545), .B1(new_n559), .B2(new_n561), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n614), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n610), .A2(new_n319), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n243), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n285), .A2(new_n287), .A3(new_n244), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n631), .A2(new_n241), .A3(new_n634), .A4(new_n605), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT95), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n634), .A2(new_n241), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT95), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n605), .A4(new_n631), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n604), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(KEYINPUT96), .A3(new_n604), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n627), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n271), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n590), .A2(new_n593), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n580), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n597), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n626), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n502), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT37), .B(G110), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  NAND2_X1  g472(.A1(new_n566), .A2(new_n544), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT32), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n625), .A2(new_n563), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n653), .B1(new_n662), .B2(new_n543), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n420), .B1(new_n419), .B2(new_n430), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n433), .A2(new_n432), .A3(new_n434), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n437), .B(new_n501), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n293), .B1(new_n668), .B2(new_n294), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n637), .A2(new_n631), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n663), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n436), .B(KEYINPUT38), .Z(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n514), .A2(new_n516), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n594), .B1(new_n676), .B2(new_n521), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n535), .B1(new_n534), .B2(new_n513), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n662), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n288), .A2(new_n289), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n612), .B2(new_n241), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n669), .B(KEYINPUT39), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n501), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n603), .B(new_n654), .C1(new_n686), .C2(KEYINPUT40), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n687), .B1(KEYINPUT40), .B2(new_n686), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n194), .ZN(G45));
  AOI211_X1 g504(.A(new_n669), .B(new_n609), .C1(new_n612), .C2(new_n241), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n663), .A2(new_n667), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT99), .B(G146), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G48));
  INV_X1    g508(.A(KEYINPUT100), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n499), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n498), .B2(new_n287), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n286), .B(new_n696), .C1(new_n496), .C2(new_n497), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n698), .A2(new_n699), .A3(new_n439), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n568), .A2(new_n599), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n614), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT41), .B(G113), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT101), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n702), .B(new_n704), .ZN(G15));
  INV_X1    g519(.A(new_n701), .ZN(new_n706));
  INV_X1    g520(.A(new_n644), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT96), .B1(new_n640), .B2(new_n604), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  NAND3_X1  g524(.A1(new_n604), .A2(new_n324), .A3(new_n700), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n568), .A2(new_n654), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n570), .ZN(G21));
  NOR2_X1   g528(.A1(new_n557), .A2(new_n547), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n555), .B2(new_n558), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n517), .A2(new_n523), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n535), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n545), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n599), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n624), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n698), .A2(new_n699), .A3(new_n439), .A4(new_n296), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n604), .A3(new_n683), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NAND3_X1  g538(.A1(new_n436), .A2(new_n437), .A3(new_n700), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n624), .A2(new_n719), .A3(new_n653), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n691), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND4_X1  g543(.A1(new_n501), .A2(new_n431), .A3(new_n435), .A4(new_n437), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n568), .A3(new_n691), .A4(new_n599), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n660), .A2(new_n661), .B1(G472), .B2(new_n542), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n720), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n691), .A4(new_n731), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  NOR3_X1   g553(.A1(new_n735), .A2(new_n730), .A3(new_n720), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n671), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n618), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT102), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n499), .B1(new_n618), .B2(new_n743), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n620), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n750), .B2(new_n749), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n615), .A3(new_n685), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n609), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n612), .A3(new_n241), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(new_n654), .C1(new_n625), .C2(new_n624), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n431), .A2(new_n435), .A3(new_n437), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT103), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n754), .A2(new_n760), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  NOR3_X1   g579(.A1(new_n568), .A2(new_n762), .A3(new_n599), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n752), .A2(new_n615), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(new_n752), .B2(new_n615), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n691), .B(new_n766), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  NOR2_X1   g586(.A1(new_n698), .A2(new_n699), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT49), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n599), .A2(new_n437), .A3(new_n615), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n774), .B2(KEYINPUT49), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n681), .A2(new_n756), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n674), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n757), .A2(new_n293), .ZN(new_n780));
  INV_X1    g594(.A(new_n700), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n762), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n736), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  INV_X1    g602(.A(G952), .ZN(new_n789));
  INV_X1    g603(.A(new_n782), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n790), .A2(new_n681), .A3(new_n720), .A4(new_n292), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n789), .B(G953), .C1(new_n791), .C2(new_n613), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n780), .A2(new_n721), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n788), .B(new_n792), .C1(new_n725), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n769), .A2(new_n770), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n615), .B2(new_n774), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n780), .A2(new_n721), .A3(new_n763), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n612), .A2(new_n241), .A3(new_n609), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n784), .A2(new_n727), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n793), .A2(new_n437), .A3(new_n675), .A4(new_n781), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT50), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n798), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n787), .B(new_n794), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n796), .A2(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n797), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n801), .B(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n803), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n612), .A2(new_n241), .A3(new_n634), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT106), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n604), .A2(new_n622), .A3(new_n626), .A4(new_n605), .ZN(new_n817));
  OAI22_X1  g631(.A1(new_n816), .A2(new_n817), .B1(new_n701), .B2(new_n614), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n723), .B1(new_n712), .B2(new_n711), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n502), .B1(new_n600), .B2(new_n655), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n643), .A2(new_n644), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n604), .A2(KEYINPUT105), .A3(new_n605), .A4(new_n613), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT105), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n627), .B1(new_n614), .B2(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n822), .A2(new_n706), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n691), .A2(new_n727), .ZN(new_n827));
  INV_X1    g641(.A(new_n631), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n241), .A2(new_n682), .A3(new_n670), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT107), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n634), .A2(new_n669), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n241), .A4(new_n631), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n827), .B1(new_n712), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n835), .A2(new_n731), .B1(new_n740), .B2(new_n671), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n821), .A2(new_n826), .A3(new_n738), .A4(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n663), .B(new_n667), .C1(new_n671), .C2(new_n691), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n653), .A2(new_n670), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n667), .A2(new_n681), .A3(new_n683), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n728), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n728), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n813), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT108), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(KEYINPUT109), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n738), .A2(new_n836), .ZN(new_n851));
  INV_X1    g665(.A(new_n711), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n604), .A2(new_n683), .ZN(new_n853));
  INV_X1    g667(.A(new_n698), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n498), .A2(new_n287), .A3(new_n697), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n615), .A3(new_n605), .A4(new_n855), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n856), .A2(new_n624), .A3(new_n719), .A4(new_n720), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n852), .A2(new_n663), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n702), .ZN(new_n859));
  INV_X1    g673(.A(new_n502), .ZN(new_n860));
  INV_X1    g674(.A(new_n655), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n736), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n817), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n814), .B(KEYINPUT106), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n858), .A2(new_n859), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n825), .A2(new_n823), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n709), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n851), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT109), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n843), .A2(new_n870), .A3(new_n845), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n850), .A2(new_n869), .A3(KEYINPUT53), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(KEYINPUT108), .B(new_n813), .C1(new_n837), .C2(new_n846), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n849), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n837), .A2(new_n846), .A3(new_n813), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n850), .A2(new_n869), .A3(new_n871), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n876), .B(new_n878), .C1(new_n879), .C2(KEYINPUT53), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT110), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT110), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n875), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n812), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n789), .A2(new_n188), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT115), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n779), .B1(new_n885), .B2(new_n887), .ZN(G75));
  NOR2_X1   g702(.A1(new_n879), .A2(KEYINPUT53), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n877), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n287), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n891), .B2(new_n432), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n397), .A2(new_n418), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n433), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n892), .B(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n188), .A2(G952), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT116), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n896), .A2(new_n899), .ZN(G51));
  INV_X1    g714(.A(new_n897), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT54), .B1(new_n889), .B2(new_n877), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n880), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n748), .B(KEYINPUT57), .Z(new_n904));
  AOI22_X1  g718(.A1(new_n903), .A2(new_n904), .B1(new_n497), .B2(new_n496), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n890), .A2(new_n287), .A3(new_n747), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT117), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n909), .B(new_n901), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(G54));
  NAND3_X1  g725(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n317), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n317), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n897), .ZN(G60));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n882), .A2(new_n884), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n606), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n919), .A2(KEYINPUT118), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT118), .B1(new_n919), .B2(new_n920), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n903), .A2(new_n606), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n898), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n651), .B(KEYINPUT119), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n890), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n587), .B(new_n586), .C1(new_n890), .C2(new_n927), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n898), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n931), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  INV_X1    g751(.A(G224), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n295), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT121), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n866), .A2(new_n868), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(G953), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n394), .B(new_n396), .C1(G898), .C2(new_n188), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  AND2_X1   g758(.A1(new_n838), .A2(new_n728), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n689), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n740), .B(new_n685), .C1(new_n613), .C2(new_n864), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n764), .A3(new_n771), .A4(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n951), .B2(KEYINPUT62), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n949), .A2(KEYINPUT123), .A3(new_n958), .A4(new_n950), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(G953), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n530), .A2(new_n551), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n301), .A2(new_n302), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n962), .B(new_n963), .Z(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT124), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n967), .B(new_n964), .C1(new_n968), .C2(G953), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n736), .A2(new_n853), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n741), .B1(new_n753), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n771), .A2(new_n973), .A3(new_n764), .A4(new_n738), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n947), .A2(new_n948), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n970), .B1(new_n976), .B2(G953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n966), .A2(new_n969), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n966), .A2(new_n969), .A3(new_n981), .A4(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT125), .Z(new_n986));
  INV_X1    g800(.A(new_n941), .ZN(new_n987));
  OAI211_X1 g801(.A(KEYINPUT126), .B(new_n986), .C1(new_n976), .C2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n974), .A2(new_n975), .A3(new_n987), .ZN(new_n990));
  INV_X1    g804(.A(new_n986), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n536), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n988), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n968), .B2(new_n941), .ZN(new_n995));
  INV_X1    g809(.A(new_n678), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n994), .B(new_n901), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n874), .A2(new_n536), .A3(new_n996), .A4(new_n985), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(G57));
endmodule


