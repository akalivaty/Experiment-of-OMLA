//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n458), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AOI211_X1 g042(.A(KEYINPUT64), .B(new_n467), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n467), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT66), .B1(new_n467), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G101), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n459), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT65), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n467), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR3_X1   g053(.A1(new_n466), .A2(new_n468), .A3(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n476), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g058(.A(G2105), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n483), .B1(G124), .B2(new_n485), .ZN(G162));
  NOR3_X1   g061(.A1(new_n461), .A2(KEYINPUT65), .A3(KEYINPUT3), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n472), .B1(new_n459), .B2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n460), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G126), .A4(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT67), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n488), .A2(new_n460), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n497), .A2(G138), .A3(new_n467), .A4(new_n473), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n498), .A2(KEYINPUT4), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n496), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT68), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n506), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT69), .B(G88), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n512), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT70), .Z(new_n523));
  INV_X1    g098(.A(new_n514), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n513), .A2(KEYINPUT71), .A3(G543), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n527), .A2(G51), .A3(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n521), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n522), .B(KEYINPUT70), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n529), .A2(new_n532), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT73), .A4(new_n525), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n509), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n543));
  OAI21_X1  g118(.A(G651), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n543), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n527), .A2(new_n528), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n514), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n540), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n527), .A2(G43), .A3(new_n528), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n524), .A2(G81), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n517), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n517), .B2(new_n564), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n524), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n509), .B2(G65), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  AOI211_X1 g148(.A(KEYINPUT75), .B(new_n569), .C1(new_n509), .C2(G65), .ZN(new_n574));
  NOR3_X1   g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n506), .A2(new_n508), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(G65), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(new_n568), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n511), .B1(new_n579), .B2(KEYINPUT75), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  AOI21_X1  g156(.A(KEYINPUT76), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n567), .B1(new_n575), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  AND2_X1   g159(.A1(new_n534), .A2(new_n537), .ZN(G286));
  NAND2_X1  g160(.A1(new_n524), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n513), .A2(G49), .A3(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n511), .ZN(new_n591));
  INV_X1    g166(.A(G86), .ZN(new_n592));
  INV_X1    g167(.A(G48), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n514), .A2(new_n592), .B1(new_n593), .B2(new_n517), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n524), .A2(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n511), .B2(new_n598), .C1(new_n599), .C2(new_n546), .ZN(G290));
  NAND3_X1  g175(.A1(new_n527), .A2(G54), .A3(new_n528), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n509), .A2(G66), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n511), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n601), .B(new_n607), .C1(new_n511), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n509), .A2(G92), .A3(new_n513), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(G171), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(new_n616), .B2(G171), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n616), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n616), .B2(G168), .ZN(G280));
  AOI22_X1  g197(.A1(new_n606), .A2(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(G148));
  NAND3_X1  g200(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(new_n616), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n615), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g205(.A(KEYINPUT66), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n461), .B2(G2105), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n467), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n499), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n485), .A2(G123), .ZN(new_n639));
  INV_X1    g214(.A(new_n476), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n467), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n639), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT16), .B(G1341), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(G14), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n652), .A2(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT17), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT78), .Z(new_n667));
  INV_X1    g242(.A(new_n662), .ZN(new_n668));
  INV_X1    g243(.A(new_n664), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n662), .B2(new_n664), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n663), .B2(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n667), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT79), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(new_n682), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n683), .B1(KEYINPUT20), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n680), .A2(new_n684), .A3(new_n682), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(KEYINPUT20), .C2(new_n685), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1991), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n691), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(G229));
  NOR2_X1   g274(.A1(G16), .A2(G22), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G166), .B2(G16), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT82), .B(G1971), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G6), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n595), .B2(new_n704), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n703), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT34), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n640), .A2(G131), .ZN(new_n716));
  NOR3_X1   g291(.A1(KEYINPUT80), .A2(G95), .A3(G2105), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT80), .B1(G95), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G119), .B2(new_n485), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT81), .ZN(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT35), .B(G1991), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G24), .B(G290), .S(G16), .Z(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1986), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n715), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT36), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n704), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n557), .B2(new_n704), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT83), .Z(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n704), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n704), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT90), .B(G1966), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT92), .Z(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n740), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT93), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n740), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n740), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2078), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n745), .B2(KEYINPUT93), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n734), .A2(new_n739), .A3(new_n746), .A4(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n740), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G140), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n467), .A2(G116), .ZN(new_n756));
  OAI21_X1  g331(.A(KEYINPUT84), .B1(G104), .B2(G2105), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n756), .A2(G2104), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(KEYINPUT84), .A2(G104), .A3(G2105), .ZN(new_n759));
  OAI22_X1  g334(.A1(new_n476), .A2(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G128), .B2(new_n485), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n754), .B1(new_n761), .B2(new_n740), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT31), .B(G11), .Z(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n740), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n740), .B1(KEYINPUT24), .B2(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(KEYINPUT24), .B2(G34), .ZN(new_n768));
  INV_X1    g343(.A(G160), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G2084), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n766), .B1(new_n740), .B2(new_n644), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n763), .B(new_n772), .C1(new_n771), .C2(new_n770), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n640), .A2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n485), .A2(G129), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n634), .A2(G105), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n775), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT89), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT27), .B(G1996), .Z(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NOR2_X1   g361(.A1(G5), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G171), .B2(G16), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G1961), .ZN(new_n789));
  AOI22_X1  g364(.A1(G1961), .A2(new_n788), .B1(new_n743), .B2(new_n744), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n773), .A2(new_n786), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  INV_X1    g368(.A(G139), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n476), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT86), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n499), .A2(G127), .ZN(new_n799));
  INV_X1    g374(.A(G115), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n461), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n797), .A2(new_n798), .B1(G2105), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G29), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G29), .B2(G33), .ZN(new_n804));
  INV_X1    g379(.A(G2072), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT88), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT87), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n751), .A2(new_n791), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n704), .A2(G20), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n566), .ZN(new_n812));
  INV_X1    g387(.A(G91), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n514), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n573), .B1(new_n572), .B2(new_n574), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n580), .A2(KEYINPUT76), .A3(new_n581), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(KEYINPUT23), .B(new_n811), .C1(new_n817), .C2(new_n704), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(KEYINPUT23), .B2(new_n811), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1956), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n704), .A2(G4), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n623), .B2(new_n704), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n736), .A2(new_n737), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT91), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n810), .A2(new_n820), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n730), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n829));
  XNOR2_X1  g404(.A(G311), .B(new_n829), .ZN(G150));
  NAND2_X1  g405(.A1(new_n623), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n546), .A2(new_n834), .B1(new_n835), .B2(new_n514), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n837), .A2(new_n511), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n557), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n836), .A2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n626), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n833), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G860), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n833), .A2(new_n843), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n841), .A2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(G145));
  NAND2_X1  g425(.A1(new_n640), .A2(G142), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n467), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G130), .B2(new_n485), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(new_n636), .Z(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n722), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n802), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n783), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G164), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n761), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n761), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G162), .B(KEYINPUT95), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n644), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n769), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n864), .A2(new_n858), .A3(new_n865), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT97), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n869), .B1(new_n874), .B2(new_n866), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  NOR3_X1   g454(.A1(G299), .A2(new_n623), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT98), .B1(new_n615), .B2(new_n817), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n623), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n628), .B(new_n843), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT99), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n879), .B1(G299), .B2(new_n623), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n615), .A2(new_n817), .A3(KEYINPUT98), .ZN(new_n889));
  AND4_X1   g464(.A1(KEYINPUT41), .A2(new_n888), .A3(new_n889), .A4(new_n883), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT100), .B1(new_n880), .B2(new_n881), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n883), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n887), .B1(new_n896), .B2(new_n885), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n886), .B1(new_n897), .B2(KEYINPUT99), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(new_n710), .ZN(new_n899));
  XNOR2_X1  g474(.A(G303), .B(new_n595), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n903), .B2(new_n898), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g484(.A(new_n908), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  OAI21_X1  g486(.A(G301), .B1(G168), .B2(KEYINPUT103), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n843), .A2(G168), .A3(KEYINPUT103), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n843), .B1(KEYINPUT103), .B2(G168), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n840), .B(new_n842), .C1(G286), .C2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G171), .B1(G286), .B2(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n913), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n911), .B1(new_n896), .B2(new_n921), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n916), .A2(new_n920), .B1(new_n882), .B2(new_n883), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n893), .A2(new_n883), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n892), .B1(new_n888), .B2(new_n889), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n895), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n890), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n916), .A2(new_n920), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n901), .B(new_n922), .C1(new_n930), .C2(new_n911), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n901), .B(KEYINPUT105), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n896), .A2(new_n921), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT104), .B1(new_n936), .B2(new_n923), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n935), .B1(new_n937), .B2(new_n922), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n933), .A2(new_n938), .A3(KEYINPUT43), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n923), .B(KEYINPUT106), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n942));
  AOI211_X1 g517(.A(new_n942), .B(new_n921), .C1(KEYINPUT41), .C2(new_n894), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n934), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n944), .A2(new_n932), .A3(new_n931), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n939), .B(KEYINPUT44), .C1(new_n940), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n933), .B2(new_n938), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n944), .A2(new_n940), .A3(new_n932), .A4(new_n931), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT107), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  AOI211_X1 g527(.A(new_n952), .B(KEYINPUT44), .C1(new_n947), .C2(new_n948), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n946), .B1(new_n951), .B2(new_n953), .ZN(G397));
  INV_X1    g529(.A(KEYINPUT114), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n496), .B2(new_n502), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(G160), .B2(G40), .ZN(new_n960));
  INV_X1    g535(.A(new_n464), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n499), .B2(G125), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT64), .B1(new_n962), .B2(new_n467), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n465), .A2(new_n458), .A3(G2105), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G40), .ZN(new_n966));
  NOR4_X1   g541(.A1(new_n965), .A2(KEYINPUT109), .A3(new_n966), .A4(new_n478), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n958), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT113), .B(G8), .Z(new_n969));
  AOI21_X1  g544(.A(new_n955), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G101), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n632), .B2(new_n633), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n640), .B2(G137), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(G40), .A3(new_n963), .A4(new_n964), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n466), .A2(new_n468), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(new_n959), .A3(G40), .A4(new_n973), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n957), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n969), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(KEYINPUT114), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n970), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n982));
  NAND3_X1  g557(.A1(G305), .A2(new_n982), .A3(G1981), .ZN(new_n983));
  INV_X1    g558(.A(G1981), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT49), .B1(new_n595), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n595), .A2(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n983), .A2(new_n990), .A3(new_n985), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n981), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n975), .A2(new_n977), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT45), .B(new_n956), .C1(new_n496), .C2(new_n502), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n957), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n956), .C1(new_n496), .C2(new_n502), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n957), .A2(KEYINPUT50), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(G2090), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT55), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1008), .A3(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(KEYINPUT116), .A2(G1976), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(KEYINPUT116), .A2(G1976), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT52), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(G288), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1976), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G288), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n968), .A2(new_n955), .A3(new_n969), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT114), .B1(new_n978), .B2(new_n979), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(KEYINPUT115), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1015), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1022), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1017), .B(new_n1024), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n993), .B(new_n1009), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1008), .B1(new_n1005), .B2(new_n969), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT124), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n981), .A2(new_n992), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n970), .A2(new_n980), .B1(new_n1016), .B2(G288), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1014), .B1(new_n1030), .B2(new_n1024), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT124), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1027), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1009), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G299), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n817), .A2(KEYINPUT57), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1956), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1004), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n975), .A2(new_n977), .B1(new_n957), .B2(new_n996), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT120), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n995), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1041), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1041), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1049));
  INV_X1    g624(.A(G2067), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1004), .A2(new_n823), .B1(new_n1050), .B2(new_n978), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n615), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1048), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT58), .B(G1341), .Z(new_n1054));
  NAND2_X1  g629(.A1(new_n968), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n1056));
  INV_X1    g631(.A(G1996), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n994), .A2(new_n997), .A3(new_n1057), .A4(new_n995), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n557), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1051), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n615), .B1(new_n1051), .B2(KEYINPUT60), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1065), .A2(new_n1066), .B1(KEYINPUT60), .B2(new_n1051), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1049), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1069), .B2(new_n1048), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1041), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(KEYINPUT61), .A3(new_n1049), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1064), .A2(new_n1067), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(KEYINPUT122), .B(new_n557), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT59), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1058), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1054), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n978), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT121), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT122), .B1(new_n1083), .B2(new_n557), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1053), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  INV_X1    g662(.A(G2078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n994), .A2(new_n997), .A3(new_n1088), .A4(new_n995), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n957), .A2(KEYINPUT108), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT108), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n956), .C1(new_n496), .C2(new_n502), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n996), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1088), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1096), .B(new_n478), .C1(G2105), .C2(new_n465), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n995), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT123), .B(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1004), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1091), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1087), .B1(new_n1101), .B2(G171), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1090), .A2(new_n1089), .B1(new_n1004), .B2(new_n1099), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1044), .A2(KEYINPUT53), .A3(new_n1088), .A4(new_n995), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(KEYINPUT125), .A3(G301), .A4(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1091), .A2(new_n1100), .A3(new_n1104), .A4(G301), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(G301), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1110));
  AND4_X1   g685(.A1(G301), .A2(new_n1091), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1087), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n737), .B1(new_n1044), .B2(new_n995), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1114), .A2(new_n1115), .B1(G2084), .B2(new_n1004), .ZN(new_n1116));
  INV_X1    g691(.A(new_n737), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n998), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(KEYINPUT118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n969), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G168), .A2(new_n979), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1118), .A2(KEYINPUT118), .B1(new_n1124), .B2(new_n771), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n1127), .B2(G8), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1123), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1121), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1113), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1037), .A2(new_n1086), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n993), .A2(new_n1016), .A3(new_n710), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n981), .B1(new_n1134), .B2(new_n988), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1009), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(new_n1033), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1133), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1120), .A2(G286), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1005), .A2(G8), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT63), .B1(new_n1141), .B2(new_n1008), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1140), .A2(new_n1026), .A3(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1033), .A2(new_n1139), .A3(new_n1035), .A4(new_n1009), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n1144), .B2(KEYINPUT119), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1026), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1146), .A2(new_n1147), .A3(new_n1035), .A4(new_n1139), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1030), .A2(new_n1024), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1032), .A3(new_n1015), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(new_n1035), .A3(new_n1009), .A4(new_n993), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1140), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1148), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1143), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1133), .A4(new_n1137), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1110), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(KEYINPUT62), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1037), .C1(KEYINPUT62), .C2(new_n1162), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1150), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1095), .B1(new_n977), .B2(new_n975), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT110), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n761), .B(new_n1050), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT111), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n861), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1166), .A2(new_n1057), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1171), .A2(new_n1172), .B1(new_n1057), .B2(new_n861), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1167), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n722), .B(new_n724), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT112), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(G290), .B(G1986), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1178), .B1(new_n1166), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1165), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1172), .B(KEYINPUT46), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1182), .A2(new_n1171), .A3(new_n1169), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G290), .A2(G1986), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1166), .A2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT48), .Z(new_n1187));
  OAI21_X1  g762(.A(new_n1184), .B1(new_n1178), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n722), .A2(new_n724), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1174), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n761), .A2(new_n1050), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1175), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1188), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1181), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g769(.A(G319), .B1(new_n659), .B2(new_n660), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g771(.A1(new_n694), .A2(new_n698), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n1199));
  XNOR2_X1  g773(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  AND3_X1   g774(.A1(new_n1200), .A2(new_n877), .A3(new_n949), .ZN(G308));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n877), .A3(new_n949), .ZN(G225));
endmodule


