

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X2 U555 ( .A1(G2105), .A2(n525), .ZN(n885) );
  NOR2_X2 U556 ( .A1(n1002), .A2(n640), .ZN(n654) );
  OR2_X2 U557 ( .A1(n635), .A2(n634), .ZN(n683) );
  NOR2_X1 U558 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U559 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U560 ( .A(n592), .B(KEYINPUT86), .ZN(n635) );
  AND2_X1 U561 ( .A1(n735), .A2(n734), .ZN(n736) );
  BUF_X1 U562 ( .A(n683), .Z(n694) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n731), .ZN(n709) );
  NOR2_X1 U564 ( .A1(n710), .A2(n709), .ZN(n711) );
  AND2_X1 U565 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U566 ( .A1(G651), .A2(n558), .ZN(n531) );
  XNOR2_X1 U567 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n522) );
  NOR2_X1 U568 ( .A1(n737), .A2(n736), .ZN(n739) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n799) );
  NOR2_X2 U570 ( .A1(n526), .A2(n525), .ZN(n889) );
  XNOR2_X1 U571 ( .A(KEYINPUT73), .B(n632), .ZN(n1002) );
  NAND2_X1 U572 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U573 ( .A1(n591), .A2(n590), .ZN(n756) );
  BUF_X1 U574 ( .A(n756), .Z(G160) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X2 U576 ( .A(n522), .B(n521), .ZN(n884) );
  NAND2_X1 U577 ( .A1(G138), .A2(n884), .ZN(n524) );
  INV_X1 U578 ( .A(G2104), .ZN(n525) );
  NAND2_X1 U579 ( .A1(G102), .A2(n885), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n524), .A2(n523), .ZN(n530) );
  INV_X1 U581 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U582 ( .A1(G114), .A2(n889), .ZN(n528) );
  NOR2_X1 U583 ( .A1(G2104), .A2(n526), .ZN(n890) );
  NAND2_X1 U584 ( .A1(G126), .A2(n890), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n530), .A2(n529), .ZN(G164) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n558) );
  XOR2_X1 U588 ( .A(KEYINPUT65), .B(n531), .Z(n794) );
  NAND2_X1 U589 ( .A1(G52), .A2(n794), .ZN(n534) );
  INV_X1 U590 ( .A(G651), .ZN(n535) );
  NOR2_X1 U591 ( .A1(G543), .A2(n535), .ZN(n532) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n532), .Z(n795) );
  NAND2_X1 U593 ( .A1(G64), .A2(n795), .ZN(n533) );
  AND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT72), .B(KEYINPUT9), .ZN(n539) );
  NOR2_X1 U596 ( .A1(n558), .A2(n535), .ZN(n798) );
  NAND2_X1 U597 ( .A1(G77), .A2(n798), .ZN(n537) );
  NAND2_X1 U598 ( .A1(G90), .A2(n799), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U600 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(G301) );
  NAND2_X1 U602 ( .A1(n799), .A2(G89), .ZN(n542) );
  XNOR2_X1 U603 ( .A(n542), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G76), .A2(n798), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT5), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G51), .A2(n794), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G63), .A2(n795), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n548), .Z(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U612 ( .A(n551), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G75), .A2(n798), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G88), .A2(n799), .ZN(n552) );
  NAND2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G50), .A2(n794), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G62), .A2(n795), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U620 ( .A1(n557), .A2(n556), .ZN(G166) );
  NAND2_X1 U621 ( .A1(n558), .A2(G87), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G49), .A2(n794), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G74), .A2(G651), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n795), .A2(n561), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(KEYINPUT81), .B(n564), .Z(G288) );
  INV_X1 U628 ( .A(G166), .ZN(G303) );
  NAND2_X1 U629 ( .A1(G73), .A2(n798), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT2), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT82), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G86), .A2(n799), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G48), .A2(n794), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G61), .A2(n795), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT83), .B(n573), .ZN(G305) );
  NAND2_X1 U639 ( .A1(n798), .A2(G72), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT70), .B(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n799), .A2(G85), .ZN(n575) );
  XOR2_X1 U642 ( .A(KEYINPUT69), .B(n575), .Z(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(KEYINPUT71), .B(n578), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G47), .A2(n794), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G60), .A2(n795), .ZN(n579) );
  AND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(G290) );
  NAND2_X1 U649 ( .A1(n884), .A2(G137), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n889), .A2(G113), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n585), .B(KEYINPUT68), .ZN(n591) );
  XOR2_X1 U653 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n587) );
  NAND2_X1 U654 ( .A1(G101), .A2(n885), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n587), .B(n586), .ZN(n589) );
  NAND2_X1 U656 ( .A1(n890), .A2(G125), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n756), .A2(G40), .ZN(n592) );
  NOR2_X1 U659 ( .A1(G164), .A2(G1384), .ZN(n633) );
  NOR2_X1 U660 ( .A1(n635), .A2(n633), .ZN(n751) );
  NAND2_X1 U661 ( .A1(G140), .A2(n884), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G104), .A2(n885), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT34), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT87), .ZN(n602) );
  XNOR2_X1 U666 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G116), .A2(n889), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G128), .A2(n890), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U672 ( .A(KEYINPUT36), .B(n603), .Z(n898) );
  XNOR2_X1 U673 ( .A(KEYINPUT37), .B(G2067), .ZN(n748) );
  NOR2_X1 U674 ( .A1(n898), .A2(n748), .ZN(n928) );
  NAND2_X1 U675 ( .A1(n751), .A2(n928), .ZN(n746) );
  NAND2_X1 U676 ( .A1(G107), .A2(n889), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G119), .A2(n890), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G131), .A2(n884), .ZN(n606) );
  XNOR2_X1 U680 ( .A(KEYINPUT89), .B(n606), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n885), .A2(G95), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n876) );
  NAND2_X1 U684 ( .A1(G1991), .A2(n876), .ZN(n621) );
  NAND2_X1 U685 ( .A1(G117), .A2(n889), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT90), .B(n611), .Z(n614) );
  NAND2_X1 U687 ( .A1(n885), .A2(G105), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT38), .B(n612), .Z(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n890), .A2(G129), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT91), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G141), .A2(n884), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n875) );
  NAND2_X1 U695 ( .A1(G1996), .A2(n875), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U697 ( .A(KEYINPUT92), .B(n622), .ZN(n931) );
  NAND2_X1 U698 ( .A1(n751), .A2(n931), .ZN(n740) );
  NAND2_X1 U699 ( .A1(n746), .A2(n740), .ZN(n737) );
  NAND2_X1 U700 ( .A1(n799), .A2(G81), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT12), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G68), .A2(n798), .ZN(n624) );
  NAND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(KEYINPUT13), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n794), .A2(G43), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n795), .A2(G56), .ZN(n629) );
  XOR2_X1 U708 ( .A(KEYINPUT14), .B(n629), .Z(n630) );
  NOR2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U710 ( .A(n633), .ZN(n634) );
  INV_X2 U711 ( .A(n683), .ZN(n676) );
  NAND2_X1 U712 ( .A1(G1996), .A2(n676), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n636), .B(KEYINPUT26), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G1341), .A2(n683), .ZN(n637) );
  XOR2_X1 U715 ( .A(n637), .B(KEYINPUT97), .Z(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G79), .A2(n798), .ZN(n642) );
  NAND2_X1 U718 ( .A1(G54), .A2(n794), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G92), .A2(n799), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G66), .A2(n795), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U723 ( .A(KEYINPUT77), .B(n645), .Z(n646) );
  NOR2_X1 U724 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT15), .B(n648), .ZN(n790) );
  INV_X1 U726 ( .A(n790), .ZN(n997) );
  NAND2_X1 U727 ( .A1(n654), .A2(n997), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n676), .A2(G2067), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G1348), .A2(n694), .ZN(n649) );
  NAND2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(KEYINPUT98), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n653), .A2(n652), .ZN(n657) );
  INV_X1 U733 ( .A(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n655), .A2(n790), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G53), .A2(n794), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G65), .A2(n795), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U739 ( .A1(G78), .A2(n798), .ZN(n661) );
  NAND2_X1 U740 ( .A1(G91), .A2(n799), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n994) );
  NAND2_X1 U743 ( .A1(n676), .A2(G2072), .ZN(n664) );
  XNOR2_X1 U744 ( .A(KEYINPUT27), .B(n664), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT95), .B(G1956), .Z(n950) );
  NAND2_X1 U746 ( .A1(n950), .A2(n683), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT96), .B(n665), .Z(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n994), .A2(n670), .ZN(n668) );
  NAND2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U751 ( .A1(n670), .A2(n994), .ZN(n671) );
  XOR2_X1 U752 ( .A(n671), .B(KEYINPUT28), .Z(n672) );
  NAND2_X1 U753 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n674), .B(KEYINPUT29), .ZN(n680) );
  XOR2_X1 U755 ( .A(G2078), .B(KEYINPUT25), .Z(n974) );
  NOR2_X1 U756 ( .A1(n974), .A2(n694), .ZN(n675) );
  XNOR2_X1 U757 ( .A(n675), .B(KEYINPUT94), .ZN(n678) );
  NOR2_X1 U758 ( .A1(n676), .A2(G1961), .ZN(n677) );
  NOR2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U760 ( .A1(G301), .A2(n682), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n681), .B(KEYINPUT99), .ZN(n692) );
  AND2_X1 U763 ( .A1(G301), .A2(n682), .ZN(n688) );
  NAND2_X1 U764 ( .A1(G8), .A2(n683), .ZN(n731) );
  NOR2_X1 U765 ( .A1(G2084), .A2(n694), .ZN(n705) );
  NOR2_X1 U766 ( .A1(n709), .A2(n705), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G8), .A2(n684), .ZN(n685) );
  XNOR2_X1 U768 ( .A(KEYINPUT30), .B(n685), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n686), .A2(G168), .ZN(n687) );
  XOR2_X1 U770 ( .A(n689), .B(KEYINPUT100), .Z(n690) );
  XNOR2_X1 U771 ( .A(KEYINPUT31), .B(n690), .ZN(n691) );
  NAND2_X1 U772 ( .A1(n692), .A2(n691), .ZN(n708) );
  AND2_X1 U773 ( .A1(G286), .A2(G8), .ZN(n693) );
  NAND2_X1 U774 ( .A1(n708), .A2(n693), .ZN(n703) );
  INV_X1 U775 ( .A(G8), .ZN(n701) );
  NOR2_X1 U776 ( .A1(G1971), .A2(n731), .ZN(n696) );
  NOR2_X1 U777 ( .A1(G2090), .A2(n694), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U779 ( .A(KEYINPUT102), .B(n697), .Z(n698) );
  NOR2_X1 U780 ( .A1(G166), .A2(n698), .ZN(n699) );
  XNOR2_X1 U781 ( .A(n699), .B(KEYINPUT103), .ZN(n700) );
  OR2_X1 U782 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U783 ( .A(n704), .B(KEYINPUT32), .ZN(n713) );
  NAND2_X1 U784 ( .A1(G8), .A2(n705), .ZN(n706) );
  XOR2_X1 U785 ( .A(KEYINPUT93), .B(n706), .Z(n707) );
  NAND2_X1 U786 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U787 ( .A(n711), .B(KEYINPUT101), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n725) );
  NOR2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n720) );
  NOR2_X1 U790 ( .A1(G1971), .A2(G303), .ZN(n714) );
  NOR2_X1 U791 ( .A1(n720), .A2(n714), .ZN(n993) );
  NAND2_X1 U792 ( .A1(n725), .A2(n993), .ZN(n717) );
  NAND2_X1 U793 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  INV_X1 U794 ( .A(n1000), .ZN(n715) );
  NOR2_X1 U795 ( .A1(n715), .A2(n731), .ZN(n716) );
  XNOR2_X1 U796 ( .A(n718), .B(KEYINPUT64), .ZN(n719) );
  NOR2_X1 U797 ( .A1(KEYINPUT33), .A2(n719), .ZN(n723) );
  NAND2_X1 U798 ( .A1(n720), .A2(KEYINPUT33), .ZN(n721) );
  NOR2_X1 U799 ( .A1(n721), .A2(n731), .ZN(n722) );
  XOR2_X1 U800 ( .A(G1981), .B(G305), .Z(n989) );
  NAND2_X1 U801 ( .A1(n724), .A2(n989), .ZN(n735) );
  NOR2_X1 U802 ( .A1(G2090), .A2(G303), .ZN(n726) );
  NAND2_X1 U803 ( .A1(G8), .A2(n726), .ZN(n727) );
  NAND2_X1 U804 ( .A1(n725), .A2(n727), .ZN(n728) );
  AND2_X1 U805 ( .A1(n728), .A2(n731), .ZN(n733) );
  NOR2_X1 U806 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XOR2_X1 U807 ( .A(n729), .B(KEYINPUT24), .Z(n730) );
  NOR2_X1 U808 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U809 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U810 ( .A(G1986), .B(G290), .ZN(n1008) );
  NAND2_X1 U811 ( .A1(n1008), .A2(n751), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n754) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n875), .ZN(n915) );
  INV_X1 U814 ( .A(n740), .ZN(n743) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n876), .ZN(n918) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U817 ( .A1(n918), .A2(n741), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U819 ( .A1(n915), .A2(n744), .ZN(n745) );
  XNOR2_X1 U820 ( .A(KEYINPUT39), .B(n745), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n748), .A2(n898), .ZN(n749) );
  XNOR2_X1 U823 ( .A(n749), .B(KEYINPUT104), .ZN(n933) );
  NAND2_X1 U824 ( .A1(n750), .A2(n933), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n755), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U827 ( .A(G2435), .B(G2446), .Z(n758) );
  XNOR2_X1 U828 ( .A(KEYINPUT105), .B(G2451), .ZN(n757) );
  XNOR2_X1 U829 ( .A(n758), .B(n757), .ZN(n759) );
  XOR2_X1 U830 ( .A(n759), .B(G2430), .Z(n761) );
  XNOR2_X1 U831 ( .A(G1348), .B(G1341), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n761), .B(n760), .ZN(n765) );
  XOR2_X1 U833 ( .A(G2438), .B(KEYINPUT107), .Z(n763) );
  XNOR2_X1 U834 ( .A(KEYINPUT106), .B(G2454), .ZN(n762) );
  XNOR2_X1 U835 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U836 ( .A(n765), .B(n764), .Z(n767) );
  XNOR2_X1 U837 ( .A(G2443), .B(G2427), .ZN(n766) );
  XNOR2_X1 U838 ( .A(n767), .B(n766), .ZN(n768) );
  AND2_X1 U839 ( .A1(n768), .A2(G14), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U841 ( .A1(G123), .A2(n890), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n769), .B(KEYINPUT78), .ZN(n770) );
  XNOR2_X1 U843 ( .A(n770), .B(KEYINPUT18), .ZN(n772) );
  NAND2_X1 U844 ( .A1(G111), .A2(n889), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U846 ( .A1(G135), .A2(n884), .ZN(n774) );
  NAND2_X1 U847 ( .A1(G99), .A2(n885), .ZN(n773) );
  NAND2_X1 U848 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U849 ( .A1(n776), .A2(n775), .ZN(n917) );
  XNOR2_X1 U850 ( .A(n917), .B(G2096), .ZN(n777) );
  XNOR2_X1 U851 ( .A(n777), .B(KEYINPUT79), .ZN(n778) );
  OR2_X1 U852 ( .A1(G2100), .A2(n778), .ZN(G156) );
  INV_X1 U853 ( .A(n994), .ZN(G299) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  INV_X1 U856 ( .A(G82), .ZN(G220) );
  NAND2_X1 U857 ( .A1(G7), .A2(G661), .ZN(n779) );
  XOR2_X1 U858 ( .A(n779), .B(KEYINPUT10), .Z(n833) );
  NAND2_X1 U859 ( .A1(n833), .A2(G567), .ZN(n780) );
  XOR2_X1 U860 ( .A(KEYINPUT11), .B(n780), .Z(G234) );
  XOR2_X1 U861 ( .A(G860), .B(KEYINPUT74), .Z(n787) );
  NOR2_X1 U862 ( .A1(n1002), .A2(n787), .ZN(n781) );
  XNOR2_X1 U863 ( .A(n781), .B(KEYINPUT75), .ZN(G153) );
  NAND2_X1 U864 ( .A1(G301), .A2(G868), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT76), .ZN(n784) );
  INV_X1 U866 ( .A(G868), .ZN(n817) );
  NAND2_X1 U867 ( .A1(n817), .A2(n790), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n784), .A2(n783), .ZN(G284) );
  NOR2_X1 U869 ( .A1(G286), .A2(n817), .ZN(n786) );
  NOR2_X1 U870 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(G297) );
  NAND2_X1 U872 ( .A1(n787), .A2(G559), .ZN(n788) );
  NAND2_X1 U873 ( .A1(n788), .A2(n997), .ZN(n789) );
  XNOR2_X1 U874 ( .A(n789), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U875 ( .A1(G559), .A2(n790), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n791), .A2(G868), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n1002), .A2(n817), .ZN(n792) );
  NAND2_X1 U878 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U879 ( .A1(G55), .A2(n794), .ZN(n797) );
  NAND2_X1 U880 ( .A1(G67), .A2(n795), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n803) );
  NAND2_X1 U882 ( .A1(G80), .A2(n798), .ZN(n801) );
  NAND2_X1 U883 ( .A1(G93), .A2(n799), .ZN(n800) );
  NAND2_X1 U884 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U885 ( .A1(n803), .A2(n802), .ZN(n816) );
  XNOR2_X1 U886 ( .A(KEYINPUT80), .B(n1002), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n997), .A2(G559), .ZN(n814) );
  XNOR2_X1 U888 ( .A(n804), .B(n814), .ZN(n805) );
  NOR2_X1 U889 ( .A1(G860), .A2(n805), .ZN(n806) );
  XNOR2_X1 U890 ( .A(n816), .B(n806), .ZN(G145) );
  XNOR2_X1 U891 ( .A(G290), .B(n1002), .ZN(n813) );
  XOR2_X1 U892 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n807) );
  XNOR2_X1 U893 ( .A(G288), .B(n807), .ZN(n808) );
  XOR2_X1 U894 ( .A(G303), .B(n808), .Z(n811) );
  XOR2_X1 U895 ( .A(G299), .B(n816), .Z(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(G305), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U898 ( .A(n813), .B(n812), .ZN(n904) );
  XOR2_X1 U899 ( .A(n904), .B(n814), .Z(n815) );
  NOR2_X1 U900 ( .A1(n817), .A2(n815), .ZN(n819) );
  AND2_X1 U901 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U902 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U905 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XOR2_X1 U906 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n822) );
  XNOR2_X1 U907 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U908 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XNOR2_X1 U909 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n825) );
  XOR2_X1 U911 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U912 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G96), .A2(n827), .ZN(n838) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n838), .ZN(n831) );
  NAND2_X1 U915 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U916 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U917 ( .A1(G108), .A2(n829), .ZN(n837) );
  NAND2_X1 U918 ( .A1(G567), .A2(n837), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n840) );
  NAND2_X1 U920 ( .A1(G483), .A2(G661), .ZN(n832) );
  NOR2_X1 U921 ( .A1(n840), .A2(n832), .ZN(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U923 ( .A(G301), .ZN(G171) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U925 ( .A(n833), .ZN(G223) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U927 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  XOR2_X1 U935 ( .A(n839), .B(KEYINPUT108), .Z(G261) );
  INV_X1 U936 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U937 ( .A(KEYINPUT109), .B(n840), .ZN(G319) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2090), .Z(n844) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U944 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1981), .B(G1966), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n860) );
  XOR2_X1 U950 ( .A(KEYINPUT111), .B(G2474), .Z(n852) );
  XNOR2_X1 U951 ( .A(G1976), .B(KEYINPUT112), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(G1971), .B(G1956), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1961), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U957 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G124), .A2(n890), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n889), .A2(G112), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G136), .A2(n884), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G100), .A2(n885), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G139), .A2(n884), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G103), .A2(n885), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G115), .A2(n889), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G127), .A2(n890), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n919) );
  XNOR2_X1 U976 ( .A(n919), .B(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n879) );
  XNOR2_X1 U979 ( .A(n917), .B(KEYINPUT46), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U982 ( .A(G164), .B(G162), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n900) );
  NAND2_X1 U984 ( .A1(G142), .A2(n884), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G106), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n888), .B(KEYINPUT45), .ZN(n895) );
  NAND2_X1 U988 ( .A1(G118), .A2(n889), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT113), .B(n893), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U993 ( .A(G160), .B(n896), .ZN(n897) );
  XOR2_X1 U994 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G395) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(G286), .Z(n903) );
  XOR2_X1 U998 ( .A(G301), .B(n997), .Z(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(n907), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n908), .B(KEYINPUT49), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n909), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n910), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(KEYINPUT117), .B(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1012 ( .A(G2090), .B(G162), .Z(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1014 ( .A(KEYINPUT51), .B(n916), .Z(n930) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n926) );
  XOR2_X1 U1016 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n922), .Z(n924) );
  XOR2_X1 U1020 ( .A(G160), .B(G2084), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(n935) );
  INV_X1 U1025 ( .A(n931), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  XOR2_X1 U1029 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n985) );
  NAND2_X1 U1030 ( .A1(n937), .A2(n985), .ZN(n938) );
  NAND2_X1 U1031 ( .A1(n938), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G23), .B(G1976), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G1986), .B(G24), .Z(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n943) );
  XNOR2_X1 U1038 ( .A(n944), .B(n943), .ZN(n948) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G21), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G1961), .B(G5), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n960) );
  XNOR2_X1 U1043 ( .A(G1348), .B(KEYINPUT59), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n949), .B(G4), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n950), .B(G20), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G6), .B(G1981), .Z(n955) );
  XNOR2_X1 U1050 ( .A(KEYINPUT125), .B(n955), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1052 ( .A(n958), .B(KEYINPUT60), .Z(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1054 ( .A(KEYINPUT127), .B(n961), .Z(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT61), .B(n962), .ZN(n963) );
  INV_X1 U1056 ( .A(G16), .ZN(n988) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n988), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n964), .A2(G11), .ZN(n1018) );
  XNOR2_X1 U1059 ( .A(G25), .B(G1991), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT119), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G32), .B(G1996), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(G28), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT120), .B(G2072), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(G33), .B(n969), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G27), .B(n974), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1071 ( .A(KEYINPUT53), .B(n977), .Z(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT54), .B(G34), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT121), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(G2084), .B(n979), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G35), .B(G2090), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n985), .B(n984), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(G29), .A2(n986), .ZN(n987) );
  XOR2_X1 U1080 ( .A(KEYINPUT122), .B(n987), .Z(n1016) );
  XOR2_X1 U1081 ( .A(n988), .B(KEYINPUT56), .Z(n1013) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT57), .B(n991), .ZN(n1011) );
  NAND2_X1 U1085 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1087 ( .A(G1956), .B(n994), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1006) );
  XOR2_X1 U1089 ( .A(G171), .B(G1961), .Z(n999) );
  XOR2_X1 U1090 ( .A(n997), .B(G1348), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G1341), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT123), .B(n1009), .Z(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(n1014), .B(KEYINPUT124), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1021), .ZN(G150) );
  INV_X1 U1105 ( .A(G150), .ZN(G311) );
endmodule

