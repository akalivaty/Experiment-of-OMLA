//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT9), .B(G234), .Z(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n191), .B(KEYINPUT72), .Z(new_n192));
  AND2_X1   g006(.A1(KEYINPUT73), .A2(G104), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT73), .A2(G104), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G107), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT74), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n196), .A3(G104), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT73), .A2(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT73), .A2(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n196), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(KEYINPUT3), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n200), .A2(new_n201), .A3(new_n206), .A4(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n198), .B1(new_n209), .B2(G101), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT64), .A2(G146), .ZN(new_n213));
  OAI21_X1  g027(.A(G143), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT64), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT64), .A2(G146), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n215), .A2(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n218), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n220), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n221), .A2(new_n223), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n233), .B2(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n218), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n220), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n198), .B(new_n236), .C1(new_n209), .C2(G101), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n211), .A2(new_n232), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(G137), .ZN(new_n242));
  INV_X1    g056(.A(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT11), .A3(G134), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n244), .A3(new_n247), .A4(new_n242), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT75), .A2(KEYINPUT4), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n209), .A2(G101), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n209), .A2(G101), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n209), .B2(G101), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n218), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n214), .A2(new_n217), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n214), .A2(KEYINPUT65), .A3(new_n217), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n218), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n224), .B2(new_n225), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n264), .A2(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n238), .B(new_n253), .C1(new_n259), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n238), .B1(new_n259), .B2(new_n269), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n252), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n258), .A2(new_n257), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n209), .A2(G101), .A3(new_n255), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n237), .A2(new_n231), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(KEYINPUT74), .B1(G107), .B2(new_n207), .ZN(new_n279));
  INV_X1    g093(.A(G101), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n201), .A4(new_n206), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n229), .A4(new_n198), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n271), .B(new_n252), .C1(new_n276), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n270), .B1(new_n273), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n287));
  XNOR2_X1  g101(.A(G110), .B(G140), .ZN(new_n288));
  INV_X1    g102(.A(G227), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(G953), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n288), .B(new_n290), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n276), .A2(new_n283), .A3(new_n252), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n252), .B1(new_n276), .B2(new_n283), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT76), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n296), .B2(new_n284), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT79), .B1(new_n297), .B2(new_n291), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n294), .A2(new_n292), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n210), .A2(new_n230), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n253), .B1(new_n300), .B2(new_n237), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT78), .B(G469), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n304), .A2(new_n190), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n299), .B1(new_n273), .B2(new_n285), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT12), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n301), .B(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n292), .B1(new_n309), .B2(new_n294), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G469), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT77), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n270), .A2(new_n291), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n284), .B2(new_n296), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n291), .B1(new_n302), .B2(new_n270), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n190), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(G469), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n192), .B1(new_n306), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G214), .B1(G237), .B2(G902), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G210), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G110), .B(G122), .Z(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT8), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G113), .ZN(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G119), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(KEYINPUT5), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G116), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT2), .B(G113), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n331), .A2(new_n334), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n281), .A2(new_n198), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n281), .B2(new_n198), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n328), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(KEYINPUT82), .B(new_n328), .C1(new_n338), .C2(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n268), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n220), .C1(new_n227), .C2(new_n228), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G224), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT7), .B1(new_n350), .B2(G953), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n338), .ZN(new_n354));
  INV_X1    g168(.A(new_n326), .ZN(new_n355));
  INV_X1    g169(.A(new_n330), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(KEYINPUT67), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(new_n336), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n355), .C1(new_n259), .C2(new_n358), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n346), .A2(KEYINPUT80), .ZN(new_n360));
  INV_X1    g174(.A(new_n348), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT80), .B1(new_n346), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n350), .A2(G953), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT7), .B1(new_n363), .B2(KEYINPUT83), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(KEYINPUT83), .B2(new_n363), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n190), .B1(new_n353), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n274), .B2(new_n275), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n326), .B1(new_n369), .B2(new_n338), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n359), .A3(KEYINPUT6), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n363), .B(KEYINPUT81), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n360), .A2(new_n362), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n360), .B2(new_n362), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(new_n326), .C1(new_n369), .C2(new_n338), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n325), .B1(new_n368), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n367), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n342), .A2(new_n343), .B1(new_n349), .B2(new_n351), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n371), .A2(new_n375), .A3(new_n377), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n324), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n323), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  NOR2_X1   g200(.A1(G237), .A2(G953), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n388));
  AOI21_X1  g202(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n247), .ZN(new_n391));
  OAI21_X1  g205(.A(G131), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT17), .ZN(new_n394));
  XOR2_X1   g208(.A(G125), .B(G140), .Z(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n395), .A2(new_n396), .B1(G140), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n215), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n394), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT18), .A2(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n390), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT84), .ZN(new_n405));
  INV_X1    g219(.A(new_n395), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n233), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n215), .B2(new_n406), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n405), .B(new_n408), .C1(new_n390), .C2(new_n403), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(G104), .Z(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n386), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n402), .A2(new_n409), .A3(KEYINPUT87), .A4(new_n412), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n393), .A2(KEYINPUT85), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n398), .A2(new_n215), .ZN(new_n418));
  AND2_X1   g232(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n419));
  NOR2_X1   g233(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  MUX2_X1   g235(.A(new_n419), .B(new_n421), .S(new_n395), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n233), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n414), .A2(new_n415), .B1(new_n413), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT88), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(KEYINPUT20), .A3(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n414), .A2(new_n415), .B1(new_n413), .B2(new_n410), .ZN(new_n432));
  OAI21_X1  g246(.A(G475), .B1(new_n432), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n426), .B2(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT15), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G953), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n189), .A2(G217), .A3(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT94), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G122), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G116), .ZN(new_n446));
  AND2_X1   g260(.A1(KEYINPUT89), .A2(G122), .ZN(new_n447));
  NOR2_X1   g261(.A1(KEYINPUT89), .A2(G122), .ZN(new_n448));
  OAI21_X1  g262(.A(G116), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(KEYINPUT90), .B(G116), .C1(new_n447), .C2(new_n448), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(new_n196), .ZN(new_n454));
  XNOR2_X1  g268(.A(G128), .B(G143), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(G134), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(new_n452), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT14), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n446), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT92), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n465), .B(new_n462), .C1(new_n451), .C2(new_n452), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n446), .A2(new_n461), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n464), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n459), .B1(new_n469), .B2(new_n196), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT89), .B(G122), .ZN(new_n471));
  AOI21_X1  g285(.A(KEYINPUT90), .B1(new_n471), .B2(G116), .ZN(new_n472));
  INV_X1    g286(.A(new_n452), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n465), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n460), .A2(KEYINPUT92), .A3(new_n463), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n477), .A2(KEYINPUT93), .A3(G107), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n458), .B1(new_n470), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n455), .A2(new_n240), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n453), .A2(new_n196), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n454), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n240), .B1(new_n455), .B2(KEYINPUT13), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n222), .A2(G128), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(KEYINPUT13), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT91), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n444), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n477), .A2(KEYINPUT93), .A3(G107), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT93), .B1(new_n477), .B2(G107), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n457), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n487), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n443), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n493), .A3(new_n190), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n488), .A2(new_n493), .A3(KEYINPUT95), .A4(new_n190), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n440), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n439), .B1(new_n494), .B2(new_n495), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(G234), .A2(G237), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G952), .A3(new_n441), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT96), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(G902), .A3(G953), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n385), .A2(new_n437), .A3(new_n500), .A4(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n187), .B1(new_n321), .B2(new_n511), .ZN(new_n512));
  AND4_X1   g326(.A1(new_n500), .A2(new_n385), .A3(new_n437), .A4(new_n510), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n304), .A2(new_n190), .A3(new_n305), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n313), .A3(new_n319), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n513), .A2(KEYINPUT97), .A3(new_n192), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n333), .A2(G128), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(KEYINPUT70), .B2(KEYINPUT23), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(KEYINPUT70), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n218), .A2(G119), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n518), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G110), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n520), .ZN(new_n525));
  XOR2_X1   g339(.A(KEYINPUT24), .B(G110), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n399), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n523), .A2(G110), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(new_n418), .A3(new_n407), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT22), .B(G137), .ZN(new_n532));
  INV_X1    g346(.A(G234), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n188), .A2(new_n533), .A3(G953), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n532), .B(new_n534), .Z(new_n535));
  XNOR2_X1  g349(.A(new_n531), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n190), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(KEYINPUT25), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n538), .A2(KEYINPUT25), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n190), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n190), .A2(G234), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n539), .A2(new_n542), .A3(G217), .A4(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(G902), .B1(new_n533), .B2(G217), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  INV_X1    g362(.A(new_n358), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n268), .A2(new_n252), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n248), .B(KEYINPUT66), .ZN(new_n552));
  INV_X1    g366(.A(new_n242), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n240), .A2(G137), .ZN(new_n554));
  OAI21_X1  g368(.A(G131), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n229), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n551), .B1(new_n550), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n549), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n358), .A3(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n387), .A2(G210), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(new_n280), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n562), .B(new_n563), .Z(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n559), .A2(KEYINPUT31), .A3(new_n560), .A4(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n560), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n358), .B1(new_n550), .B2(new_n556), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT28), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT28), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n564), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT68), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n567), .B2(new_n568), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n581));
  INV_X1    g395(.A(new_n578), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n548), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n559), .A2(new_n560), .ZN(new_n586));
  INV_X1    g400(.A(new_n564), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n572), .A2(new_n574), .A3(new_n564), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n574), .A2(KEYINPUT69), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT69), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n560), .B2(new_n573), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n572), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n587), .A2(new_n589), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n190), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n585), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n547), .B1(new_n584), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n512), .A2(new_n516), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND3_X1  g417(.A1(new_n577), .A2(KEYINPUT68), .A3(new_n578), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n580), .B2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n321), .A2(new_n608), .A3(new_n547), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n382), .A2(new_n324), .A3(new_n383), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n324), .B1(new_n382), .B2(new_n383), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n322), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n509), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n488), .A2(new_n493), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n488), .A2(new_n493), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n190), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G478), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n494), .A2(G478), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n614), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT99), .B(new_n622), .C1(new_n620), .C2(G478), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n624), .A2(new_n625), .A3(new_n437), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n609), .A2(new_n613), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  NOR4_X1   g443(.A1(new_n612), .A2(new_n500), .A3(new_n509), .A4(new_n436), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n609), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(new_n535), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n531), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n545), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n544), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n606), .A2(new_n607), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n512), .A2(new_n516), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G110), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  OAI211_X1 g458(.A(new_n192), .B(new_n638), .C1(new_n306), .C2(new_n320), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n498), .A2(new_n499), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n503), .B(KEYINPUT101), .Z(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n508), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n646), .A2(new_n437), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT32), .B1(new_n604), .B2(new_n605), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n585), .A2(new_n599), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n385), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n645), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n218), .ZN(G30));
  OAI21_X1  g471(.A(new_n436), .B1(new_n498), .B2(new_n499), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n610), .A2(new_n611), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n659), .B(new_n660), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n650), .B(KEYINPUT39), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n321), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n658), .B(new_n661), .C1(new_n664), .C2(KEYINPUT40), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n638), .A2(new_n323), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n587), .B1(new_n570), .B2(new_n571), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n669), .A2(new_n565), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n584), .A2(new_n585), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT104), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n584), .A2(new_n675), .A3(new_n585), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n665), .A2(new_n666), .A3(new_n677), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NOR4_X1   g494(.A1(new_n624), .A2(new_n625), .A3(new_n437), .A4(new_n650), .ZN(new_n681));
  INV_X1    g495(.A(new_n192), .ZN(new_n682));
  INV_X1    g496(.A(new_n638), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n311), .A2(KEYINPUT77), .A3(new_n312), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n318), .B1(new_n317), .B2(G469), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n682), .B(new_n683), .C1(new_n686), .C2(new_n514), .ZN(new_n687));
  INV_X1    g501(.A(new_n655), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n681), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  NAND2_X1  g504(.A1(new_n304), .A2(new_n190), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n514), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n191), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n626), .A3(new_n601), .A4(new_n613), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n601), .A3(new_n630), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  AOI21_X1  g513(.A(new_n312), .B1(new_n304), .B2(new_n190), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n306), .A2(new_n700), .A3(new_n191), .A4(new_n612), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n584), .A2(new_n600), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n646), .A2(new_n509), .A3(new_n683), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n437), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  INV_X1    g519(.A(new_n658), .ZN(new_n706));
  INV_X1    g520(.A(new_n547), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n595), .A2(new_n587), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n569), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n578), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n707), .A2(new_n607), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n701), .A2(new_n510), .A3(new_n706), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  NAND2_X1  g527(.A1(new_n621), .A2(new_n623), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT99), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n621), .A2(new_n614), .A3(new_n623), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n436), .A3(new_n716), .A4(new_n651), .ZN(new_n717));
  INV_X1    g531(.A(new_n191), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n692), .A2(new_n718), .A3(new_n514), .A4(new_n385), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n638), .A2(new_n710), .A3(new_n607), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n345), .ZN(G27));
  OAI21_X1  g536(.A(new_n548), .B1(new_n580), .B2(new_n582), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n585), .A2(new_n599), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(new_n707), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n725), .B1(new_n724), .B2(new_n707), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n317), .A2(G469), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n191), .B1(new_n514), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n610), .A2(new_n611), .A3(new_n323), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n728), .A2(new_n732), .A3(new_n717), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n601), .A2(new_n730), .A3(new_n731), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n717), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n734), .C1(new_n735), .C2(new_n717), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n733), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n247), .ZN(G33));
  INV_X1    g555(.A(new_n652), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n743));
  INV_X1    g557(.A(new_n732), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(KEYINPUT107), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n743), .A2(new_n601), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  NOR2_X1   g561(.A1(new_n624), .A2(new_n625), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n437), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT43), .Z(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n608), .A3(new_n638), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT44), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n307), .A2(new_n310), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(G469), .ZN(new_n755));
  NAND2_X1  g569(.A1(G469), .A2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n514), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n718), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(new_n662), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n731), .B(KEYINPUT108), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n718), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n659), .A2(new_n322), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n702), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n547), .A3(new_n681), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  INV_X1    g587(.A(G952), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n750), .A2(new_n648), .A3(new_n711), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n774), .B(G953), .C1(new_n775), .C2(new_n701), .ZN(new_n776));
  INV_X1    g590(.A(new_n677), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n693), .A2(new_n191), .A3(new_n770), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n707), .A3(new_n504), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n626), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n726), .A2(new_n727), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n648), .A2(new_n750), .A3(new_n782), .A4(new_n778), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT48), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n776), .B(new_n781), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT115), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n322), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n775), .A2(new_n661), .A3(new_n694), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n779), .A2(new_n436), .A3(new_n748), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n767), .B(new_n768), .C1(new_n192), .C2(new_n693), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n750), .A2(new_n648), .A3(new_n711), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n762), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n720), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n750), .A2(new_n648), .A3(new_n800), .A4(new_n778), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n792), .A2(new_n793), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n794), .A2(new_n799), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(KEYINPUT51), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n788), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n788), .B(KEYINPUT116), .C1(new_n804), .C2(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n658), .A2(new_n612), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n730), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n638), .A2(new_n650), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n677), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n681), .A2(new_n701), .A3(new_n800), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n687), .A2(new_n742), .A3(new_n688), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n689), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n721), .A2(new_n656), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT113), .A3(new_n689), .A4(new_n815), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n820), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n437), .B1(new_n653), .B2(new_n654), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n731), .A2(new_n500), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n687), .A2(KEYINPUT112), .A3(new_n651), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT112), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n515), .A2(new_n192), .A3(new_n638), .A4(new_n651), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n702), .A2(new_n500), .A3(new_n437), .A4(new_n731), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n744), .A2(new_n681), .A3(new_n800), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n746), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n740), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n641), .A2(new_n631), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n641), .B2(new_n631), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n626), .A2(new_n613), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n626), .A2(KEYINPUT110), .A3(new_n613), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n609), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n847), .A2(new_n602), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n695), .A2(new_n704), .A3(new_n712), .A4(new_n698), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n838), .A2(new_n842), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(new_n841), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n641), .A2(new_n631), .A3(new_n839), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n848), .A2(new_n853), .A3(new_n854), .A4(new_n849), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n740), .A2(new_n837), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n818), .A2(new_n823), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n852), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n811), .B1(new_n851), .B2(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n826), .A2(new_n852), .A3(new_n850), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n857), .B2(new_n860), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n865), .B2(new_n811), .ZN(new_n866));
  OAI22_X1  g680(.A1(new_n810), .A2(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n749), .A2(new_n547), .A3(new_n682), .A4(new_n323), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n869), .A2(KEYINPUT109), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(KEYINPUT109), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n693), .B(KEYINPUT49), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n677), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n870), .A2(new_n661), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n874), .ZN(G75));
  NOR2_X1   g689(.A1(new_n851), .A2(new_n861), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(G210), .A3(G902), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n371), .A2(new_n377), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(new_n375), .Z(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT55), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT56), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n883), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n877), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n774), .A2(G953), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT118), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n884), .A2(new_n887), .A3(new_n890), .ZN(G51));
  OAI211_X1 g705(.A(new_n857), .B(new_n852), .C1(new_n824), .C2(new_n825), .ZN(new_n892));
  INV_X1    g706(.A(new_n860), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n893), .B2(new_n850), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT54), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n897), .B(new_n811), .C1(new_n851), .C2(new_n861), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n756), .B(KEYINPUT57), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n304), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n900), .B2(new_n304), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n876), .A2(G902), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(new_n755), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n890), .B1(new_n904), .B2(new_n906), .ZN(G54));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n426), .B1(new_n909), .B2(G475), .ZN(new_n910));
  INV_X1    g724(.A(G475), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n905), .A2(new_n908), .A3(new_n911), .A4(new_n427), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n889), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(KEYINPUT121), .B(new_n889), .C1(new_n910), .C2(new_n912), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n617), .A2(new_n619), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT122), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n896), .A2(new_n898), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n889), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n922), .B2(new_n889), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n866), .B2(new_n919), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G63));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  AND2_X1   g743(.A1(new_n876), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n636), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n889), .C1(new_n536), .C2(new_n930), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT61), .B1(new_n931), .B2(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G66));
  OAI21_X1  g748(.A(G953), .B1(new_n506), .B2(new_n350), .ZN(new_n935));
  INV_X1    g749(.A(new_n855), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n881), .B1(G898), .B2(new_n441), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NOR2_X1   g753(.A1(new_n557), .A2(new_n558), .ZN(new_n940));
  XNOR2_X1  g754(.A(KEYINPUT125), .B(KEYINPUT126), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(new_n422), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n764), .A2(new_n772), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n780), .B1(new_n500), .B2(new_n436), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(new_n601), .A3(new_n663), .A4(new_n731), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n821), .A2(new_n689), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n679), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT62), .Z(new_n950));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n944), .B1(new_n951), .B2(new_n441), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n945), .A2(new_n746), .ZN(new_n953));
  INV_X1    g767(.A(new_n740), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n782), .A2(new_n812), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n954), .B(new_n948), .C1(new_n761), .C2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n441), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n649), .A2(G953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n952), .B1(new_n959), .B2(new_n944), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n289), .B2(new_n649), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n951), .B2(new_n855), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n587), .B1(new_n559), .B2(new_n560), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n890), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n586), .A2(new_n564), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n953), .A2(new_n855), .A3(new_n956), .ZN(new_n969));
  INV_X1    g783(.A(new_n964), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n865), .A2(new_n968), .A3(new_n966), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n972), .B1(new_n964), .B2(new_n973), .ZN(G57));
endmodule


