//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n551, new_n552, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n591, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n459), .B1(new_n448), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(new_n464), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n462), .A2(new_n473), .A3(G137), .A4(new_n464), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n464), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n472), .A2(new_n474), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n462), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  INV_X1    g056(.A(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n470), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI211_X1 g074(.A(KEYINPUT70), .B(new_n498), .C1(new_n499), .C2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT5), .B1(new_n499), .B2(KEYINPUT70), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND2_X1  g091(.A1(new_n505), .A2(KEYINPUT72), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n518), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n512), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n510), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(G89), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n521), .A2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(new_n520), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  INV_X1    g109(.A(new_n512), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n526), .A2(G90), .B1(G52), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n539), .B(new_n540), .C1(new_n531), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n541), .B1(new_n517), .B2(new_n519), .ZN(new_n543));
  INV_X1    g118(.A(new_n540), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT73), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n545), .A3(G651), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n526), .A2(G81), .B1(G43), .B2(new_n535), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n512), .B2(new_n554), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n512), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(new_n556), .B1(new_n526), .B2(G91), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n507), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G299));
  OAI21_X1  g135(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n526), .A2(G87), .B1(G49), .B2(new_n535), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT74), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(G288));
  AOI22_X1  g142(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n568), .A2(new_n507), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n510), .A2(new_n570), .B1(new_n512), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n569), .A2(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n507), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n526), .A2(G85), .B1(G47), .B2(new_n535), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G301), .A2(G868), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(G92), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n505), .A2(G66), .ZN(new_n582));
  INV_X1    g157(.A(G79), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n499), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n578), .B1(new_n587), .B2(G868), .ZN(G284));
  OAI21_X1  g163(.A(new_n578), .B1(new_n587), .B2(G868), .ZN(G321));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G286), .A2(new_n590), .ZN(new_n591));
  XOR2_X1   g166(.A(G299), .B(KEYINPUT75), .Z(new_n592));
  AOI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n590), .ZN(G280));
  XNOR2_X1  g168(.A(G280), .B(KEYINPUT76), .ZN(G297));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n587), .B1(new_n595), .B2(G860), .ZN(G148));
  NAND2_X1  g171(.A1(new_n587), .A2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT77), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n480), .A2(G123), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n482), .A2(G135), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n464), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT79), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2096), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n462), .A2(new_n475), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G156));
  XNOR2_X1  g189(.A(KEYINPUT15), .B(G2435), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT82), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2427), .B(G2430), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(KEYINPUT14), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT81), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2451), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n621), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G14), .C1(new_n630), .C2(new_n628), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(G401));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  XNOR2_X1  g211(.A(G2067), .B(G2678), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT17), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n638), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(G227));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1961), .B(G1966), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT20), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n657), .C1(new_n648), .C2(new_n656), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G229));
  AND2_X1   g241(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n667));
  NOR2_X1   g242(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(G6), .A2(G16), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n569), .A2(new_n572), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(G16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT32), .ZN(new_n673));
  INV_X1    g248(.A(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  MUX2_X1   g250(.A(G23), .B(new_n563), .S(G16), .Z(new_n676));
  XOR2_X1   g251(.A(KEYINPUT33), .B(G1976), .Z(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR2_X1   g254(.A1(G16), .A2(G22), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G166), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT87), .B(G1971), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND4_X1  g258(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(KEYINPUT34), .ZN(new_n686));
  MUX2_X1   g261(.A(G24), .B(G290), .S(G16), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT86), .B(G1986), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G25), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n480), .A2(G119), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n482), .A2(G131), .ZN(new_n693));
  OR2_X1    g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n694), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n685), .A2(new_n686), .A3(new_n689), .A4(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n667), .B(new_n669), .S(new_n701), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n690), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n480), .A2(G128), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n482), .A2(G140), .ZN(new_n706));
  OR2_X1    g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n707), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(new_n690), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT89), .B(G2067), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n587), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G4), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(G1348), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n548), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G16), .B2(G19), .ZN(new_n721));
  INV_X1    g296(.A(G1341), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n690), .B1(KEYINPUT24), .B2(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(KEYINPUT24), .B2(G34), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n477), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n690), .A2(G32), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT26), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n475), .A2(G105), .ZN(new_n736));
  INV_X1    g311(.A(G141), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n470), .B2(new_n737), .ZN(new_n738));
  AOI211_X1 g313(.A(new_n735), .B(new_n738), .C1(G129), .C2(new_n480), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n733), .B1(new_n739), .B2(new_n690), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT93), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n732), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n714), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n714), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n744), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT95), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n725), .A2(new_n726), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n690), .A2(G33), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT25), .Z(new_n753));
  INV_X1    g328(.A(G139), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n754), .B2(new_n470), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT91), .Z(new_n756));
  AOI22_X1  g331(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n756), .B1(G2105), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n690), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G2072), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n743), .B2(new_n742), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n690), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n690), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT29), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n760), .A2(G2072), .B1(G2090), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT99), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT100), .B(G1956), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT94), .B(G28), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT30), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(new_n690), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n773), .B1(new_n775), .B2(new_n777), .C1(new_n607), .C2(new_n690), .ZN(new_n778));
  NOR2_X1   g353(.A1(G27), .A2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(G29), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT96), .B(G2078), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n782), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n762), .A2(new_n766), .A3(new_n772), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n730), .A2(new_n731), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT92), .Z(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n745), .B2(new_n747), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n765), .A2(G2090), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n714), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n786), .A2(new_n789), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n727), .A2(new_n749), .A3(new_n750), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n702), .A2(new_n799), .ZN(G311));
  INV_X1    g375(.A(G311), .ZN(G150));
  NOR2_X1   g376(.A1(new_n586), .A2(new_n595), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT38), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT102), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n526), .A2(G93), .B1(G55), .B2(new_n535), .ZN(new_n805));
  INV_X1    g380(.A(new_n519), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n498), .B1(new_n501), .B2(G543), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT70), .B1(new_n499), .B2(KEYINPUT71), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n518), .B1(new_n809), .B2(new_n500), .ZN(new_n810));
  OAI21_X1  g385(.A(G67), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n507), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n805), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G67), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n517), .B2(new_n519), .ZN(new_n817));
  INV_X1    g392(.A(new_n812), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n814), .B(G651), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n804), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n546), .A2(new_n547), .ZN(new_n822));
  OAI21_X1  g397(.A(G651), .B1(new_n817), .B2(new_n818), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT101), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n824), .A2(KEYINPUT102), .A3(new_n819), .A4(new_n805), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n546), .B(new_n547), .C1(new_n815), .C2(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n803), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  AOI21_X1  g405(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n821), .A2(new_n825), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT104), .Z(G145));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n480), .A2(G130), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n464), .A2(G118), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G142), .B2(new_n482), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n611), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n697), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(KEYINPUT107), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n709), .B(new_n496), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n739), .ZN(new_n849));
  INV_X1    g424(.A(new_n759), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n846), .A2(KEYINPUT107), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n849), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n759), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n849), .B(KEYINPUT105), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n850), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n847), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n477), .B(new_n486), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n607), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n858), .A2(KEYINPUT106), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n855), .ZN(new_n864));
  INV_X1    g439(.A(new_n847), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n851), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n860), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n862), .B1(new_n860), .B2(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n839), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n872), .A2(KEYINPUT40), .A3(new_n868), .A4(new_n867), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n871), .A2(new_n873), .ZN(G395));
  XOR2_X1   g449(.A(new_n828), .B(new_n597), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n586), .A2(G299), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n581), .A2(new_n559), .A3(new_n557), .A4(new_n585), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n828), .B(new_n597), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT41), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(G305), .ZN(new_n887));
  XOR2_X1   g462(.A(G303), .B(new_n563), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n885), .B(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n889), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n833), .A2(new_n590), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(G295));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n883), .A2(new_n882), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n534), .A2(G286), .A3(new_n536), .ZN(new_n901));
  AOI21_X1  g476(.A(G286), .B1(new_n534), .B2(new_n536), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n826), .A2(new_n827), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n826), .B2(new_n827), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n828), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n826), .A2(new_n903), .A3(new_n827), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n878), .A3(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n900), .B(KEYINPUT108), .C1(new_n904), .C2(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n914), .B2(new_n889), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n908), .A2(new_n890), .A3(new_n912), .A4(new_n913), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n899), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n906), .A2(new_n912), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n889), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n916), .A3(new_n899), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n917), .A2(KEYINPUT44), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n914), .A2(new_n889), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n899), .A3(new_n868), .A4(new_n916), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n916), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n923), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n915), .A2(new_n916), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n923), .A3(new_n920), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT44), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(G397));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n476), .A2(new_n466), .A3(G40), .A4(new_n468), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n496), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n496), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n940), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT49), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n671), .A2(new_n674), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n671), .A2(new_n674), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(G305), .A2(G1981), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT49), .A3(new_n949), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n952), .A2(G8), .A3(new_n946), .A4(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1976), .ZN(new_n956));
  INV_X1    g531(.A(G288), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n949), .B(KEYINPUT116), .ZN(new_n959));
  AOI211_X1 g534(.A(new_n938), .B(new_n947), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT114), .A4(G1976), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n563), .B2(new_n956), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n946), .A2(G8), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n565), .A2(new_n956), .A3(new_n566), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n955), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n964), .B2(KEYINPUT52), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(new_n969), .A3(KEYINPUT52), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n943), .A2(new_n974), .A3(new_n945), .ZN(new_n975));
  INV_X1    g550(.A(G2090), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n496), .B2(new_n941), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n939), .A2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT45), .B1(new_n496), .B2(new_n941), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n981), .A2(new_n939), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1971), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n986));
  NAND2_X1  g561(.A1(G303), .A2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND4_X1  g565(.A1(G303), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(G8), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n960), .B1(new_n973), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n975), .A2(new_n731), .A3(new_n978), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n975), .A2(KEYINPUT118), .A3(new_n978), .A4(new_n731), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n943), .B2(new_n945), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n939), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n496), .A2(new_n944), .A3(new_n941), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n944), .B1(new_n496), .B2(new_n941), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT117), .A3(new_n940), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n980), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1001), .B1(new_n795), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G168), .A2(G8), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n996), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n795), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n999), .A2(new_n1000), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(KEYINPUT119), .A3(G8), .A4(G168), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n972), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n970), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n939), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g599(.A1(new_n1024), .A2(G2090), .B1(G1971), .B2(new_n983), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n992), .B1(new_n1025), .B2(G8), .ZN(new_n1026));
  NOR4_X1   g601(.A1(new_n1020), .A2(new_n994), .A3(new_n1026), .A4(new_n968), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT63), .B1(new_n1018), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n994), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT63), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(new_n985), .B2(new_n993), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n973), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1017), .B2(new_n1013), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n995), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT120), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n946), .A2(G2067), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1348), .B1(new_n975), .B2(new_n978), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT60), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n587), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1039), .ZN(new_n1044));
  INV_X1    g619(.A(G2067), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n947), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1046), .A3(KEYINPUT60), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT123), .A3(new_n586), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1043), .A2(new_n1048), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1040), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1037), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1041), .A2(new_n1042), .A3(new_n587), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n586), .B1(new_n1047), .B2(KEYINPUT123), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT124), .A3(new_n1050), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G299), .B(KEYINPUT57), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1956), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1059));
  INV_X1    g634(.A(new_n982), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n940), .A2(new_n1060), .A3(new_n980), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT122), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1024), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1058), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n983), .A2(new_n1062), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1066), .A2(KEYINPUT61), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT58), .B(G1341), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n947), .A2(new_n1073), .B1(G1996), .B2(new_n1061), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1074), .A2(new_n548), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1074), .B2(new_n548), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n1079));
  AND4_X1   g654(.A1(new_n1079), .A2(new_n1071), .A3(new_n1065), .A4(KEYINPUT61), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1072), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1052), .A2(new_n1057), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1065), .B1(new_n1083), .B2(new_n586), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1071), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n975), .A2(new_n978), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n745), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1061), .B2(G2078), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1004), .A2(new_n980), .A3(new_n1009), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(G301), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n981), .A2(new_n982), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n476), .A2(KEYINPUT125), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n476), .A2(KEYINPUT125), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(G40), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1098), .A2(new_n465), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1089), .A2(new_n1091), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1087), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1092), .A2(G301), .A3(new_n1094), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1087), .B1(new_n1102), .B2(G171), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1027), .B(new_n1104), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1014), .A2(new_n1015), .A3(G168), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1111), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1016), .A2(G286), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(G8), .A3(new_n1111), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1115), .B2(KEYINPUT51), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1086), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n938), .B1(new_n1011), .B2(G168), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1112), .B1(new_n1121), .B2(new_n1114), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT62), .B1(new_n1122), .B2(new_n1113), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1027), .A2(new_n1095), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT120), .B(new_n995), .C1(new_n1028), .C2(new_n1033), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1036), .A2(new_n1118), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1060), .A2(KEYINPUT110), .A3(new_n939), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT110), .B1(new_n1060), .B2(new_n939), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n739), .B(G1996), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n709), .B(new_n1045), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n696), .B(new_n699), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G290), .A2(G1986), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1137), .B(new_n1139), .C1(KEYINPUT111), .C2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1140), .A2(KEYINPUT111), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1130), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1127), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1996), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1130), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT46), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1130), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1132), .A2(new_n739), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT47), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1151), .A2(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(KEYINPUT127), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1148), .A2(new_n1139), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1154), .A2(KEYINPUT48), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1154), .A2(KEYINPUT48), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n697), .A2(new_n699), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1133), .A2(new_n1157), .B1(G2067), .B2(new_n709), .ZN(new_n1158));
  AOI22_X1  g733(.A1(new_n1155), .A2(new_n1156), .B1(new_n1130), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1152), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1144), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g736(.A1(G227), .A2(new_n460), .ZN(new_n1163));
  AND3_X1   g737(.A1(new_n665), .A2(new_n633), .A3(new_n1163), .ZN(new_n1164));
  OAI221_X1 g738(.A(new_n1164), .B1(new_n917), .B2(new_n921), .C1(new_n869), .C2(new_n870), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


