//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT67), .A3(G101), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n464), .A2(new_n466), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G124), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n486), .A2(new_n489), .A3(new_n467), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OR3_X1    g071(.A1(new_n496), .A2(G100), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(G100), .B2(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n467), .A2(G112), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(new_n498), .A3(G2104), .A4(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n492), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  NAND4_X1  g077(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n467), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n487), .A2(G138), .A3(new_n467), .A4(new_n505), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G114), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G2105), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n511), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n512));
  AND2_X1   g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n464), .A2(new_n466), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT6), .B(G651), .Z(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G166));
  NAND2_X1  g105(.A1(new_n523), .A2(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(new_n522), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n528), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G89), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n528), .A2(KEYINPUT72), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT6), .B(G651), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(G543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G51), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n541), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND2_X1  g125(.A1(new_n535), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n525), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n539), .A2(G90), .ZN(new_n554));
  INV_X1    g129(.A(G52), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n546), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(G171));
  AND2_X1   g132(.A1(new_n535), .A2(G56), .ZN(new_n558));
  AND2_X1   g133(.A1(G68), .A2(G543), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n547), .A2(G43), .B1(G81), .B2(new_n539), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G188));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n546), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n546), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n525), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G91), .B2(new_n539), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n574), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G166), .ZN(G303));
  OAI21_X1  g155(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n542), .A2(G49), .A3(G543), .A4(new_n545), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n539), .A2(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(KEYINPUT74), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n581), .A2(new_n586), .A3(new_n582), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n585), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n532), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT75), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n594), .A3(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(G48), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n532), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n543), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n593), .A2(new_n595), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n535), .A2(G60), .ZN(new_n601));
  NAND2_X1  g176(.A1(G72), .A2(G543), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n525), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n539), .A2(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n546), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n539), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  INV_X1    g186(.A(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n546), .A2(new_n612), .B1(new_n525), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT76), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n609), .B1(new_n619), .B2(G868), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n494), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n467), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(G123), .B2(new_n491), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT81), .Z(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n487), .A2(new_n473), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(G2100), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n643), .B1(KEYINPUT80), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(KEYINPUT80), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n638), .B(new_n646), .C1(new_n647), .C2(new_n643), .ZN(G156));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2435), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n659), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n669), .ZN(new_n674));
  AND3_X1   g249(.A1(new_n674), .A2(KEYINPUT17), .A3(new_n671), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n674), .B2(KEYINPUT17), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n675), .A2(new_n676), .A3(new_n670), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n682), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n687), .B1(new_n682), .B2(new_n685), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n690), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT21), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT84), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  AND3_X1   g274(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G16), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G16), .B2(G23), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT33), .B(G1976), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(G6), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G305), .B2(G16), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  OAI211_X1 g284(.A(new_n704), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n706), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1971), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n491), .A2(G119), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n494), .A2(G131), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n467), .A2(G107), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(KEYINPUT85), .A2(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(KEYINPUT85), .A2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  MUX2_X1   g299(.A(G25), .B(new_n721), .S(new_n724), .Z(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT35), .B(G1991), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n706), .A2(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n607), .B2(new_n706), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n716), .A2(new_n731), .B1(KEYINPUT86), .B2(new_n732), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n733), .A2(KEYINPUT86), .A3(new_n732), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(KEYINPUT86), .B2(new_n732), .ZN(new_n735));
  INV_X1    g310(.A(new_n724), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(G34), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n483), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n563), .A2(new_n706), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n706), .B2(G19), .ZN(new_n746));
  INV_X1    g321(.A(G1341), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n746), .A2(new_n747), .B1(new_n743), .B2(new_n742), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n744), .B(new_n748), .C1(new_n747), .C2(new_n746), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n706), .A2(G20), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT92), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n623), .B2(new_n706), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1956), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G33), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n494), .A2(G139), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  INV_X1    g335(.A(G127), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n485), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  INV_X1    g338(.A(G103), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n470), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n762), .A2(G2105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n756), .B1(new_n769), .B2(G29), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n770), .A2(G2072), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(KEYINPUT89), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n706), .A2(G5), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G171), .B2(new_n706), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT90), .Z(new_n776));
  AOI21_X1  g351(.A(new_n772), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n736), .A2(G26), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  OR2_X1    g354(.A1(G104), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n781));
  INV_X1    g356(.A(G128), .ZN(new_n782));
  INV_X1    g357(.A(G140), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n781), .B1(new_n490), .B2(new_n782), .C1(new_n783), .C2(new_n493), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(G29), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n776), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G1961), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n771), .A2(KEYINPUT89), .B1(new_n788), .B2(new_n787), .ZN(new_n792));
  INV_X1    g367(.A(G1348), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n619), .A2(new_n706), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G4), .B2(new_n706), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n736), .A2(G35), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n736), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT29), .Z(new_n798));
  INV_X1    g373(.A(G2090), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n793), .A2(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n777), .A2(new_n791), .A3(new_n792), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n804));
  OR2_X1    g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NAND2_X1  g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G1966), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G21), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G168), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n807), .B1(new_n808), .B2(new_n811), .C1(new_n637), .C2(new_n736), .ZN(new_n812));
  NOR2_X1   g387(.A1(G164), .A2(new_n736), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G27), .B2(new_n736), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT91), .B(G2078), .Z(new_n815));
  AOI22_X1  g390(.A1(new_n811), .A2(new_n808), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n770), .A2(G2072), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT26), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n822), .A2(new_n823), .B1(G105), .B2(new_n473), .ZN(new_n824));
  INV_X1    g399(.A(G129), .ZN(new_n825));
  INV_X1    g400(.A(G141), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n824), .B1(new_n490), .B2(new_n825), .C1(new_n826), .C2(new_n493), .ZN(new_n827));
  MUX2_X1   g402(.A(G32), .B(new_n827), .S(G29), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT27), .B(G1996), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n818), .A2(new_n819), .A3(new_n830), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n795), .A2(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n755), .A2(new_n801), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n734), .A2(new_n735), .A3(new_n833), .ZN(G150));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n835));
  XNOR2_X1  g410(.A(G150), .B(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n539), .A2(G93), .ZN(new_n837));
  INV_X1    g412(.A(G55), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n546), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n535), .A2(G67), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n839), .B1(new_n842), .B2(G651), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n562), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n562), .A2(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n619), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n853));
  AOI21_X1  g428(.A(G860), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  INV_X1    g430(.A(new_n845), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT37), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(G145));
  XNOR2_X1  g434(.A(new_n786), .B(new_n827), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n512), .A2(new_n861), .A3(new_n514), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n512), .B2(new_n514), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n509), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n768), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT98), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n865), .A2(KEYINPUT97), .A3(new_n768), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n515), .A2(KEYINPUT96), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n512), .A2(new_n861), .A3(new_n514), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n870), .A2(new_n871), .B1(new_n507), .B2(new_n508), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n860), .B(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n869), .B1(new_n873), .B2(new_n769), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n501), .B(new_n641), .Z(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n867), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n867), .B2(new_n875), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n494), .A2(G142), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT99), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n491), .A2(G130), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n467), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n721), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n637), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n483), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n879), .A2(new_n880), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(new_n875), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n866), .B(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n876), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n878), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n890), .A2(new_n891), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT40), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n890), .A2(new_n900), .A3(new_n897), .A4(new_n891), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(G395));
  XNOR2_X1  g477(.A(new_n623), .B(new_n618), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT41), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n848), .B(new_n628), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n607), .B(G303), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n700), .B(G305), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(KEYINPUT100), .B(KEYINPUT42), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT101), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n913), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n908), .A2(KEYINPUT101), .A3(new_n913), .ZN(new_n917));
  OAI21_X1  g492(.A(G868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g494(.A(new_n918), .B1(G868), .B2(new_n845), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  XNOR2_X1  g496(.A(G286), .B(G171), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n848), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n903), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n904), .A2(new_n923), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n911), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT102), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n911), .B1(new_n925), .B2(new_n926), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n928), .B2(new_n931), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n921), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n931), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT44), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(new_n477), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n487), .B2(G125), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n480), .B1(new_n941), .B2(new_n467), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(G40), .A3(new_n482), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT104), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n481), .A2(new_n946), .A3(G40), .A4(new_n482), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(KEYINPUT103), .B(G1384), .Z(new_n949));
  AOI21_X1  g524(.A(KEYINPUT45), .B1(new_n864), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n786), .B(new_n788), .ZN(new_n953));
  INV_X1    g528(.A(G1996), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n827), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n721), .B(new_n726), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(G290), .A2(G1986), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n959), .A2(KEYINPUT105), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1976), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT52), .B1(G288), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n948), .A2(new_n967), .A3(new_n864), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n700), .A2(G1976), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G8), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT110), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n968), .A2(G8), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(new_n965), .A3(new_n969), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n593), .A2(new_n978), .A3(new_n595), .A4(new_n599), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  INV_X1    g555(.A(new_n599), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n592), .B1(new_n981), .B2(KEYINPUT112), .ZN(new_n983));
  OAI21_X1  g558(.A(G1981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(KEYINPUT113), .A2(KEYINPUT49), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n980), .B(new_n984), .C1(KEYINPUT113), .C2(KEYINPUT49), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n974), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n973), .A2(new_n977), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n517), .A2(new_n967), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n948), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT106), .B(G1971), .Z(new_n996));
  AND2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n864), .A2(new_n998), .A3(new_n967), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT107), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n864), .A2(new_n1001), .A3(new_n998), .A4(new_n967), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n799), .A4(new_n948), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n999), .A2(KEYINPUT107), .B1(KEYINPUT50), .B2(new_n991), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(new_n799), .A3(new_n948), .A4(new_n1002), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n997), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1010), .B2(KEYINPUT109), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1012), .B(new_n997), .C1(new_n1009), .C2(new_n1006), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT55), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n990), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT50), .B1(new_n872), .B2(G1384), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n948), .B(new_n1019), .C1(KEYINPUT50), .C2(new_n991), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(G2090), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1021), .B2(new_n997), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1016), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n948), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT119), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT119), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1007), .A2(new_n1027), .A3(new_n948), .A4(new_n1002), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n995), .A2(G2078), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1029), .A2(new_n773), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n517), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT114), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n992), .B1(new_n872), .B2(G1384), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n517), .A2(new_n1036), .A3(KEYINPUT45), .A4(new_n967), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n945), .A2(new_n947), .ZN(new_n1039));
  OR4_X1    g614(.A1(new_n1031), .A2(new_n1038), .A3(new_n1039), .A4(G2078), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G171), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n808), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1046), .B(new_n808), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1004), .A2(new_n743), .A3(new_n948), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT51), .B1(new_n1049), .B2(G8), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1007), .A2(new_n948), .A3(new_n1002), .ZN(new_n1051));
  AOI22_X1  g626(.A1(KEYINPUT115), .A2(new_n1044), .B1(new_n1051), .B2(new_n743), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT124), .B1(new_n1052), .B2(new_n1047), .ZN(new_n1053));
  AND4_X1   g628(.A1(KEYINPUT124), .A2(new_n1045), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1054));
  OAI21_X1  g629(.A(G168), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1050), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1049), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1045), .A2(KEYINPUT124), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1061), .B1(new_n1065), .B2(new_n1058), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1043), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1050), .ZN(new_n1068));
  AOI21_X1  g643(.A(G286), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1058), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1058), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1060), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(KEYINPUT62), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1042), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G299), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n574), .A2(KEYINPUT57), .A3(new_n577), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT117), .B(G1956), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n1020), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n993), .A2(new_n994), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT56), .B(G2072), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT118), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1083), .A2(new_n948), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1080), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1082), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n618), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1029), .A2(new_n793), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n968), .A2(G2067), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1348), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1091), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n619), .A3(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1090), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1092), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1103), .B(KEYINPUT123), .Z(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT120), .B(G1996), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n948), .A2(new_n993), .A3(new_n994), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  AOI22_X1  g684(.A1(new_n1107), .A2(new_n1108), .B1(new_n968), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1083), .A2(KEYINPUT121), .A3(new_n948), .A4(new_n1106), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n562), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1102), .A2(KEYINPUT59), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n968), .A2(new_n1109), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1111), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n563), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1113), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1104), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1080), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1082), .A2(new_n1080), .A3(new_n1086), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1114), .A2(new_n1120), .A3(new_n1122), .A4(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1094), .B1(new_n1101), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(G171), .B(KEYINPUT54), .Z(new_n1130));
  NOR2_X1   g705(.A1(new_n943), .A2(KEYINPUT125), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n943), .A2(KEYINPUT125), .ZN(new_n1132));
  INV_X1    g707(.A(G40), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1031), .A2(new_n1133), .A3(G2078), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n479), .A3(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n950), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1130), .B1(new_n994), .B2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1041), .A2(new_n1130), .B1(new_n1032), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1076), .A2(new_n1129), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1024), .B1(new_n1075), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1049), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1141));
  INV_X1    g716(.A(new_n997), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1012), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1142), .B(KEYINPUT109), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(G8), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1141), .B1(new_n1148), .B2(new_n1016), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT116), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1018), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1016), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1146), .A2(G8), .A3(new_n1017), .A4(new_n1147), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n977), .A2(new_n989), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n976), .B1(new_n975), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1141), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1152), .A2(new_n1153), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT116), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1049), .A2(G8), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(G286), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1153), .A2(new_n1157), .A3(new_n1023), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1151), .A2(new_n1160), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1153), .A2(new_n990), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n989), .A2(new_n964), .A3(new_n585), .A4(new_n587), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n980), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n974), .B2(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n963), .B1(new_n1140), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n726), .B(new_n721), .C1(new_n956), .C2(new_n952), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n786), .A2(G2067), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1173), .A2(KEYINPUT126), .A3(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT126), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(new_n952), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(new_n953), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n952), .B1(new_n1178), .B2(new_n827), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n952), .A2(KEYINPUT46), .A3(new_n954), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT46), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1181), .B1(new_n951), .B2(G1996), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n952), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT48), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n958), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1177), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT127), .B1(new_n1172), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT127), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1188), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1042), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1071), .A2(KEYINPUT62), .A3(new_n1073), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT62), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1076), .A2(new_n1129), .A3(new_n1138), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1192), .B1(new_n1198), .B2(new_n1024), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1190), .B(new_n1191), .C1(new_n1199), .C2(new_n963), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1189), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g776(.A1(new_n937), .A2(new_n932), .ZN(new_n1203));
  NOR4_X1   g777(.A1(G229), .A2(new_n461), .A3(G401), .A4(G227), .ZN(new_n1204));
  AND3_X1   g778(.A1(new_n1203), .A2(new_n1204), .A3(new_n898), .ZN(G308));
  NAND3_X1  g779(.A1(new_n1203), .A2(new_n1204), .A3(new_n898), .ZN(G225));
endmodule


