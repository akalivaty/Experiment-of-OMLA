//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT64), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G169), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n249));
  INV_X1    g0049(.A(G223), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G226), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n252), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G87), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n249), .A3(G274), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n249), .A2(G232), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n247), .B1(new_n260), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n259), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT16), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G20), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G159), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT76), .ZN(new_n277));
  XNOR2_X1  g0077(.A(G58), .B(G68), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(G20), .ZN(new_n279));
  AND2_X1   g0079(.A1(G58), .A2(G68), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(G20), .C1(new_n280), .C2(new_n201), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n276), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G20), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n255), .A2(new_n256), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n274), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n219), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT7), .B1(new_n288), .B2(new_n210), .ZN(new_n294));
  NOR4_X1   g0094(.A1(new_n255), .A2(new_n256), .A3(new_n285), .A4(G20), .ZN(new_n295));
  OAI21_X1  g0095(.A(G68), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(G20), .B1(new_n280), .B2(new_n201), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT76), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n281), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n276), .A4(new_n299), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n291), .A2(new_n293), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT77), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT65), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n292), .A2(KEYINPUT65), .A3(new_n219), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G58), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n310), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT8), .B(G58), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT8), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G58), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(KEYINPUT8), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT66), .ZN(new_n318));
  OR3_X1    g0118(.A1(new_n310), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n209), .A2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n307), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n302), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n314), .A2(new_n302), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n273), .B1(new_n301), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n291), .A2(new_n300), .A3(new_n293), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n314), .A2(new_n302), .A3(new_n322), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n323), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n272), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT18), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G190), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n260), .A2(new_n268), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n259), .B2(new_n267), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n329), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT17), .A4(new_n339), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n328), .A2(new_n334), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n332), .A2(new_n333), .ZN(new_n347));
  AOI211_X1 g0147(.A(KEYINPUT18), .B(new_n272), .C1(new_n329), .C2(new_n331), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n342), .A2(new_n343), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT78), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n275), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n318), .A2(new_n319), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n210), .A2(G33), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n304), .A2(new_n308), .ZN(new_n356));
  NOR3_X1   g0156(.A1(new_n305), .A2(new_n210), .A3(G1), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n355), .A2(new_n356), .B1(new_n202), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n320), .A2(G50), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT67), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(new_n309), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(KEYINPUT9), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT70), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n249), .A2(new_n265), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n264), .B1(new_n253), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n286), .A2(G222), .A3(new_n251), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n288), .A2(G77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n286), .A2(G1698), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n250), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G190), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(new_n337), .B2(new_n371), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT9), .B1(new_n358), .B2(new_n361), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n363), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n371), .A2(new_n270), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT68), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n358), .A2(new_n361), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(G169), .C2(new_n371), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n346), .A2(new_n351), .A3(new_n380), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G238), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n264), .B1(new_n387), .B2(new_n364), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n253), .A2(new_n251), .ZN(new_n389));
  INV_X1    g0189(.A(G232), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n391), .C1(new_n255), .C2(new_n256), .ZN(new_n392));
  AND3_X1   g0192(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n249), .B1(new_n396), .B2(KEYINPUT72), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT72), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n388), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT13), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT13), .B(new_n388), .C1(new_n397), .C2(new_n399), .ZN(new_n403));
  OAI21_X1  g0203(.A(G169), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT14), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(G169), .C1(new_n402), .C2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n397), .A2(new_n399), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(KEYINPUT13), .C1(new_n409), .C2(new_n388), .ZN(new_n410));
  INV_X1    g0210(.A(new_n403), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT73), .B1(new_n400), .B2(new_n401), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(G179), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n275), .A2(G50), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n210), .A2(G33), .A3(G77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n284), .A2(G20), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n356), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT74), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT11), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  INV_X1    g0222(.A(new_n308), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT65), .B1(new_n292), .B2(new_n219), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n418), .B(new_n422), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n420), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n425), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(new_n356), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT11), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n307), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT12), .B1(new_n307), .B2(G68), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n357), .A2(new_n293), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n284), .B1(new_n209), .B2(G20), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n430), .A2(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n426), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT75), .A4(new_n434), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n414), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(G190), .ZN(new_n442));
  OAI21_X1  g0242(.A(G200), .B1(new_n402), .B2(new_n403), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n316), .A2(new_n317), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n275), .B1(G20), .B2(G77), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n354), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(new_n293), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n432), .A2(G77), .A3(new_n320), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(G77), .B2(new_n307), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n286), .A2(G232), .A3(new_n251), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n288), .A2(G107), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n368), .C2(new_n387), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n370), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT69), .ZN(new_n457));
  INV_X1    g0257(.A(new_n264), .ZN(new_n458));
  INV_X1    g0258(.A(new_n364), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(G244), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n456), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n452), .B1(new_n463), .B2(G200), .ZN(new_n464));
  OAI21_X1  g0264(.A(G190), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n270), .B1(new_n461), .B2(new_n462), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n467), .A2(new_n452), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n247), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n441), .A2(new_n444), .A3(new_n466), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n386), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT6), .A2(G107), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT79), .A2(KEYINPUT6), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n207), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI22_X1  g0279(.A1(new_n478), .A2(new_n479), .B1(KEYINPUT79), .B2(KEYINPUT6), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(G20), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n275), .A2(G77), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT80), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G107), .B1(new_n294), .B2(new_n295), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT80), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n293), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n307), .A2(G97), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n309), .B1(new_n209), .B2(G33), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G97), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT81), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT81), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n487), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n251), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n286), .A2(G250), .A3(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n370), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT5), .B(G41), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n262), .A2(G1), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(G274), .A3(new_n249), .A4(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(G1), .A2(G13), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(new_n504), .B1(new_n507), .B2(new_n248), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(G257), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT82), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(G190), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(G200), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n492), .A2(new_n494), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n513), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT82), .B1(new_n502), .B2(new_n509), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n247), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n502), .A2(new_n509), .A3(new_n270), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n491), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n249), .A2(G274), .A3(new_n504), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n209), .A2(G45), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n249), .A2(G250), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT83), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT83), .ZN(new_n528));
  OAI211_X1 g0328(.A(G244), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n529));
  OAI211_X1 g0329(.A(G238), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n527), .A2(new_n528), .B1(new_n370), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(G169), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n527), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n370), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n535), .A2(new_n270), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n447), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n489), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n286), .A2(new_n210), .A3(G68), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n354), .B2(new_n205), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n207), .A2(G87), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT19), .B1(new_n393), .B2(new_n394), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n210), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n293), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n447), .A2(new_n357), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n540), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n528), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT83), .B1(new_n522), .B2(new_n524), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n536), .B(G190), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT84), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n535), .A2(new_n555), .A3(G190), .A4(new_n536), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n337), .B1(new_n535), .B2(new_n536), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n423), .A2(new_n424), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n209), .A2(G33), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n559), .A2(G87), .A3(new_n560), .A4(new_n307), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n548), .A2(new_n549), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n538), .A2(new_n550), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n516), .A2(new_n521), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT91), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n210), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT22), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT88), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n286), .A2(new_n210), .A3(new_n569), .A4(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  INV_X1    g0374(.A(G116), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n354), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(KEYINPUT89), .B1(new_n210), .B2(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT23), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT23), .ZN(new_n579));
  OAI211_X1 g0379(.A(KEYINPUT89), .B(new_n579), .C1(new_n210), .C2(G107), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n573), .A2(new_n574), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n574), .B1(new_n573), .B2(new_n581), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n293), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n357), .A2(new_n206), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n585), .B(KEYINPUT25), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n489), .B2(G107), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n589));
  OAI211_X1 g0389(.A(G250), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n370), .B1(new_n508), .B2(G264), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(new_n335), .A3(new_n505), .ZN(new_n594));
  AOI21_X1  g0394(.A(G200), .B1(new_n593), .B2(new_n505), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n566), .B1(new_n588), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n505), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n337), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n593), .A2(new_n335), .A3(new_n505), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n601), .A2(KEYINPUT91), .A3(new_n584), .A4(new_n587), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n286), .A2(G257), .A3(new_n251), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n288), .A2(G303), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n370), .ZN(new_n608));
  AND2_X1   g0408(.A1(KEYINPUT5), .A2(G41), .ZN(new_n609));
  NOR2_X1   g0409(.A1(KEYINPUT5), .A2(G41), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n504), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(G270), .A3(new_n249), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n612), .A2(KEYINPUT85), .A3(new_n505), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT85), .B1(new_n612), .B2(new_n505), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n608), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n575), .A2(G20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n293), .A2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(G20), .B1(G33), .B2(G283), .ZN(new_n619));
  INV_X1    g0419(.A(G33), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G97), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n621), .A3(KEYINPUT86), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT86), .B1(new_n619), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n618), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT20), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT20), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n618), .C1(new_n623), .C2(new_n624), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n616), .A2(G1), .A3(new_n305), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n575), .B1(new_n209), .B2(G33), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n432), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n615), .A2(new_n632), .A3(G169), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n612), .A2(new_n505), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT85), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n612), .A2(new_n505), .A3(KEYINPUT85), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n370), .B2(new_n607), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(G179), .A3(new_n632), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n615), .A2(new_n632), .A3(KEYINPUT21), .A4(G169), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n635), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n608), .B(G190), .C1(new_n613), .C2(new_n614), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n639), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n337), .B1(new_n647), .B2(new_n608), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT87), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n615), .A2(G200), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT87), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n644), .A4(new_n645), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n598), .A2(KEYINPUT90), .A3(G169), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n593), .A2(G179), .A3(new_n505), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT90), .B1(new_n598), .B2(G169), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n588), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n603), .A2(new_n643), .A3(new_n653), .A4(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n473), .A2(new_n565), .A3(new_n659), .ZN(G372));
  AND3_X1   g0460(.A1(new_n469), .A2(new_n452), .A3(new_n467), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n440), .B2(new_n414), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n350), .A2(new_n444), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n349), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n380), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(new_n385), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n516), .A2(new_n521), .A3(new_n564), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n643), .A2(new_n658), .B1(new_n597), .B2(new_n602), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT26), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n557), .A2(new_n563), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n535), .A2(new_n536), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n247), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n533), .A2(new_n270), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n550), .A3(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n671), .A2(new_n519), .A3(new_n520), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n494), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n493), .B1(new_n487), .B2(new_n490), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n670), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n519), .A2(new_n520), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n564), .A3(KEYINPUT26), .A4(new_n491), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n669), .A2(new_n683), .A3(new_n675), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n666), .B1(new_n473), .B2(new_n685), .ZN(G369));
  AND2_X1   g0486(.A1(new_n643), .A2(new_n653), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n306), .A2(new_n688), .A3(new_n210), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G213), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n306), .A2(new_n210), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(KEYINPUT93), .B(G343), .Z(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n632), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n643), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n603), .A2(new_n658), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n588), .A2(new_n697), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n695), .A2(new_n696), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n658), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n643), .A2(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n658), .A2(new_n697), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n213), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n217), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(new_n491), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n670), .B1(new_n676), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n492), .A2(new_n494), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n681), .A2(new_n564), .A3(new_n724), .A4(KEYINPUT26), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n642), .A2(new_n641), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n658), .A2(new_n728), .A3(new_n635), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n603), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n675), .B1(new_n730), .B2(new_n565), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT29), .B(new_n706), .C1(new_n727), .C2(new_n731), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n667), .A2(new_n668), .B1(new_n550), .B2(new_n538), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n697), .B1(new_n733), .B2(new_n683), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n732), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(G330), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n512), .A2(new_n513), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n640), .A2(G179), .A3(new_n533), .A4(new_n593), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n608), .B(G179), .C1(new_n613), .C2(new_n614), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n535), .A2(new_n536), .A3(new_n593), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(KEYINPUT30), .A3(new_n512), .A4(new_n513), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n510), .A2(new_n598), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n640), .A2(G179), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n533), .A2(KEYINPUT94), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n533), .A2(KEYINPUT94), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n740), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n750), .B2(new_n697), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n667), .A2(new_n703), .A3(new_n687), .A4(new_n706), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n736), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n735), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n721), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR2_X1   g0559(.A1(new_n305), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n209), .B1(new_n760), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n716), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n715), .A2(new_n288), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT95), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(G355), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT95), .B1(new_n207), .B2(G87), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n766), .A2(new_n767), .B1(G116), .B2(new_n213), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n245), .A2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n715), .A2(new_n286), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n262), .B2(new_n218), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n219), .B1(G20), .B2(new_n247), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n210), .B1(new_n782), .B2(G190), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G97), .ZN(new_n785));
  NAND3_X1  g0585(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(new_n335), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n785), .B1(new_n788), .B2(new_n284), .C1(new_n202), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT97), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n210), .B2(G190), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n337), .A2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n335), .A2(KEYINPUT97), .A3(G20), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G107), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n794), .A2(G20), .A3(G190), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G87), .ZN(new_n801));
  NAND2_X1  g0601(.A1(G20), .A2(G179), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n802), .A2(new_n335), .A3(G200), .ZN(new_n803));
  NOR3_X1   g0603(.A1(new_n802), .A2(G190), .A3(G200), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G58), .A2(new_n803), .B1(new_n804), .B2(G77), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n798), .A2(new_n801), .A3(new_n286), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT32), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n793), .A2(new_n782), .A3(new_n795), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(new_n809), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n808), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n812));
  OR4_X1    g0612(.A1(new_n791), .A2(new_n806), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n804), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  INV_X1    g0615(.A(G303), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n814), .A2(new_n815), .B1(new_n799), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n286), .B(new_n817), .C1(G322), .C2(new_n803), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n809), .A2(G329), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n796), .ZN(new_n821));
  INV_X1    g0621(.A(G317), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n822), .A2(KEYINPUT33), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(KEYINPUT33), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n787), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n789), .A2(G326), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n783), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n813), .B1(new_n821), .B2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT98), .Z(new_n830));
  INV_X1    g0630(.A(new_n779), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n763), .B1(new_n774), .B2(new_n781), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT99), .ZN(new_n833));
  INV_X1    g0633(.A(new_n778), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n700), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n702), .A2(new_n763), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(G330), .B2(new_n700), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  INV_X1    g0639(.A(KEYINPUT100), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n452), .A2(new_n840), .A3(new_n697), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n449), .A2(new_n451), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT100), .B1(new_n842), .B2(new_n706), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n465), .B2(new_n464), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n470), .A3(new_n706), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n733), .B2(new_n683), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n468), .A2(new_n469), .A3(new_n706), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n845), .B2(new_n661), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n848), .B1(new_n734), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n763), .B1(new_n852), .B2(new_n756), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n756), .B2(new_n852), .ZN(new_n854));
  INV_X1    g0654(.A(new_n803), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n855), .A2(new_n827), .B1(new_n799), .B2(new_n206), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n286), .B(new_n856), .C1(G116), .C2(new_n804), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n797), .A2(G87), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n857), .B(new_n858), .C1(new_n815), .C2(new_n808), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n785), .B1(new_n788), .B2(new_n820), .C1(new_n816), .C2(new_n790), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G143), .A2(new_n803), .B1(new_n804), .B2(G159), .ZN(new_n861));
  INV_X1    g0661(.A(G150), .ZN(new_n862));
  INV_X1    g0662(.A(G137), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n861), .B1(new_n788), .B2(new_n862), .C1(new_n863), .C2(new_n790), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT34), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n797), .A2(G68), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n286), .B1(new_n783), .B2(new_n310), .C1(new_n799), .C2(new_n202), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G132), .B2(new_n809), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n864), .A2(new_n865), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n859), .A2(new_n860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n779), .ZN(new_n873));
  INV_X1    g0673(.A(new_n763), .ZN(new_n874));
  INV_X1    g0674(.A(G77), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n779), .A2(new_n776), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n873), .B(new_n877), .C1(new_n851), .C2(new_n777), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n854), .A2(new_n878), .ZN(G384));
  NOR2_X1   g0679(.A1(new_n760), .A2(new_n209), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n440), .A2(new_n697), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n441), .A2(new_n444), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n439), .A2(new_n442), .A3(new_n443), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n440), .B(new_n697), .C1(new_n883), .C2(new_n414), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n750), .A2(new_n697), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT31), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n659), .A2(new_n565), .A3(new_n697), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n885), .B(new_n851), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n329), .A2(new_n331), .A3(new_n339), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n332), .ZN(new_n897));
  INV_X1    g0697(.A(new_n695), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n301), .B2(new_n326), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AND4_X1   g0700(.A1(new_n895), .A2(new_n327), .A3(new_n899), .A4(new_n340), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n349), .B2(new_n350), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n894), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT103), .ZN(new_n905));
  INV_X1    g0705(.A(new_n899), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n344), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n327), .A2(new_n899), .A3(new_n340), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n327), .A2(new_n899), .A3(new_n895), .A4(new_n340), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n893), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT103), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n291), .A2(new_n356), .A3(new_n300), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n898), .B1(new_n914), .B2(new_n326), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n273), .B1(new_n914), .B2(new_n326), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n915), .A3(new_n340), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n344), .A2(new_n916), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n912), .A2(new_n913), .B1(KEYINPUT38), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n892), .B1(new_n905), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n344), .A2(new_n916), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n910), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n924), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n922), .A2(new_n923), .B1(new_n892), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n753), .A2(new_n754), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n472), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n736), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n930), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n732), .B(new_n472), .C1(new_n734), .C2(KEYINPUT29), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n666), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT39), .B1(new_n921), .B2(new_n905), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n926), .A2(new_n927), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n414), .A2(new_n440), .A3(new_n706), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT101), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n849), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n885), .B1(new_n847), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n926), .A2(new_n927), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n945), .A2(new_n946), .B1(new_n349), .B2(new_n898), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n937), .B(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n880), .B1(new_n934), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n934), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n477), .A2(new_n480), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT35), .ZN(new_n953));
  OAI211_X1 g0753(.A(G116), .B(new_n220), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT36), .Z(new_n956));
  NOR3_X1   g0756(.A1(new_n217), .A2(new_n875), .A3(new_n280), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n284), .A2(G50), .ZN(new_n958));
  OAI211_X1 g0758(.A(G1), .B(new_n305), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(G367));
  OAI221_X1 g0760(.A(new_n780), .B1(new_n213), .B2(new_n447), .C1(new_n771), .C2(new_n237), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n799), .A2(new_n575), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n962), .A2(KEYINPUT46), .B1(new_n815), .B2(new_n790), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT46), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n288), .B1(new_n814), .B2(new_n820), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G303), .B2(new_n803), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n784), .A2(G107), .B1(G294), .B2(new_n787), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G97), .A2(new_n797), .B1(new_n809), .B2(G317), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n783), .A2(new_n284), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n855), .A2(new_n862), .B1(new_n799), .B2(new_n310), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(G143), .C2(new_n789), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G50), .A2(new_n804), .B1(new_n787), .B2(G159), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT112), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n974), .C1(new_n863), .C2(new_n808), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n797), .A2(G77), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n286), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT113), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n969), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  OAI211_X1 g0780(.A(new_n763), .B(new_n961), .C1(new_n980), .C2(new_n831), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n697), .A2(new_n562), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n564), .A2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n984), .A2(KEYINPUT106), .B1(new_n675), .B2(new_n983), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n984), .A2(KEYINPUT106), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n982), .B1(new_n834), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n516), .A2(new_n521), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n724), .A2(new_n697), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n681), .B2(new_n991), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n713), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n996));
  XOR2_X1   g0796(.A(new_n995), .B(new_n996), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n713), .A2(new_n994), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT45), .Z(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n709), .A3(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n995), .B(new_n996), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n998), .B(KEYINPUT45), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n702), .B(new_n708), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(KEYINPUT110), .B(new_n711), .C1(new_n708), .C2(new_n710), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT110), .B2(new_n711), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(new_n702), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n758), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n716), .B(KEYINPUT41), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT111), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1008), .A2(new_n1013), .A3(new_n1010), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n762), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n993), .A2(new_n711), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n521), .B1(new_n993), .B2(new_n658), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n706), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT107), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(KEYINPUT107), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT43), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1021), .A2(new_n1022), .A3(new_n1028), .A4(new_n987), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n709), .A2(new_n993), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(KEYINPUT108), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1030), .B1(new_n709), .B2(new_n993), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT108), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1027), .A2(new_n1035), .A3(new_n1031), .A4(new_n1029), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n989), .B1(new_n1015), .B2(new_n1037), .ZN(G387));
  AOI21_X1  g0838(.A(new_n286), .B1(new_n809), .B2(G326), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n799), .A2(new_n827), .B1(new_n783), .B2(new_n820), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G303), .A2(new_n804), .B1(new_n803), .B2(G317), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n789), .A2(G322), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n815), .C2(new_n788), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT48), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1040), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1039), .B1(new_n575), .B2(new_n796), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT115), .B1(new_n790), .B2(new_n811), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n862), .B2(new_n808), .C1(new_n353), .C2(new_n788), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n855), .A2(new_n202), .B1(new_n814), .B2(new_n284), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n783), .A2(new_n447), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n286), .B1(new_n799), .B2(new_n875), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n789), .A2(G159), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1055), .B1(KEYINPUT115), .B2(new_n1056), .C1(new_n205), .C2(new_n796), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1048), .A2(new_n1049), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n779), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n718), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n764), .A2(new_n1060), .B1(new_n206), .B2(new_n715), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n234), .A2(new_n262), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n445), .A2(new_n202), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n718), .B(new_n262), .C1(new_n284), .C2(new_n875), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n770), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n874), .B1(new_n1067), .B2(new_n780), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1059), .B(new_n1068), .C1(new_n708), .C2(new_n834), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1006), .B(new_n701), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1070), .A2(new_n758), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1007), .A2(new_n757), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n716), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1069), .B1(new_n761), .B2(new_n1007), .C1(new_n1075), .C2(new_n1076), .ZN(G393));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1004), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1073), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n716), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1004), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n993), .A2(new_n778), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n242), .A2(new_n770), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n780), .B1(new_n205), .B2(new_n213), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n763), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n288), .B1(new_n814), .B2(new_n827), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n788), .A2(new_n816), .B1(new_n783), .B2(new_n575), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G283), .C2(new_n800), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G311), .A2(new_n803), .B1(new_n789), .B2(G317), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  NAND2_X1  g0890(.A1(new_n809), .A2(G322), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1088), .A2(new_n1090), .A3(new_n798), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n783), .A2(new_n875), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n286), .B1(new_n799), .B2(new_n284), .C1(new_n814), .C2(new_n312), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G50), .C2(new_n787), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n809), .A2(G143), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n858), .A3(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G159), .A2(new_n803), .B1(new_n789), .B2(G150), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1085), .B1(new_n1100), .B2(new_n779), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1081), .A2(new_n762), .B1(new_n1082), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1080), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1080), .A2(new_n1102), .A3(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n776), .B1(new_n938), .B2(new_n940), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n353), .A2(new_n876), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n814), .A2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n288), .B(new_n1111), .C1(G132), .C2(new_n803), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n799), .A2(new_n862), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT53), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1113), .A2(new_n1114), .B1(new_n787), .B2(G137), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G50), .A2(new_n797), .B1(new_n809), .B2(G125), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n784), .A2(G159), .B1(G128), .B2(new_n789), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1114), .B2(new_n1113), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G97), .A2(new_n804), .B1(new_n803), .B2(G116), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n801), .A2(new_n1120), .A3(new_n288), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n867), .C1(new_n827), .C2(new_n808), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1093), .B1(G107), .B2(new_n787), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n820), .B2(new_n790), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1117), .A2(new_n1119), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n874), .B(new_n1109), .C1(new_n1125), .C2(new_n779), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1108), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(G330), .B(new_n851), .C1(new_n890), .C2(new_n891), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n882), .A2(new_n884), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n913), .B(new_n894), .C1(new_n902), .C2(new_n903), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n920), .A2(KEYINPUT38), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n912), .A2(new_n913), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n939), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n940), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1135), .A2(new_n1136), .B1(new_n945), .B2(new_n941), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n941), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n851), .B(new_n706), .C1(new_n727), .C2(new_n731), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n944), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1129), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1130), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n846), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n944), .B1(new_n684), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n941), .B1(new_n1145), .B2(new_n1129), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n938), .B2(new_n940), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n921), .A2(new_n905), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n697), .B1(new_n733), .B2(new_n726), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n944), .B1(new_n1149), .B2(new_n851), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1148), .B(new_n941), .C1(new_n1150), .C2(new_n1129), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n755), .A2(new_n851), .A3(new_n885), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1147), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1143), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1127), .B1(new_n1154), .B2(new_n761), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n755), .A2(new_n472), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n935), .A2(new_n666), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1152), .A2(new_n1150), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1145), .B1(new_n1152), .B2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n717), .B1(new_n1154), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n935), .A2(new_n666), .A3(new_n1157), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1145), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n885), .B1(new_n755), .B2(new_n851), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1130), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1150), .A2(new_n1152), .A3(new_n1159), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1143), .A2(new_n1169), .A3(new_n1153), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT118), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1137), .A2(new_n1142), .A3(new_n1130), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1152), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1162), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AND4_X1   g0974(.A1(KEYINPUT118), .A2(new_n1174), .A3(new_n716), .A4(new_n1170), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1156), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1174), .A2(new_n716), .A3(new_n1170), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT118), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1163), .A2(KEYINPUT118), .A3(new_n1170), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(KEYINPUT119), .A3(new_n1156), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1178), .A2(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(new_n948), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n384), .A2(new_n898), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n380), .A2(new_n385), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1187), .B1(new_n380), .B2(new_n385), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n892), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n923), .B1(new_n1148), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n928), .A2(new_n892), .ZN(new_n1196));
  OAI211_X1 g0996(.A(G330), .B(new_n1193), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1193), .B1(new_n929), .B2(G330), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1186), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1193), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1129), .A2(new_n850), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n931), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1196), .B1(new_n1203), .B2(KEYINPUT40), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(new_n736), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n948), .A3(new_n1197), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1200), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n776), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n288), .A2(new_n261), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n800), .A2(G77), .B1(new_n539), .B2(new_n804), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(G107), .B2(new_n803), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n797), .A2(G58), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n970), .B1(G97), .B2(new_n787), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n575), .B2(new_n790), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G283), .C2(new_n809), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1210), .B1(new_n1217), .B2(KEYINPUT58), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT120), .Z(new_n1219));
  AOI211_X1 g1019(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n811), .B2(new_n796), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n799), .A2(new_n1110), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G128), .B2(new_n803), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n804), .A2(G137), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n789), .A2(G125), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n784), .A2(G150), .B1(G132), .B2(new_n787), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1221), .B1(new_n1227), .B2(KEYINPUT59), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1217), .A2(KEYINPUT58), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n831), .B1(new_n1219), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT121), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n874), .B(new_n1232), .C1(new_n202), .C2(new_n876), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1207), .A2(new_n762), .B1(new_n1208), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1170), .A2(new_n1158), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1205), .A2(new_n948), .A3(new_n1197), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n948), .B1(new_n1205), .B2(new_n1197), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(KEYINPUT57), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n716), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1235), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1234), .B1(new_n1239), .B2(new_n1240), .ZN(G375));
  OAI21_X1  g1041(.A(new_n762), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n874), .B1(new_n284), .B2(new_n876), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT122), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n976), .A2(new_n288), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT123), .Z(new_n1246));
  AOI21_X1  g1046(.A(new_n1053), .B1(G294), .B2(new_n789), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n575), .B2(new_n788), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n800), .A2(G97), .B1(G107), .B2(new_n804), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n820), .B2(new_n855), .C1(new_n816), .C2(new_n808), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1246), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(KEYINPUT124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n789), .A2(G132), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n783), .B2(new_n202), .C1(new_n788), .C2(new_n1110), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n800), .A2(G159), .B1(G150), .B2(new_n804), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n809), .A2(G128), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n288), .B1(G137), .B2(new_n803), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1255), .A2(new_n1213), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1252), .B1(new_n1254), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(KEYINPUT124), .B2(new_n1251), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1244), .B1(new_n831), .B2(new_n1260), .C1(new_n885), .C2(new_n777), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1242), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1167), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1162), .A2(new_n1010), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1156), .A2(new_n1179), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  OR3_X1    g1070(.A1(new_n1270), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n1233), .A2(new_n1208), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n761), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1200), .A2(new_n1206), .B1(new_n1158), .B2(new_n1170), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n717), .B1(new_n1275), .B2(KEYINPUT57), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1207), .A2(new_n1235), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT57), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1276), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n696), .A2(G213), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT125), .Z(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1269), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1263), .B1(new_n1169), .B2(new_n1286), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1167), .A2(KEYINPUT60), .A3(new_n1164), .A4(new_n1168), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n716), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1262), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n854), .A3(new_n878), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(G384), .A3(new_n1262), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G375), .B1(new_n1178), .B2(new_n1184), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1275), .A2(new_n1010), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1268), .B1(new_n1234), .B2(new_n1296), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1285), .B(new_n1294), .C1(new_n1295), .C2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1282), .A2(G2897), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(KEYINPUT126), .A3(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT126), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1301), .B1(new_n1293), .B2(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1297), .B1(G378), .B2(new_n1280), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(new_n1282), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT119), .B1(new_n1183), .B2(new_n1156), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1177), .B(new_n1155), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1280), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1297), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1315), .A3(new_n1285), .A4(new_n1294), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1299), .A2(new_n1300), .A3(new_n1309), .A4(new_n1316), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(G393), .B(new_n838), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(G387), .A2(new_n1266), .ZN(new_n1320));
  AOI211_X1 g1120(.A(KEYINPUT111), .B(new_n1009), .C1(new_n1079), .C2(new_n758), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1013), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n761), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1036), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G390), .B1(new_n1325), .B2(new_n989), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1319), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(G387), .A2(new_n1266), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1325), .A2(new_n989), .A3(G390), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n1329), .A3(new_n1318), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1327), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1317), .A2(new_n1331), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1328), .A2(new_n1329), .A3(new_n1318), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1318), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1314), .A2(new_n1285), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1336), .B2(new_n1307), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1298), .A2(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1314), .A2(KEYINPUT63), .A3(new_n1285), .A4(new_n1294), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1335), .A2(new_n1337), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1332), .A2(new_n1341), .ZN(G405));
  OAI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1327), .A2(new_n1344), .A3(new_n1330), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1280), .A2(new_n1268), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1295), .A2(new_n1346), .A3(new_n1294), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1294), .B1(new_n1295), .B2(new_n1346), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1343), .A2(new_n1345), .A3(new_n1348), .A4(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1349), .ZN(new_n1351));
  OAI211_X1 g1151(.A(new_n1331), .B(KEYINPUT127), .C1(new_n1347), .C2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(G402));
endmodule


