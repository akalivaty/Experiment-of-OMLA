//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n464), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT67), .B1(new_n466), .B2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(new_n468), .A3(KEYINPUT3), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n479), .A2(new_n481), .A3(new_n472), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n483), .A2(G137), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n479), .A2(new_n481), .A3(new_n472), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n489), .B2(new_n485), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n468), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G101), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n478), .A2(new_n491), .A3(new_n493), .ZN(G160));
  NOR2_X1   g069(.A1(new_n489), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G136), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n463), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n482), .A2(KEYINPUT69), .A3(new_n464), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n489), .B2(new_n463), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(G124), .B2(new_n503), .ZN(G162));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  AND3_X1   g081(.A1(new_n483), .A2(G138), .A3(new_n484), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n473), .B1(new_n471), .B2(new_n472), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n483), .A2(G138), .A3(new_n484), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT4), .B1(new_n489), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(G126), .A2(G2105), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n479), .A2(new_n481), .A3(new_n472), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G114), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G2105), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n517), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n505), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  AOI211_X1 g096(.A(KEYINPUT70), .B(new_n519), .C1(new_n510), .C2(new_n512), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(G164));
  OR2_X1    g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  OR2_X1    g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G88), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n529), .A2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g117(.A(new_n533), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n526), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n535), .A2(G89), .ZN(new_n547));
  NAND2_X1  g122(.A1(G63), .A2(G651), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G168));
  NAND2_X1  g125(.A1(new_n526), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n528), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n524), .A2(new_n525), .B1(new_n531), .B2(new_n532), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G90), .B1(new_n533), .B2(G52), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n555), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  AOI22_X1  g135(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n528), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n533), .A2(G43), .ZN(new_n563));
  INV_X1    g138(.A(G81), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n536), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n536), .A2(KEYINPUT72), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT72), .B1(new_n536), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n546), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n573), .A2(new_n574), .B1(G651), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n533), .A2(G53), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  OAI21_X1  g157(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n533), .A2(G49), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n536), .ZN(G288));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n524), .B2(new_n525), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT73), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT73), .B(G651), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n556), .A2(G86), .B1(new_n533), .B2(G48), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n528), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n533), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n536), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  OR3_X1    g178(.A1(G171), .A2(KEYINPUT74), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT74), .B1(G171), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n556), .A2(G92), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT10), .Z(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n546), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n612), .ZN(G284));
  OAI211_X1 g188(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n612), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT75), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n612), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g200(.A1(new_n508), .A2(new_n509), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n492), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n503), .A2(G123), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT76), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n495), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n463), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n631), .A2(new_n638), .A3(new_n639), .ZN(G156));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  INV_X1    g238(.A(new_n656), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1971), .B(G1976), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  AOI211_X1 g252(.A(new_n675), .B(new_n677), .C1(new_n670), .C2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT78), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G24), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n601), .B2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n686), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(G6), .A2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G305), .B2(new_n686), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n686), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n686), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT82), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n696), .A2(new_n697), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n694), .A2(new_n698), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n690), .B1(new_n706), .B2(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n495), .A2(G131), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT79), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n503), .A2(G119), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n463), .C2(G107), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT80), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n709), .B1(new_n715), .B2(G29), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT81), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n707), .B(new_n719), .C1(KEYINPUT34), .C2(new_n706), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n708), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n503), .A2(G128), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G116), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n464), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n495), .B2(G140), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n730), .A2(new_n731), .A3(G29), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n731), .B1(new_n730), .B2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n723), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2067), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n708), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n708), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT88), .Z(new_n739));
  INV_X1    g314(.A(G2078), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n708), .A2(G33), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT25), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G139), .B2(new_n495), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n463), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2072), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT84), .ZN(new_n753));
  NAND2_X1  g328(.A1(G160), .A2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT24), .B2(new_n755), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(G2084), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n495), .A2(G141), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT26), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n762), .A2(new_n763), .B1(G105), .B2(new_n492), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G129), .B2(new_n503), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n708), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n708), .B2(G32), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT85), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n750), .A2(new_n751), .ZN(new_n772));
  AND4_X1   g347(.A1(new_n753), .A2(new_n758), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT86), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT86), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G35), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G162), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT29), .B(G2090), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI21_X1  g355(.A(G2084), .B1(new_n754), .B2(new_n757), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G4), .A2(G16), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n612), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G16), .A2(G19), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n566), .B2(G16), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G1341), .Z(new_n789));
  NOR2_X1   g364(.A1(G168), .A2(new_n686), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n686), .B2(G21), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G28), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT30), .ZN(new_n795));
  AOI21_X1  g370(.A(G29), .B1(new_n794), .B2(KEYINPUT30), .ZN(new_n796));
  OR2_X1    g371(.A1(KEYINPUT31), .A2(G11), .ZN(new_n797));
  NAND2_X1  g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n789), .A2(new_n793), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n791), .A2(new_n792), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT87), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n786), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n686), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n686), .ZN(new_n805));
  INV_X1    g380(.A(G1961), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n708), .B2(new_n637), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT89), .B(KEYINPUT23), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n686), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G299), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1956), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n770), .B2(new_n768), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n803), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n775), .A2(new_n782), .A3(new_n815), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n721), .A2(new_n743), .A3(new_n774), .A4(new_n816), .ZN(G311));
  XNOR2_X1  g392(.A(G311), .B(KEYINPUT90), .ZN(G150));
  AOI22_X1  g393(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(new_n528), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n556), .A2(G93), .B1(new_n533), .B2(G55), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n566), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n822), .A2(new_n566), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  INV_X1    g408(.A(new_n612), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n620), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT92), .Z(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n828), .B1(new_n839), .B2(new_n841), .ZN(G145));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n749), .A2(KEYINPUT95), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n766), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n519), .B1(new_n510), .B2(new_n512), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n729), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G118), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n464), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n851), .A2(new_n850), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n852), .A2(new_n853), .B1(new_n495), .B2(G142), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n503), .A2(new_n855), .A3(G130), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n503), .B2(G130), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT98), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n629), .ZN(new_n860));
  INV_X1    g435(.A(new_n715), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n848), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(new_n715), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT99), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n848), .A3(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G162), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n637), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n843), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n843), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n869), .ZN(new_n877));
  AOI21_X1  g452(.A(G37), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  AOI21_X1  g453(.A(KEYINPUT40), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n878), .B(KEYINPUT40), .C1(new_n880), .C2(new_n873), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n879), .A2(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(new_n832), .B(new_n622), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n834), .A2(new_n617), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n612), .A2(G299), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n834), .A2(KEYINPUT101), .A3(new_n617), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n891), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n889), .B1(new_n899), .B2(new_n884), .ZN(new_n900));
  XNOR2_X1  g475(.A(G288), .B(KEYINPUT103), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G303), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n905));
  XOR2_X1   g480(.A(new_n904), .B(new_n905), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n900), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G868), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n824), .A2(new_n603), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G331));
  XOR2_X1   g485(.A(G331), .B(KEYINPUT105), .Z(G295));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n912));
  OAI21_X1  g487(.A(G301), .B1(new_n912), .B2(G168), .ZN(new_n913));
  NAND2_X1  g488(.A1(G168), .A2(new_n912), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n832), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n832), .A2(new_n915), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(new_n887), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n896), .A2(new_n918), .A3(new_n897), .A4(new_n898), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n904), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n921), .A2(G37), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n904), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(KEYINPUT41), .B(new_n893), .C1(new_n916), .C2(new_n917), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n904), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n888), .B2(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n921), .A2(G37), .A3(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n929), .A2(KEYINPUT108), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n929), .B2(KEYINPUT108), .ZN(new_n931));
  OAI221_X1 g506(.A(KEYINPUT44), .B1(KEYINPUT43), .B2(new_n924), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n922), .B2(new_n923), .ZN(new_n934));
  NOR4_X1   g509(.A1(new_n921), .A2(new_n928), .A3(KEYINPUT43), .A4(G37), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT107), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT107), .B(new_n937), .C1(new_n934), .C2(new_n935), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n938), .B2(new_n940), .ZN(G397));
  INV_X1    g516(.A(KEYINPUT127), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n506), .B1(new_n482), .B2(new_n507), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n483), .A2(new_n506), .A3(G138), .A4(new_n484), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n944), .B1(new_n470), .B2(new_n474), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n520), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT109), .ZN(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n513), .B2(new_n520), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n478), .A2(G40), .A3(new_n491), .A4(new_n493), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n715), .B(new_n718), .Z(new_n958));
  XNOR2_X1  g533(.A(new_n729), .B(G2067), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n766), .B(G1996), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n601), .B(G1986), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT120), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n946), .A2(new_n966), .A3(new_n947), .ZN(new_n967));
  NAND3_X1  g542(.A1(G160), .A2(new_n967), .A3(G40), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n947), .B1(new_n521), .B2(new_n522), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(KEYINPUT50), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G2084), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n955), .B1(new_n953), .B2(new_n948), .ZN(new_n972));
  OAI211_X1 g547(.A(KEYINPUT45), .B(new_n947), .C1(new_n521), .C2(new_n522), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n970), .A2(new_n971), .B1(new_n792), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G8), .ZN(new_n976));
  NOR2_X1   g551(.A1(G168), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n965), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n792), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n846), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n955), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n946), .A2(KEYINPUT70), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n846), .A2(new_n505), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n985), .B2(new_n966), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(G2084), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT120), .A3(new_n977), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n979), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(KEYINPUT51), .B(new_n978), .C1(new_n975), .C2(new_n976), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(G8), .C1(new_n987), .C2(G286), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  INV_X1    g570(.A(G2090), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n982), .B(new_n996), .C1(new_n985), .C2(new_n966), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n969), .A2(new_n953), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n846), .A2(new_n953), .A3(G1384), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n955), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1971), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT110), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n693), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n997), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G303), .A2(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1009));
  NOR2_X1   g584(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT112), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1003), .A2(G8), .A3(new_n1007), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n700), .A2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT115), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  INV_X1    g600(.A(new_n493), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n476), .B1(new_n626), .B2(new_n465), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n464), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n950), .A2(new_n1028), .A3(G40), .A4(new_n491), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1029), .B2(G8), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1025), .B(G8), .C1(new_n955), .C2(new_n948), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1021), .B(new_n1024), .C1(new_n1030), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT49), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G305), .A2(G1981), .ZN(new_n1035));
  INV_X1    g610(.A(G1981), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n592), .A2(new_n1036), .A3(new_n594), .A4(new_n593), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(KEYINPUT49), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n1030), .A2(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1033), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n955), .A2(new_n948), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT114), .B1(new_n1044), .B2(new_n976), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1031), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1043), .B1(new_n1046), .B2(new_n1021), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n955), .B1(KEYINPUT50), .B2(new_n948), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n966), .B(new_n947), .C1(new_n521), .C2(new_n522), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(G2090), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1052), .B2(new_n1002), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1020), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1001), .B(new_n740), .C1(new_n985), .C2(KEYINPUT45), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n986), .A2(new_n806), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT53), .A4(new_n740), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G171), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1056), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n994), .A2(new_n995), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1045), .A2(new_n1031), .B1(G1976), .B2(new_n700), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1033), .B(new_n1041), .C1(new_n1067), .C2(new_n1043), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n975), .A2(new_n976), .A3(G286), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT63), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1055), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1071), .B2(new_n1020), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1054), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1007), .A2(G8), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1003), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT63), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1041), .A2(new_n1022), .A3(new_n700), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1079), .A2(new_n1037), .B1(new_n1031), .B2(new_n1045), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1073), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1051), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT116), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1051), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT57), .B1(new_n578), .B2(KEYINPUT117), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(G299), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n999), .A2(new_n1001), .A3(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(KEYINPUT118), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1086), .B1(new_n1051), .B2(new_n1083), .ZN(new_n1094));
  AOI211_X1 g669(.A(KEYINPUT116), .B(G1956), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1090), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1090), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n1103), .B2(new_n982), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1029), .A2(G2067), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n612), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1001), .B(new_n1111), .C1(new_n985), .C2(KEYINPUT45), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1113), .B1(new_n1029), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n999), .A2(KEYINPUT119), .A3(new_n1111), .A4(new_n1001), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1117), .B2(new_n566), .ZN(new_n1118));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n829), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1104), .A2(new_n1120), .A3(new_n1105), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n612), .B2(new_n1122), .ZN(new_n1123));
  NOR4_X1   g698(.A1(new_n1104), .A2(new_n1120), .A3(new_n834), .A4(new_n1105), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1118), .A2(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1096), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1109), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n976), .B1(new_n975), .B2(G168), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n979), .A2(new_n988), .B1(new_n1133), .B2(new_n991), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1056), .B1(new_n1134), .B2(new_n990), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT124), .B1(new_n1062), .B2(G171), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n740), .A2(KEYINPUT53), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1000), .A2(new_n955), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n986), .A2(new_n806), .B1(new_n954), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1059), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1141), .B2(G171), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(G301), .A4(new_n1059), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1136), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1140), .A2(G301), .A3(new_n1059), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1140), .A2(new_n1149), .A3(new_n1059), .A4(G301), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(new_n1063), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n1137), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1151), .B2(new_n1137), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1135), .B(new_n1146), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1082), .B1(new_n1132), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1066), .B1(new_n1156), .B2(KEYINPUT125), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1073), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1068), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n993), .A2(new_n1146), .A3(new_n1020), .A4(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1154), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1151), .A2(new_n1152), .A3(new_n1137), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI221_X1 g738(.A(new_n1126), .B1(new_n1118), .B2(new_n1119), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1108), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1158), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n964), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n956), .A2(new_n1111), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT46), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n959), .A2(new_n766), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n957), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n861), .A2(new_n718), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n961), .A2(new_n1176), .B1(G2067), .B2(new_n730), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n956), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT126), .Z(new_n1179));
  INV_X1    g754(.A(new_n962), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n957), .A2(G1986), .A3(G290), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1180), .A2(new_n956), .B1(KEYINPUT48), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(KEYINPUT48), .B2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1175), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n942), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n964), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1065), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1156), .A2(KEYINPUT125), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1184), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(KEYINPUT127), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1185), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g767(.A1(new_n876), .A2(new_n878), .ZN(new_n1194));
  NOR4_X1   g768(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1195));
  AND3_X1   g769(.A1(new_n1194), .A2(new_n936), .A3(new_n1195), .ZN(G308));
  NAND3_X1  g770(.A1(new_n1194), .A2(new_n936), .A3(new_n1195), .ZN(G225));
endmodule


