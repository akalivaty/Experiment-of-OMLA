

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788;

  XNOR2_X1 U373 ( .A(n575), .B(KEYINPUT32), .ZN(n649) );
  XNOR2_X1 U374 ( .A(n558), .B(n557), .ZN(n773) );
  XNOR2_X1 U375 ( .A(n526), .B(n362), .ZN(n571) );
  NOR2_X2 U376 ( .A1(n670), .A2(n759), .ZN(n671) );
  OR2_X2 U377 ( .A1(n787), .A2(n786), .ZN(n465) );
  NAND2_X1 U378 ( .A1(n448), .A2(n693), .ZN(n779) );
  XNOR2_X1 U379 ( .A(n402), .B(n625), .ZN(n448) );
  NAND2_X1 U380 ( .A1(n383), .A2(n450), .ZN(n382) );
  XNOR2_X1 U381 ( .A(n469), .B(KEYINPUT86), .ZN(n684) );
  XNOR2_X1 U382 ( .A(n601), .B(n492), .ZN(n605) );
  AND2_X1 U383 ( .A1(n441), .A2(n439), .ZN(n438) );
  XNOR2_X1 U384 ( .A(n475), .B(n474), .ZN(n547) );
  XNOR2_X1 U385 ( .A(G146), .B(G125), .ZN(n508) );
  XNOR2_X1 U386 ( .A(KEYINPUT3), .B(G119), .ZN(n475) );
  NAND2_X1 U387 ( .A1(n744), .A2(n447), .ZN(n445) );
  NAND2_X1 U388 ( .A1(n684), .A2(n415), .ZN(n414) );
  AND2_X1 U389 ( .A1(n413), .A2(n416), .ZN(n412) );
  AND2_X1 U390 ( .A1(n467), .A2(n418), .ZN(n415) );
  NOR2_X1 U391 ( .A1(n756), .A2(G902), .ZN(n541) );
  INV_X1 U392 ( .A(G113), .ZN(n474) );
  XNOR2_X1 U393 ( .A(n508), .B(n507), .ZN(n529) );
  INV_X1 U394 ( .A(KEYINPUT10), .ZN(n507) );
  XNOR2_X1 U395 ( .A(n552), .B(n551), .ZN(n558) );
  NAND2_X1 U396 ( .A1(n438), .A2(n445), .ZN(n601) );
  NOR2_X1 U397 ( .A1(n440), .A2(n446), .ZN(n439) );
  INV_X1 U398 ( .A(n701), .ZN(n446) );
  XOR2_X1 U399 ( .A(G137), .B(KEYINPUT69), .Z(n556) );
  XNOR2_X1 U400 ( .A(n515), .B(n514), .ZN(n552) );
  INV_X1 U401 ( .A(G134), .ZN(n514) );
  XNOR2_X1 U402 ( .A(n431), .B(KEYINPUT91), .ZN(n430) );
  XOR2_X1 U403 ( .A(G131), .B(G140), .Z(n561) );
  INV_X1 U404 ( .A(G210), .ZN(n437) );
  AND2_X1 U405 ( .A1(n636), .A2(n468), .ZN(n467) );
  INV_X1 U406 ( .A(KEYINPUT47), .ZN(n468) );
  INV_X1 U407 ( .A(KEYINPUT77), .ZN(n418) );
  OR2_X1 U408 ( .A1(n684), .A2(n420), .ZN(n413) );
  NOR2_X1 U409 ( .A1(KEYINPUT77), .A2(KEYINPUT47), .ZN(n420) );
  INV_X1 U410 ( .A(KEYINPUT15), .ZN(n485) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT101), .ZN(n486) );
  NOR2_X1 U412 ( .A1(n616), .A2(n353), .ZN(n617) );
  XNOR2_X1 U413 ( .A(n382), .B(n381), .ZN(n380) );
  INV_X1 U414 ( .A(G237), .ZN(n487) );
  OR2_X1 U415 ( .A1(n744), .A2(n442), .ZN(n441) );
  NAND2_X1 U416 ( .A1(n351), .A2(n443), .ZN(n442) );
  INV_X1 U417 ( .A(n590), .ZN(n424) );
  XNOR2_X1 U418 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n550) );
  OR2_X1 U419 ( .A1(n745), .A2(G902), .ZN(n568) );
  XNOR2_X1 U420 ( .A(n579), .B(KEYINPUT66), .ZN(n711) );
  NAND2_X1 U421 ( .A1(n354), .A2(n434), .ZN(n390) );
  NOR2_X1 U422 ( .A1(n377), .A2(n759), .ZN(n376) );
  NAND2_X1 U423 ( .A1(n700), .A2(n673), .ZN(n378) );
  NOR2_X1 U424 ( .A1(n379), .A2(G472), .ZN(n377) );
  XNOR2_X1 U425 ( .A(n461), .B(n460), .ZN(n766) );
  XNOR2_X1 U426 ( .A(G104), .B(G101), .ZN(n461) );
  XNOR2_X1 U427 ( .A(G110), .B(G107), .ZN(n460) );
  XNOR2_X1 U428 ( .A(n476), .B(n547), .ZN(n765) );
  XNOR2_X1 U429 ( .A(n529), .B(n472), .ZN(n471) );
  XNOR2_X1 U430 ( .A(n530), .B(KEYINPUT83), .ZN(n472) );
  XNOR2_X1 U431 ( .A(G128), .B(G119), .ZN(n527) );
  XOR2_X1 U432 ( .A(G140), .B(G110), .Z(n528) );
  XOR2_X1 U433 ( .A(KEYINPUT7), .B(G107), .Z(n518) );
  INV_X1 U434 ( .A(G146), .ZN(n559) );
  XNOR2_X1 U435 ( .A(n766), .B(KEYINPUT74), .ZN(n563) );
  NAND2_X1 U436 ( .A1(n449), .A2(n624), .ZN(n402) );
  INV_X1 U437 ( .A(KEYINPUT116), .ZN(n603) );
  NOR2_X1 U438 ( .A1(n602), .A2(n601), .ZN(n403) );
  AND2_X1 U439 ( .A1(n394), .A2(n406), .ZN(n393) );
  NAND2_X1 U440 ( .A1(n664), .A2(n673), .ZN(n397) );
  INV_X2 U441 ( .A(G953), .ZN(n781) );
  XNOR2_X1 U442 ( .A(n454), .B(n451), .ZN(n506) );
  INV_X1 U443 ( .A(G475), .ZN(n435) );
  NAND2_X1 U444 ( .A1(n436), .A2(n433), .ZN(n411) );
  AND2_X1 U445 ( .A1(n419), .A2(n417), .ZN(n416) );
  OR2_X1 U446 ( .A1(n467), .A2(n418), .ZN(n417) );
  NAND2_X1 U447 ( .A1(n356), .A2(KEYINPUT47), .ZN(n419) );
  INV_X1 U448 ( .A(KEYINPUT93), .ZN(n381) );
  XNOR2_X1 U449 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n477) );
  NAND2_X1 U450 ( .A1(n447), .A2(n662), .ZN(n444) );
  XNOR2_X1 U451 ( .A(n502), .B(KEYINPUT20), .ZN(n536) );
  XNOR2_X1 U452 ( .A(n429), .B(n428), .ZN(n544) );
  XNOR2_X1 U453 ( .A(KEYINPUT78), .B(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U454 ( .A(G116), .B(G101), .ZN(n428) );
  XNOR2_X1 U455 ( .A(G131), .B(G146), .ZN(n542) );
  INV_X1 U456 ( .A(n662), .ZN(n443) );
  NAND2_X1 U457 ( .A1(n760), .A2(n662), .ZN(n431) );
  INV_X1 U458 ( .A(n779), .ZN(n391) );
  INV_X1 U459 ( .A(KEYINPUT48), .ZN(n462) );
  XNOR2_X1 U460 ( .A(n465), .B(n598), .ZN(n464) );
  AND2_X1 U461 ( .A1(n352), .A2(n683), .ZN(n618) );
  XNOR2_X1 U462 ( .A(n425), .B(KEYINPUT21), .ZN(n714) );
  AND2_X1 U463 ( .A1(n536), .A2(G221), .ZN(n425) );
  XNOR2_X1 U464 ( .A(n368), .B(KEYINPUT1), .ZN(n710) );
  INV_X1 U465 ( .A(G902), .ZN(n554) );
  XNOR2_X1 U466 ( .A(n456), .B(n455), .ZN(n454) );
  XNOR2_X1 U467 ( .A(G104), .B(G122), .ZN(n456) );
  XNOR2_X1 U468 ( .A(G143), .B(G113), .ZN(n455) );
  XNOR2_X1 U469 ( .A(n453), .B(n452), .ZN(n451) );
  XNOR2_X1 U470 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n453) );
  XNOR2_X1 U471 ( .A(KEYINPUT105), .B(KEYINPUT107), .ZN(n452) );
  XOR2_X1 U472 ( .A(KEYINPUT108), .B(KEYINPUT106), .Z(n504) );
  XNOR2_X1 U473 ( .A(n484), .B(n483), .ZN(n744) );
  XNOR2_X1 U474 ( .A(n765), .B(n563), .ZN(n484) );
  NOR2_X1 U475 ( .A1(n373), .A2(n371), .ZN(n370) );
  NAND2_X1 U476 ( .A1(n372), .A2(n645), .ZN(n371) );
  NOR2_X1 U477 ( .A1(n732), .A2(n374), .ZN(n373) );
  NAND2_X1 U478 ( .A1(n458), .A2(n457), .ZN(n609) );
  AND2_X1 U479 ( .A1(n627), .A2(n585), .ZN(n610) );
  AND2_X1 U480 ( .A1(n390), .A2(n397), .ZN(n384) );
  XNOR2_X1 U481 ( .A(n534), .B(n470), .ZN(n756) );
  XNOR2_X1 U482 ( .A(n471), .B(n535), .ZN(n470) );
  XNOR2_X1 U483 ( .A(n407), .B(n520), .ZN(n751) );
  XNOR2_X1 U484 ( .A(n521), .B(n519), .ZN(n407) );
  XOR2_X1 U485 ( .A(KEYINPUT9), .B(KEYINPUT109), .Z(n516) );
  XNOR2_X1 U486 ( .A(n560), .B(n559), .ZN(n562) );
  AND2_X1 U487 ( .A1(n760), .A2(n358), .ZN(n399) );
  INV_X1 U488 ( .A(n604), .ZN(n450) );
  XNOR2_X1 U489 ( .A(n403), .B(n361), .ZN(n383) );
  XNOR2_X1 U490 ( .A(n635), .B(n634), .ZN(n688) );
  XNOR2_X1 U491 ( .A(n609), .B(KEYINPUT111), .ZN(n683) );
  NOR2_X1 U492 ( .A1(n607), .A2(n606), .ZN(n469) );
  NOR2_X1 U493 ( .A1(n629), .A2(n644), .ZN(n630) );
  XNOR2_X1 U494 ( .A(n577), .B(n576), .ZN(n366) );
  INV_X1 U495 ( .A(KEYINPUT94), .ZN(n576) );
  NAND2_X1 U496 ( .A1(n395), .A2(n393), .ZN(n577) );
  XNOR2_X1 U497 ( .A(n666), .B(n665), .ZN(n667) );
  INV_X1 U498 ( .A(KEYINPUT56), .ZN(n408) );
  XOR2_X1 U499 ( .A(n490), .B(n489), .Z(n351) );
  AND2_X1 U500 ( .A1(n355), .A2(n640), .ZN(n352) );
  OR2_X1 U501 ( .A1(n682), .A2(n615), .ZN(n353) );
  AND2_X1 U502 ( .A1(n433), .A2(n379), .ZN(n354) );
  AND2_X2 U503 ( .A1(n392), .A2(n364), .ZN(n664) );
  NOR2_X1 U504 ( .A1(n779), .A2(n400), .ZN(n696) );
  AND2_X1 U505 ( .A1(n600), .A2(n599), .ZN(n355) );
  AND2_X1 U506 ( .A1(KEYINPUT90), .A2(n705), .ZN(n356) );
  AND2_X1 U507 ( .A1(n378), .A2(n376), .ZN(n357) );
  AND2_X1 U508 ( .A1(n693), .A2(KEYINPUT2), .ZN(n358) );
  AND2_X1 U509 ( .A1(n714), .A2(n424), .ZN(n599) );
  AND2_X1 U510 ( .A1(n441), .A2(n444), .ZN(n359) );
  AND2_X1 U511 ( .A1(n397), .A2(n388), .ZN(n360) );
  INV_X1 U512 ( .A(n673), .ZN(n379) );
  XOR2_X1 U513 ( .A(n603), .B(KEYINPUT36), .Z(n361) );
  XOR2_X1 U514 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n362) );
  XOR2_X1 U515 ( .A(n744), .B(n743), .Z(n363) );
  OR2_X1 U516 ( .A1(n443), .A2(n697), .ZN(n364) );
  XNOR2_X1 U517 ( .A(KEYINPUT100), .B(KEYINPUT63), .ZN(n365) );
  AND2_X1 U518 ( .A1(n669), .A2(G953), .ZN(n759) );
  INV_X1 U519 ( .A(n759), .ZN(n398) );
  INV_X1 U520 ( .A(n644), .ZN(n375) );
  NAND2_X1 U521 ( .A1(n366), .A2(n578), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n700), .A2(n437), .ZN(n436) );
  XNOR2_X2 U523 ( .A(n401), .B(KEYINPUT79), .ZN(n700) );
  NAND2_X1 U524 ( .A1(n367), .A2(n459), .ZN(n639) );
  NAND2_X1 U525 ( .A1(n637), .A2(n636), .ZN(n367) );
  XNOR2_X1 U526 ( .A(n368), .B(KEYINPUT113), .ZN(n592) );
  NOR2_X1 U527 ( .A1(n711), .A2(n368), .ZN(n627) );
  XNOR2_X2 U528 ( .A(n568), .B(n567), .ZN(n368) );
  NAND2_X1 U529 ( .A1(n370), .A2(n369), .ZN(n647) );
  NAND2_X1 U530 ( .A1(n732), .A2(KEYINPUT34), .ZN(n369) );
  NAND2_X1 U531 ( .A1(n644), .A2(KEYINPUT34), .ZN(n372) );
  NAND2_X1 U532 ( .A1(n375), .A2(n426), .ZN(n374) );
  XNOR2_X1 U533 ( .A(n643), .B(KEYINPUT33), .ZN(n732) );
  NOR2_X1 U534 ( .A1(n700), .A2(n555), .ZN(n434) );
  INV_X1 U535 ( .A(n382), .ZN(n691) );
  NAND2_X1 U536 ( .A1(n617), .A2(n380), .ZN(n404) );
  NAND2_X1 U537 ( .A1(n357), .A2(n384), .ZN(n386) );
  NAND2_X1 U538 ( .A1(n385), .A2(n360), .ZN(n387) );
  AND2_X1 U539 ( .A1(n357), .A2(n390), .ZN(n385) );
  NAND2_X1 U540 ( .A1(n386), .A2(n365), .ZN(n389) );
  NAND2_X1 U541 ( .A1(n389), .A2(n387), .ZN(G57) );
  INV_X1 U542 ( .A(n365), .ZN(n388) );
  NAND2_X1 U543 ( .A1(n430), .A2(n391), .ZN(n392) );
  NOR2_X1 U544 ( .A1(n571), .A2(n640), .ZN(n396) );
  INV_X1 U545 ( .A(n640), .ZN(n394) );
  INV_X1 U546 ( .A(n571), .ZN(n395) );
  NAND2_X1 U547 ( .A1(n396), .A2(n574), .ZN(n575) );
  NAND2_X1 U548 ( .A1(n399), .A2(n448), .ZN(n401) );
  INV_X1 U549 ( .A(n760), .ZN(n400) );
  XNOR2_X1 U550 ( .A(n773), .B(n565), .ZN(n745) );
  NAND2_X1 U551 ( .A1(n605), .A2(n499), .ZN(n501) );
  NOR2_X2 U552 ( .A1(n711), .A2(n633), .ZN(n709) );
  XNOR2_X1 U553 ( .A(n548), .B(n549), .ZN(n553) );
  NAND2_X1 U554 ( .A1(n423), .A2(n599), .ZN(n422) );
  XNOR2_X2 U555 ( .A(G143), .B(G128), .ZN(n515) );
  XNOR2_X1 U556 ( .A(n486), .B(n485), .ZN(n663) );
  XNOR2_X1 U557 ( .A(n404), .B(KEYINPUT71), .ZN(n466) );
  NAND2_X1 U558 ( .A1(n405), .A2(n651), .ZN(n652) );
  NAND2_X1 U559 ( .A1(n650), .A2(KEYINPUT44), .ZN(n405) );
  BUF_X2 U560 ( .A(n710), .Z(n406) );
  XNOR2_X1 U561 ( .A(n409), .B(n408), .ZN(G51) );
  NAND2_X1 U562 ( .A1(n410), .A2(n398), .ZN(n409) );
  XNOR2_X1 U563 ( .A(n411), .B(n363), .ZN(n410) );
  NAND2_X1 U564 ( .A1(n414), .A2(n412), .ZN(n616) );
  XNOR2_X1 U565 ( .A(n422), .B(n421), .ZN(n593) );
  INV_X1 U566 ( .A(KEYINPUT28), .ZN(n421) );
  NOR2_X1 U567 ( .A1(n715), .A2(n591), .ZN(n423) );
  INV_X1 U568 ( .A(KEYINPUT34), .ZN(n426) );
  NAND2_X1 U569 ( .A1(n672), .A2(n554), .ZN(n427) );
  XNOR2_X1 U570 ( .A(n591), .B(KEYINPUT6), .ZN(n640) );
  XNOR2_X2 U571 ( .A(n427), .B(n555), .ZN(n591) );
  NAND2_X1 U572 ( .A1(n433), .A2(n432), .ZN(n668) );
  NOR2_X1 U573 ( .A1(n700), .A2(n435), .ZN(n432) );
  INV_X1 U574 ( .A(n664), .ZN(n433) );
  NOR2_X1 U575 ( .A1(n664), .A2(n700), .ZN(n755) );
  NAND2_X1 U576 ( .A1(n359), .A2(n445), .ZN(n586) );
  INV_X1 U577 ( .A(n444), .ZN(n440) );
  INV_X1 U578 ( .A(n351), .ZN(n447) );
  XNOR2_X1 U579 ( .A(n463), .B(n462), .ZN(n449) );
  INV_X1 U580 ( .A(n608), .ZN(n457) );
  INV_X1 U581 ( .A(n611), .ZN(n458) );
  XNOR2_X1 U582 ( .A(n459), .B(G101), .ZN(G3) );
  NAND2_X1 U583 ( .A1(n466), .A2(n464), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n542), .B(G137), .ZN(n543) );
  XNOR2_X1 U585 ( .A(n544), .B(n543), .ZN(n549) );
  XNOR2_X1 U586 ( .A(n562), .B(n561), .ZN(n564) );
  INV_X1 U587 ( .A(KEYINPUT0), .ZN(n500) );
  XNOR2_X1 U588 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n745), .B(n746), .ZN(n747) );
  XNOR2_X1 U590 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X2 U591 ( .A(G122), .B(G116), .ZN(n517) );
  XNOR2_X1 U592 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n473) );
  XNOR2_X1 U593 ( .A(n517), .B(n473), .ZN(n476) );
  XNOR2_X1 U594 ( .A(n508), .B(n477), .ZN(n480) );
  NAND2_X1 U595 ( .A1(n781), .A2(G224), .ZN(n478) );
  XNOR2_X1 U596 ( .A(n478), .B(KEYINPUT18), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n515), .B(n550), .ZN(n481) );
  XNOR2_X1 U599 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U600 ( .A(n663), .ZN(n662) );
  NAND2_X1 U601 ( .A1(n554), .A2(n487), .ZN(n491) );
  NAND2_X1 U602 ( .A1(n491), .A2(G210), .ZN(n490) );
  INV_X1 U603 ( .A(KEYINPUT87), .ZN(n488) );
  XNOR2_X1 U604 ( .A(n488), .B(KEYINPUT102), .ZN(n489) );
  NAND2_X1 U605 ( .A1(n491), .A2(G214), .ZN(n701) );
  XNOR2_X1 U606 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n492) );
  NAND2_X1 U607 ( .A1(G234), .A2(G237), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n493), .B(KEYINPUT14), .ZN(n728) );
  NOR2_X1 U609 ( .A1(G902), .A2(n781), .ZN(n495) );
  NOR2_X1 U610 ( .A1(G953), .A2(G952), .ZN(n494) );
  NOR2_X1 U611 ( .A1(n495), .A2(n494), .ZN(n496) );
  NAND2_X1 U612 ( .A1(n728), .A2(n496), .ZN(n580) );
  INV_X1 U613 ( .A(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U614 ( .A(n497), .B(G898), .ZN(n767) );
  AND2_X1 U615 ( .A1(n767), .A2(G953), .ZN(n498) );
  NOR2_X1 U616 ( .A1(n580), .A2(n498), .ZN(n499) );
  XNOR2_X2 U617 ( .A(n501), .B(n500), .ZN(n628) );
  NAND2_X1 U618 ( .A1(n663), .A2(G234), .ZN(n502) );
  NOR2_X1 U619 ( .A1(G953), .A2(G237), .ZN(n545) );
  NAND2_X1 U620 ( .A1(G214), .A2(n545), .ZN(n503) );
  XOR2_X1 U621 ( .A(n504), .B(n503), .Z(n505) );
  XNOR2_X1 U622 ( .A(n506), .B(n505), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n561), .B(n529), .ZN(n772) );
  XNOR2_X1 U624 ( .A(n509), .B(n772), .ZN(n666) );
  NAND2_X1 U625 ( .A1(n666), .A2(n554), .ZN(n511) );
  XNOR2_X1 U626 ( .A(KEYINPUT13), .B(G475), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n511), .B(n510), .ZN(n608) );
  NAND2_X1 U628 ( .A1(G234), .A2(n781), .ZN(n513) );
  XOR2_X1 U629 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n512) );
  XNOR2_X1 U630 ( .A(n513), .B(n512), .ZN(n531) );
  NAND2_X1 U631 ( .A1(G217), .A2(n531), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n552), .B(n516), .ZN(n520) );
  XNOR2_X1 U633 ( .A(n517), .B(n518), .ZN(n519) );
  NOR2_X1 U634 ( .A1(G902), .A2(n751), .ZN(n523) );
  INV_X1 U635 ( .A(G478), .ZN(n522) );
  XNOR2_X1 U636 ( .A(n523), .B(n522), .ZN(n611) );
  OR2_X1 U637 ( .A1(n457), .A2(n611), .ZN(n524) );
  INV_X1 U638 ( .A(n524), .ZN(n594) );
  AND2_X1 U639 ( .A1(n714), .A2(n594), .ZN(n525) );
  NAND2_X1 U640 ( .A1(n628), .A2(n525), .ZN(n526) );
  XNOR2_X1 U641 ( .A(n528), .B(n527), .ZN(n535) );
  INV_X1 U642 ( .A(KEYINPUT23), .ZN(n530) );
  NAND2_X1 U643 ( .A1(n531), .A2(G221), .ZN(n533) );
  XNOR2_X1 U644 ( .A(n556), .B(KEYINPUT24), .ZN(n532) );
  XOR2_X1 U645 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n538) );
  NAND2_X1 U646 ( .A1(G217), .A2(n536), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U648 ( .A(n539), .B(KEYINPUT25), .ZN(n540) );
  XNOR2_X2 U649 ( .A(n541), .B(n540), .ZN(n715) );
  NAND2_X1 U650 ( .A1(n545), .A2(G210), .ZN(n546) );
  XNOR2_X1 U651 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U652 ( .A(n550), .B(KEYINPUT70), .ZN(n551) );
  XNOR2_X1 U653 ( .A(n553), .B(n558), .ZN(n672) );
  INV_X1 U654 ( .A(G472), .ZN(n555) );
  INV_X1 U655 ( .A(n591), .ZN(n631) );
  NOR2_X1 U656 ( .A1(n578), .A2(n631), .ZN(n569) );
  INV_X1 U657 ( .A(n556), .ZN(n557) );
  NAND2_X1 U658 ( .A1(G227), .A2(n781), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U660 ( .A(G469), .B(KEYINPUT73), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT72), .ZN(n567) );
  NAND2_X1 U662 ( .A1(n569), .A2(n406), .ZN(n570) );
  OR2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n648) );
  XOR2_X1 U664 ( .A(G110), .B(KEYINPUT117), .Z(n572) );
  XNOR2_X1 U665 ( .A(n648), .B(n572), .ZN(G12) );
  INV_X1 U666 ( .A(KEYINPUT99), .ZN(n573) );
  XNOR2_X1 U667 ( .A(n406), .B(n573), .ZN(n604) );
  NOR2_X1 U668 ( .A1(n604), .A2(n578), .ZN(n574) );
  XNOR2_X1 U669 ( .A(n649), .B(G119), .ZN(G21) );
  INV_X1 U670 ( .A(n715), .ZN(n600) );
  INV_X1 U671 ( .A(n600), .ZN(n578) );
  INV_X1 U672 ( .A(KEYINPUT46), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n715), .A2(n714), .ZN(n579) );
  INV_X1 U674 ( .A(n580), .ZN(n582) );
  NAND2_X1 U675 ( .A1(G953), .A2(G900), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n631), .A2(n701), .ZN(n583) );
  XNOR2_X1 U678 ( .A(KEYINPUT30), .B(n583), .ZN(n584) );
  NOR2_X1 U679 ( .A1(n590), .A2(n584), .ZN(n585) );
  XNOR2_X1 U680 ( .A(n586), .B(KEYINPUT38), .ZN(n702) );
  NAND2_X1 U681 ( .A1(n610), .A2(n702), .ZN(n588) );
  INV_X1 U682 ( .A(KEYINPUT39), .ZN(n587) );
  XNOR2_X1 U683 ( .A(n588), .B(n587), .ZN(n626) );
  NOR2_X1 U684 ( .A1(n626), .A2(n609), .ZN(n589) );
  XNOR2_X1 U685 ( .A(n589), .B(KEYINPUT40), .ZN(n787) );
  NAND2_X1 U686 ( .A1(n593), .A2(n592), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U688 ( .A1(n704), .A2(n524), .ZN(n596) );
  XNOR2_X1 U689 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n595) );
  XNOR2_X1 U690 ( .A(n596), .B(n595), .ZN(n733) );
  NOR2_X1 U691 ( .A1(n607), .A2(n733), .ZN(n597) );
  XNOR2_X1 U692 ( .A(n597), .B(KEYINPUT42), .ZN(n786) );
  XNOR2_X1 U693 ( .A(n618), .B(KEYINPUT115), .ZN(n602) );
  INV_X1 U694 ( .A(n605), .ZN(n606) );
  AND2_X1 U695 ( .A1(n611), .A2(n608), .ZN(n679) );
  INV_X1 U696 ( .A(n679), .ZN(n689) );
  NAND2_X1 U697 ( .A1(n689), .A2(n609), .ZN(n636) );
  INV_X1 U698 ( .A(n636), .ZN(n705) );
  INV_X1 U699 ( .A(n610), .ZN(n613) );
  AND2_X1 U700 ( .A1(n457), .A2(n611), .ZN(n645) );
  INV_X1 U701 ( .A(n586), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n645), .A2(n622), .ZN(n612) );
  NOR2_X1 U703 ( .A1(n613), .A2(n612), .ZN(n682) );
  AND2_X1 U704 ( .A1(KEYINPUT47), .A2(n705), .ZN(n614) );
  NOR2_X1 U705 ( .A1(KEYINPUT90), .A2(n614), .ZN(n615) );
  XNOR2_X1 U706 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n621) );
  INV_X1 U707 ( .A(n710), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n618), .A2(n701), .ZN(n619) );
  NOR2_X1 U709 ( .A1(n641), .A2(n619), .ZN(n620) );
  XNOR2_X1 U710 ( .A(n621), .B(n620), .ZN(n623) );
  NOR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n694) );
  INV_X1 U712 ( .A(n694), .ZN(n624) );
  INV_X1 U713 ( .A(KEYINPUT92), .ZN(n625) );
  OR2_X1 U714 ( .A1(n626), .A2(n689), .ZN(n693) );
  INV_X1 U715 ( .A(n627), .ZN(n629) );
  INV_X1 U716 ( .A(n628), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n630), .B(KEYINPUT104), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n632), .A2(n591), .ZN(n675) );
  OR2_X1 U719 ( .A1(n406), .A2(n591), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n709), .A2(n375), .ZN(n635) );
  INV_X1 U721 ( .A(KEYINPUT31), .ZN(n634) );
  NAND2_X1 U722 ( .A1(n675), .A2(n688), .ZN(n637) );
  INV_X1 U723 ( .A(KEYINPUT110), .ZN(n638) );
  XNOR2_X1 U724 ( .A(n639), .B(n638), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U726 ( .A1(n642), .A2(n711), .ZN(n643) );
  XNOR2_X1 U727 ( .A(KEYINPUT85), .B(KEYINPUT35), .ZN(n646) );
  XNOR2_X2 U728 ( .A(n647), .B(n646), .ZN(n785) );
  AND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n785), .A2(n655), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n652), .B(KEYINPUT95), .ZN(n659) );
  INV_X1 U732 ( .A(KEYINPUT44), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n785), .A2(n653), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(KEYINPUT65), .ZN(n657) );
  XNOR2_X1 U735 ( .A(n655), .B(KEYINPUT96), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U738 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n660) );
  XNOR2_X2 U739 ( .A(n661), .B(n660), .ZN(n760) );
  INV_X1 U740 ( .A(KEYINPUT2), .ZN(n697) );
  XNOR2_X1 U741 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n668), .B(n667), .ZN(n670) );
  INV_X1 U743 ( .A(G952), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U745 ( .A(KEYINPUT62), .B(n672), .Z(n673) );
  INV_X1 U746 ( .A(n683), .ZN(n686) );
  NOR2_X1 U747 ( .A1(n686), .A2(n675), .ZN(n674) );
  XOR2_X1 U748 ( .A(G104), .B(n674), .Z(G6) );
  NOR2_X1 U749 ( .A1(n689), .A2(n675), .ZN(n677) );
  XNOR2_X1 U750 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U752 ( .A(G107), .B(n678), .ZN(G9) );
  XOR2_X1 U753 ( .A(G128), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U754 ( .A1(n679), .A2(n684), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n681), .B(n680), .ZN(G30) );
  XOR2_X1 U756 ( .A(G143), .B(n682), .Z(G45) );
  NAND2_X1 U757 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n685), .B(G146), .ZN(G48) );
  NOR2_X1 U759 ( .A1(n686), .A2(n688), .ZN(n687) );
  XOR2_X1 U760 ( .A(G113), .B(n687), .Z(G15) );
  NOR2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U762 ( .A(G116), .B(n690), .Z(G18) );
  XNOR2_X1 U763 ( .A(n691), .B(G125), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U765 ( .A(G134), .B(n693), .ZN(G36) );
  XOR2_X1 U766 ( .A(G140), .B(n694), .Z(n695) );
  XNOR2_X1 U767 ( .A(KEYINPUT118), .B(n695), .ZN(G42) );
  XNOR2_X1 U768 ( .A(KEYINPUT89), .B(n697), .ZN(n698) );
  NOR2_X1 U769 ( .A1(n696), .A2(n698), .ZN(n699) );
  NOR2_X1 U770 ( .A1(n700), .A2(n699), .ZN(n738) );
  NOR2_X1 U771 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U772 ( .A1(n524), .A2(n703), .ZN(n707) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U775 ( .A1(n708), .A2(n732), .ZN(n726) );
  INV_X1 U776 ( .A(n709), .ZN(n722) );
  XOR2_X1 U777 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n713) );
  NAND2_X1 U778 ( .A1(n711), .A2(n406), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n713), .B(n712), .ZN(n719) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n717) );
  XNOR2_X1 U781 ( .A(KEYINPUT119), .B(KEYINPUT49), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U784 ( .A1(n720), .A2(n591), .ZN(n721) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U786 ( .A(KEYINPUT51), .B(n723), .ZN(n724) );
  NOR2_X1 U787 ( .A1(n733), .A2(n724), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U789 ( .A(KEYINPUT52), .B(n727), .ZN(n730) );
  NAND2_X1 U790 ( .A1(G952), .A2(n728), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U792 ( .A1(G953), .A2(n731), .ZN(n736) );
  NOR2_X1 U793 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U794 ( .A(n734), .B(KEYINPUT121), .ZN(n735) );
  NAND2_X1 U795 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U796 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U797 ( .A(KEYINPUT53), .B(n739), .ZN(G75) );
  XOR2_X1 U798 ( .A(KEYINPUT88), .B(KEYINPUT54), .Z(n740) );
  XNOR2_X1 U799 ( .A(n740), .B(KEYINPUT98), .ZN(n742) );
  XOR2_X1 U800 ( .A(KEYINPUT97), .B(KEYINPUT55), .Z(n741) );
  XNOR2_X1 U801 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U802 ( .A1(n755), .A2(G469), .ZN(n748) );
  XOR2_X1 U803 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n746) );
  NOR2_X1 U804 ( .A1(n759), .A2(n749), .ZN(G54) );
  NAND2_X1 U805 ( .A1(n755), .A2(G478), .ZN(n753) );
  INV_X1 U806 ( .A(KEYINPUT123), .ZN(n750) );
  XNOR2_X1 U807 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U808 ( .A(n753), .B(n752), .ZN(n754) );
  NOR2_X1 U809 ( .A1(n759), .A2(n754), .ZN(G63) );
  NAND2_X1 U810 ( .A1(n755), .A2(G217), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(n756), .ZN(n758) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(G66) );
  NAND2_X1 U813 ( .A1(n760), .A2(n781), .ZN(n764) );
  NAND2_X1 U814 ( .A1(G953), .A2(G224), .ZN(n761) );
  XNOR2_X1 U815 ( .A(KEYINPUT61), .B(n761), .ZN(n762) );
  NAND2_X1 U816 ( .A1(n762), .A2(n767), .ZN(n763) );
  NAND2_X1 U817 ( .A1(n764), .A2(n763), .ZN(n771) );
  XOR2_X1 U818 ( .A(n766), .B(n765), .Z(n769) );
  NOR2_X1 U819 ( .A1(n767), .A2(n781), .ZN(n768) );
  NOR2_X1 U820 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(G69) );
  XOR2_X1 U822 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n775) );
  XNOR2_X1 U823 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U824 ( .A(n775), .B(n774), .ZN(n780) );
  XNOR2_X1 U825 ( .A(G227), .B(n780), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U827 ( .A1(n777), .A2(G953), .ZN(n778) );
  XNOR2_X1 U828 ( .A(n778), .B(KEYINPUT126), .ZN(n784) );
  XNOR2_X1 U829 ( .A(n780), .B(n779), .ZN(n782) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n784), .A2(n783), .ZN(G72) );
  XNOR2_X1 U832 ( .A(n785), .B(G122), .ZN(G24) );
  XOR2_X1 U833 ( .A(G137), .B(n786), .Z(G39) );
  XNOR2_X1 U834 ( .A(G131), .B(KEYINPUT127), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n788), .B(n787), .ZN(G33) );
endmodule

